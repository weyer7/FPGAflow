magic
tech sky130A
magscale 1 2
timestamp 1745537824
<< viali >>
rect 6101 28713 6135 28747
rect 6561 28713 6595 28747
rect 9873 28713 9907 28747
rect 3341 28577 3375 28611
rect 4905 28509 4939 28543
rect 5917 28509 5951 28543
rect 6377 28509 6411 28543
rect 8125 28509 8159 28543
rect 8677 28509 8711 28543
rect 9505 28509 9539 28543
rect 9689 28509 9723 28543
rect 12357 28509 12391 28543
rect 12541 28509 12575 28543
rect 17049 28509 17083 28543
rect 17233 28509 17267 28543
rect 4721 28441 4755 28475
rect 7880 28441 7914 28475
rect 8953 28441 8987 28475
rect 5089 28373 5123 28407
rect 6745 28373 6779 28407
rect 8493 28373 8527 28407
rect 12449 28373 12483 28407
rect 17141 28373 17175 28407
rect 4629 28169 4663 28203
rect 6193 28169 6227 28203
rect 6929 28169 6963 28203
rect 7389 28169 7423 28203
rect 9137 28169 9171 28203
rect 9321 28169 9355 28203
rect 18061 28169 18095 28203
rect 2780 28101 2814 28135
rect 4261 28101 4295 28135
rect 6561 28101 6595 28135
rect 8024 28101 8058 28135
rect 16313 28101 16347 28135
rect 1685 28033 1719 28067
rect 1869 28033 1903 28067
rect 4470 28033 4504 28067
rect 4721 28033 4755 28067
rect 4997 28033 5031 28067
rect 5549 28033 5583 28067
rect 5687 28033 5721 28067
rect 5825 28033 5859 28067
rect 5917 28033 5951 28067
rect 6009 28033 6043 28067
rect 6377 28033 6411 28067
rect 6653 28033 6687 28067
rect 6745 28033 6779 28067
rect 7205 28033 7239 28067
rect 10434 28033 10468 28067
rect 10977 28033 11011 28067
rect 11805 28033 11839 28067
rect 12633 28033 12667 28067
rect 12889 28033 12923 28067
rect 14473 28033 14507 28067
rect 14740 28033 14774 28067
rect 16497 28033 16531 28067
rect 16681 28033 16715 28067
rect 16937 28033 16971 28067
rect 19277 28033 19311 28067
rect 19533 28033 19567 28067
rect 2513 27965 2547 27999
rect 3985 27965 4019 27999
rect 4353 27965 4387 27999
rect 4813 27965 4847 27999
rect 7757 27965 7791 27999
rect 10701 27965 10735 27999
rect 11069 27965 11103 27999
rect 12449 27965 12483 27999
rect 19625 27965 19659 27999
rect 20177 27965 20211 27999
rect 5181 27897 5215 27931
rect 1685 27829 1719 27863
rect 3893 27829 3927 27863
rect 4813 27829 4847 27863
rect 11345 27829 11379 27863
rect 14013 27829 14047 27863
rect 15853 27829 15887 27863
rect 16129 27829 16163 27863
rect 18153 27829 18187 27863
rect 3157 27625 3191 27659
rect 4537 27625 4571 27659
rect 6193 27625 6227 27659
rect 12909 27625 12943 27659
rect 16221 27625 16255 27659
rect 4813 27557 4847 27591
rect 6285 27557 6319 27591
rect 10425 27557 10459 27591
rect 13921 27557 13955 27591
rect 16405 27557 16439 27591
rect 17693 27557 17727 27591
rect 1409 27489 1443 27523
rect 3065 27489 3099 27523
rect 9689 27489 9723 27523
rect 10333 27489 10367 27523
rect 10701 27489 10735 27523
rect 11253 27489 11287 27523
rect 13553 27489 13587 27523
rect 14657 27489 14691 27523
rect 17233 27489 17267 27523
rect 18337 27489 18371 27523
rect 1676 27421 1710 27455
rect 2973 27421 3007 27455
rect 3433 27421 3467 27455
rect 3617 27421 3651 27455
rect 4353 27421 4387 27455
rect 4813 27421 4847 27455
rect 4997 27421 5031 27455
rect 6193 27421 6227 27455
rect 7389 27421 7423 27455
rect 10793 27421 10827 27455
rect 11509 27421 11543 27455
rect 13645 27421 13679 27455
rect 13737 27421 13771 27455
rect 15761 27421 15795 27455
rect 17325 27421 17359 27455
rect 17785 27421 17819 27455
rect 3249 27353 3283 27387
rect 6561 27353 6595 27387
rect 7656 27353 7690 27387
rect 13921 27353 13955 27387
rect 14105 27353 14139 27387
rect 16037 27353 16071 27387
rect 16237 27353 16271 27387
rect 2789 27285 2823 27319
rect 3801 27285 3835 27319
rect 6469 27285 6503 27319
rect 8769 27285 8803 27319
rect 12633 27285 12667 27319
rect 15117 27285 15151 27319
rect 1685 27081 1719 27115
rect 2053 27081 2087 27115
rect 3157 27081 3191 27115
rect 7941 27081 7975 27115
rect 15761 27081 15795 27115
rect 20821 27081 20855 27115
rect 4721 27013 4755 27047
rect 8109 27013 8143 27047
rect 8309 27013 8343 27047
rect 13353 27013 13387 27047
rect 13553 27013 13587 27047
rect 13813 27013 13847 27047
rect 14013 27013 14047 27047
rect 18429 27013 18463 27047
rect 18858 27013 18892 27047
rect 1961 26945 1995 26979
rect 2237 26945 2271 26979
rect 2421 26945 2455 26979
rect 2605 26945 2639 26979
rect 2697 26945 2731 26979
rect 2973 26945 3007 26979
rect 3249 26945 3283 26979
rect 4537 26945 4571 26979
rect 5273 26945 5307 26979
rect 7205 26945 7239 26979
rect 9229 26945 9263 26979
rect 9321 26945 9355 26979
rect 9505 26945 9539 26979
rect 12449 26945 12483 26979
rect 12909 26945 12943 26979
rect 14289 26945 14323 26979
rect 15485 26945 15519 26979
rect 15945 26945 15979 26979
rect 16221 26945 16255 26979
rect 18337 26945 18371 26979
rect 18521 26945 18555 26979
rect 18613 26945 18647 26979
rect 21005 26945 21039 26979
rect 1685 26877 1719 26911
rect 2881 26877 2915 26911
rect 9965 26877 9999 26911
rect 12817 26877 12851 26911
rect 14197 26877 14231 26911
rect 14657 26877 14691 26911
rect 16129 26877 16163 26911
rect 17141 26877 17175 26911
rect 20637 26877 20671 26911
rect 21189 26877 21223 26911
rect 2789 26809 2823 26843
rect 9505 26809 9539 26843
rect 13093 26809 13127 26843
rect 17509 26809 17543 26843
rect 19993 26809 20027 26843
rect 1869 26741 1903 26775
rect 2973 26741 3007 26775
rect 4905 26741 4939 26775
rect 5181 26741 5215 26775
rect 7113 26741 7147 26775
rect 8125 26741 8159 26775
rect 10609 26741 10643 26775
rect 12633 26741 12667 26775
rect 13185 26741 13219 26775
rect 13369 26741 13403 26775
rect 13645 26741 13679 26775
rect 13829 26741 13863 26775
rect 14933 26741 14967 26775
rect 15945 26741 15979 26775
rect 17601 26741 17635 26775
rect 20085 26741 20119 26775
rect 1869 26537 1903 26571
rect 4077 26537 4111 26571
rect 4537 26537 4571 26571
rect 5549 26537 5583 26571
rect 6469 26537 6503 26571
rect 6561 26537 6595 26571
rect 7389 26537 7423 26571
rect 7849 26537 7883 26571
rect 8217 26537 8251 26571
rect 13737 26537 13771 26571
rect 15485 26537 15519 26571
rect 16313 26537 16347 26571
rect 16497 26537 16531 26571
rect 16681 26537 16715 26571
rect 19625 26537 19659 26571
rect 7205 26469 7239 26503
rect 13185 26469 13219 26503
rect 4261 26401 4295 26435
rect 5273 26401 5307 26435
rect 6837 26401 6871 26435
rect 6930 26401 6964 26435
rect 8401 26401 8435 26435
rect 14105 26401 14139 26435
rect 1685 26333 1719 26367
rect 2053 26333 2087 26367
rect 2881 26333 2915 26367
rect 3065 26333 3099 26367
rect 3985 26333 4019 26367
rect 4629 26333 4663 26367
rect 4787 26333 4821 26367
rect 4905 26333 4939 26367
rect 4997 26333 5031 26367
rect 5089 26333 5123 26367
rect 5733 26333 5767 26367
rect 6193 26333 6227 26367
rect 6285 26333 6319 26367
rect 6719 26333 6753 26367
rect 7021 26333 7055 26367
rect 7481 26333 7515 26367
rect 7573 26333 7607 26367
rect 7849 26333 7883 26367
rect 7941 26333 7975 26367
rect 8493 26333 8527 26367
rect 8585 26333 8619 26367
rect 8677 26333 8711 26367
rect 10445 26333 10479 26367
rect 10701 26333 10735 26367
rect 10793 26333 10827 26367
rect 12541 26333 12575 26367
rect 13461 26333 13495 26367
rect 15853 26333 15887 26367
rect 15945 26333 15979 26367
rect 16313 26333 16347 26367
rect 18438 26333 18472 26367
rect 18705 26333 18739 26367
rect 19625 26333 19659 26367
rect 19809 26333 19843 26367
rect 5917 26265 5951 26299
rect 6469 26265 6503 26299
rect 11060 26265 11094 26299
rect 13093 26265 13127 26299
rect 13185 26265 13219 26299
rect 13553 26265 13587 26299
rect 14350 26265 14384 26299
rect 16865 26265 16899 26299
rect 16957 26265 16991 26299
rect 17233 26265 17267 26299
rect 1501 26197 1535 26231
rect 2881 26197 2915 26231
rect 6009 26197 6043 26231
rect 9321 26197 9355 26231
rect 12173 26197 12207 26231
rect 13369 26197 13403 26231
rect 13753 26197 13787 26231
rect 13921 26197 13955 26231
rect 17049 26197 17083 26231
rect 17325 26197 17359 26231
rect 2053 25993 2087 26027
rect 2237 25993 2271 26027
rect 4077 25993 4111 26027
rect 5549 25993 5583 26027
rect 6745 25993 6779 26027
rect 7205 25993 7239 26027
rect 8953 25993 8987 26027
rect 9321 25993 9355 26027
rect 11253 25993 11287 26027
rect 12985 25993 13019 26027
rect 13737 25993 13771 26027
rect 14105 25993 14139 26027
rect 14473 25993 14507 26027
rect 16129 25993 16163 26027
rect 17509 25993 17543 26027
rect 21097 25993 21131 26027
rect 2881 25925 2915 25959
rect 6377 25925 6411 25959
rect 7389 25925 7423 25959
rect 13185 25925 13219 25959
rect 15485 25925 15519 25959
rect 16313 25925 16347 25959
rect 20729 25925 20763 25959
rect 20929 25925 20963 25959
rect 1869 25857 1903 25891
rect 2145 25857 2179 25891
rect 2421 25857 2455 25891
rect 3341 25857 3375 25891
rect 3433 25857 3467 25891
rect 3801 25857 3835 25891
rect 4261 25857 4295 25891
rect 4353 25857 4387 25891
rect 5273 25857 5307 25891
rect 6561 25857 6595 25891
rect 7113 25857 7147 25891
rect 8125 25857 8159 25891
rect 8217 25857 8251 25891
rect 8309 25857 8343 25891
rect 8493 25857 8527 25891
rect 8769 25857 8803 25891
rect 9505 25857 9539 25891
rect 9597 25857 9631 25891
rect 11161 25857 11195 25891
rect 11345 25857 11379 25891
rect 12081 25857 12115 25891
rect 12725 25857 12759 25891
rect 13553 25857 13587 25891
rect 13645 25857 13679 25891
rect 14289 25857 14323 25891
rect 14565 25857 14599 25891
rect 15761 25857 15795 25891
rect 15945 25857 15979 25891
rect 16405 25857 16439 25891
rect 17141 25857 17175 25891
rect 17325 25857 17359 25891
rect 20637 25857 20671 25891
rect 21189 25857 21223 25891
rect 21373 25857 21407 25891
rect 2605 25789 2639 25823
rect 4445 25789 4479 25823
rect 4537 25789 4571 25823
rect 5365 25789 5399 25823
rect 5549 25789 5583 25823
rect 9321 25789 9355 25823
rect 13277 25789 13311 25823
rect 17049 25789 17083 25823
rect 17233 25789 17267 25823
rect 18153 25789 18187 25823
rect 19993 25789 20027 25823
rect 3985 25721 4019 25755
rect 12817 25721 12851 25755
rect 17601 25721 17635 25755
rect 1685 25653 1719 25687
rect 2789 25653 2823 25687
rect 3709 25653 3743 25687
rect 7389 25653 7423 25687
rect 7849 25653 7883 25687
rect 13001 25653 13035 25687
rect 13369 25653 13403 25687
rect 13461 25653 13495 25687
rect 15945 25653 15979 25687
rect 20913 25653 20947 25687
rect 21189 25653 21223 25687
rect 4261 25449 4295 25483
rect 4629 25449 4663 25483
rect 5733 25449 5767 25483
rect 13093 25449 13127 25483
rect 16313 25449 16347 25483
rect 19625 25449 19659 25483
rect 21097 25449 21131 25483
rect 1501 25381 1535 25415
rect 5825 25381 5859 25415
rect 1869 25313 1903 25347
rect 5365 25313 5399 25347
rect 6745 25313 6779 25347
rect 6837 25313 6871 25347
rect 7297 25313 7331 25347
rect 9689 25313 9723 25347
rect 11713 25313 11747 25347
rect 13185 25313 13219 25347
rect 19717 25313 19751 25347
rect 21741 25313 21775 25347
rect 1685 25245 1719 25279
rect 1777 25245 1811 25279
rect 1961 25245 1995 25279
rect 3893 25245 3927 25279
rect 3985 25245 4019 25279
rect 4353 25245 4387 25279
rect 4813 25245 4847 25279
rect 4905 25245 4939 25279
rect 4997 25245 5031 25279
rect 5089 25245 5123 25279
rect 5273 25245 5307 25279
rect 5641 25245 5675 25279
rect 5917 25245 5951 25279
rect 6101 25245 6135 25279
rect 6377 25245 6411 25279
rect 6469 25245 6503 25279
rect 8125 25245 8159 25279
rect 10149 25245 10183 25279
rect 15577 25245 15611 25279
rect 19349 25245 19383 25279
rect 19625 25245 19659 25279
rect 21189 25245 21223 25279
rect 10416 25177 10450 25211
rect 11980 25177 12014 25211
rect 16497 25177 16531 25211
rect 19984 25177 20018 25211
rect 4537 25109 4571 25143
rect 6193 25109 6227 25143
rect 6561 25109 6595 25143
rect 7941 25109 7975 25143
rect 8217 25109 8251 25143
rect 9137 25109 9171 25143
rect 11529 25109 11563 25143
rect 13829 25109 13863 25143
rect 15485 25109 15519 25143
rect 16129 25109 16163 25143
rect 16297 25109 16331 25143
rect 19441 25109 19475 25143
rect 2697 24905 2731 24939
rect 7665 24905 7699 24939
rect 8677 24905 8711 24939
rect 16497 24905 16531 24939
rect 19993 24905 20027 24939
rect 2865 24837 2899 24871
rect 3065 24837 3099 24871
rect 5549 24837 5583 24871
rect 1685 24769 1719 24803
rect 1869 24769 1903 24803
rect 2053 24769 2087 24803
rect 4077 24769 4111 24803
rect 4445 24769 4479 24803
rect 4629 24769 4663 24803
rect 5365 24769 5399 24803
rect 5641 24769 5675 24803
rect 5825 24769 5859 24803
rect 6009 24769 6043 24803
rect 6377 24769 6411 24803
rect 6561 24769 6595 24803
rect 6745 24769 6779 24803
rect 6837 24769 6871 24803
rect 6929 24769 6963 24803
rect 7297 24769 7331 24803
rect 7481 24769 7515 24803
rect 7573 24769 7607 24803
rect 7849 24769 7883 24803
rect 8033 24769 8067 24803
rect 8217 24769 8251 24803
rect 8401 24769 8435 24803
rect 8585 24769 8619 24803
rect 9790 24769 9824 24803
rect 10241 24769 10275 24803
rect 10425 24769 10459 24803
rect 12725 24769 12759 24803
rect 14657 24769 14691 24803
rect 15384 24769 15418 24803
rect 18254 24769 18288 24803
rect 18521 24769 18555 24803
rect 18613 24769 18647 24803
rect 18869 24769 18903 24803
rect 20637 24769 20671 24803
rect 4353 24701 4387 24735
rect 5917 24701 5951 24735
rect 8125 24701 8159 24735
rect 10057 24701 10091 24735
rect 11529 24701 11563 24735
rect 15117 24701 15151 24735
rect 1501 24633 1535 24667
rect 3893 24633 3927 24667
rect 5365 24633 5399 24667
rect 13369 24633 13403 24667
rect 17141 24633 17175 24667
rect 2053 24565 2087 24599
rect 2881 24565 2915 24599
rect 4261 24565 4295 24599
rect 4537 24565 4571 24599
rect 7113 24565 7147 24599
rect 7389 24565 7423 24599
rect 10333 24565 10367 24599
rect 12173 24565 12207 24599
rect 20085 24565 20119 24599
rect 2973 24361 3007 24395
rect 3433 24361 3467 24395
rect 8033 24361 8067 24395
rect 8309 24361 8343 24395
rect 12449 24361 12483 24395
rect 16865 24361 16899 24395
rect 18705 24361 18739 24395
rect 21097 24361 21131 24395
rect 2789 24293 2823 24327
rect 1409 24225 1443 24259
rect 2881 24225 2915 24259
rect 6377 24225 6411 24259
rect 6469 24225 6503 24259
rect 6561 24225 6595 24259
rect 12357 24225 12391 24259
rect 16405 24225 16439 24259
rect 17509 24225 17543 24259
rect 19717 24225 19751 24259
rect 21741 24225 21775 24259
rect 1676 24157 1710 24191
rect 3065 24157 3099 24191
rect 3157 24157 3191 24191
rect 3341 24157 3375 24191
rect 6009 24157 6043 24191
rect 6653 24157 6687 24191
rect 6837 24157 6871 24191
rect 7757 24157 7791 24191
rect 7941 24157 7975 24191
rect 8309 24157 8343 24191
rect 8401 24157 8435 24191
rect 8677 24157 8711 24191
rect 12090 24157 12124 24191
rect 12633 24157 12667 24191
rect 12725 24157 12759 24191
rect 12817 24157 12851 24191
rect 13001 24157 13035 24191
rect 13093 24157 13127 24191
rect 13553 24157 13587 24191
rect 14105 24157 14139 24191
rect 16129 24157 16163 24191
rect 16497 24157 16531 24191
rect 16957 24157 16991 24191
rect 18797 24157 18831 24191
rect 8953 24089 8987 24123
rect 12449 24089 12483 24123
rect 14372 24089 14406 24123
rect 19962 24089 19996 24123
rect 5825 24021 5859 24055
rect 6193 24021 6227 24055
rect 7757 24021 7791 24055
rect 10241 24021 10275 24055
rect 10977 24021 11011 24055
rect 12909 24021 12943 24055
rect 13369 24021 13403 24055
rect 13461 24021 13495 24055
rect 15485 24021 15519 24055
rect 15577 24021 15611 24055
rect 21189 24021 21223 24055
rect 1501 23817 1535 23851
rect 2789 23817 2823 23851
rect 3341 23817 3375 23851
rect 4813 23817 4847 23851
rect 7021 23817 7055 23851
rect 7205 23817 7239 23851
rect 14657 23817 14691 23851
rect 15301 23817 15335 23851
rect 15469 23817 15503 23851
rect 16129 23817 16163 23851
rect 2605 23749 2639 23783
rect 4454 23749 4488 23783
rect 5948 23749 5982 23783
rect 9873 23749 9907 23783
rect 10241 23749 10275 23783
rect 12716 23749 12750 23783
rect 15669 23749 15703 23783
rect 1685 23681 1719 23715
rect 1961 23681 1995 23715
rect 2513 23681 2547 23715
rect 2697 23681 2731 23715
rect 2973 23681 3007 23715
rect 8217 23681 8251 23715
rect 10057 23681 10091 23715
rect 10517 23681 10551 23715
rect 10977 23681 11011 23715
rect 11161 23681 11195 23715
rect 11253 23681 11287 23715
rect 12081 23681 12115 23715
rect 14841 23681 14875 23715
rect 15025 23681 15059 23715
rect 15117 23681 15151 23715
rect 15945 23681 15979 23715
rect 16221 23681 16255 23715
rect 19441 23681 19475 23715
rect 3157 23613 3191 23647
rect 4721 23613 4755 23647
rect 6193 23613 6227 23647
rect 10425 23613 10459 23647
rect 12449 23613 12483 23647
rect 14473 23613 14507 23647
rect 19533 23613 19567 23647
rect 19809 23613 19843 23647
rect 7573 23545 7607 23579
rect 8401 23545 8435 23579
rect 11529 23545 11563 23579
rect 13829 23545 13863 23579
rect 1777 23477 1811 23511
rect 7205 23477 7239 23511
rect 10793 23477 10827 23511
rect 13921 23477 13955 23511
rect 15485 23477 15519 23511
rect 15761 23477 15795 23511
rect 3893 23273 3927 23307
rect 3985 23273 4019 23307
rect 12817 23273 12851 23307
rect 12909 23273 12943 23307
rect 13093 23273 13127 23307
rect 21557 23273 21591 23307
rect 20637 23205 20671 23239
rect 3801 23137 3835 23171
rect 7849 23137 7883 23171
rect 9689 23137 9723 23171
rect 13461 23137 13495 23171
rect 13921 23137 13955 23171
rect 19257 23137 19291 23171
rect 20821 23137 20855 23171
rect 3249 23069 3283 23103
rect 4077 23069 4111 23103
rect 5273 23069 5307 23103
rect 7481 23069 7515 23103
rect 7665 23069 7699 23103
rect 9229 23069 9263 23103
rect 9597 23069 9631 23103
rect 9781 23069 9815 23103
rect 9873 23069 9907 23103
rect 12541 23069 12575 23103
rect 12817 23069 12851 23103
rect 13553 23069 13587 23103
rect 14105 23069 14139 23103
rect 14657 23069 14691 23103
rect 15393 23069 15427 23103
rect 17141 23069 17175 23103
rect 17417 23069 17451 23103
rect 20913 23069 20947 23103
rect 21373 23069 21407 23103
rect 13061 23001 13095 23035
rect 13277 23001 13311 23035
rect 17662 23001 17696 23035
rect 19502 23001 19536 23035
rect 2697 22933 2731 22967
rect 9045 22933 9079 22967
rect 9413 22933 9447 22967
rect 12633 22933 12667 22967
rect 18797 22933 18831 22967
rect 21281 22933 21315 22967
rect 6837 22729 6871 22763
rect 8769 22729 8803 22763
rect 9321 22729 9355 22763
rect 10793 22729 10827 22763
rect 11713 22729 11747 22763
rect 11805 22729 11839 22763
rect 14381 22729 14415 22763
rect 16405 22729 16439 22763
rect 18981 22729 19015 22763
rect 21281 22729 21315 22763
rect 2504 22661 2538 22695
rect 9658 22661 9692 22695
rect 10885 22661 10919 22695
rect 15494 22661 15528 22695
rect 16037 22661 16071 22695
rect 16926 22661 16960 22695
rect 18245 22661 18279 22695
rect 19257 22661 19291 22695
rect 19625 22661 19659 22695
rect 2237 22593 2271 22627
rect 5080 22593 5114 22627
rect 6653 22593 6687 22627
rect 7656 22593 7690 22627
rect 9413 22593 9447 22627
rect 11069 22593 11103 22627
rect 11161 22593 11195 22627
rect 11897 22593 11931 22627
rect 12449 22593 12483 22627
rect 12541 22593 12575 22627
rect 15853 22593 15887 22627
rect 16129 22593 16163 22627
rect 16221 22593 16255 22627
rect 16681 22593 16715 22627
rect 19165 22593 19199 22627
rect 19349 22593 19383 22627
rect 19533 22593 19567 22627
rect 21189 22593 21223 22627
rect 22201 22593 22235 22627
rect 4445 22525 4479 22559
rect 4813 22525 4847 22559
rect 6469 22525 6503 22559
rect 7389 22525 7423 22559
rect 8861 22525 8895 22559
rect 11529 22525 11563 22559
rect 13645 22525 13679 22559
rect 15761 22525 15795 22559
rect 18797 22525 18831 22559
rect 20269 22525 20303 22559
rect 21373 22525 21407 22559
rect 21833 22525 21867 22559
rect 22109 22525 22143 22559
rect 3617 22457 3651 22491
rect 6193 22457 6227 22491
rect 9229 22457 9263 22491
rect 12725 22457 12759 22491
rect 20821 22457 20855 22491
rect 3893 22389 3927 22423
rect 10885 22389 10919 22423
rect 11345 22389 11379 22423
rect 12081 22389 12115 22423
rect 12265 22389 12299 22423
rect 13093 22389 13127 22423
rect 18061 22389 18095 22423
rect 2789 22185 2823 22219
rect 5549 22185 5583 22219
rect 7573 22185 7607 22219
rect 7757 22185 7791 22219
rect 12449 22185 12483 22219
rect 13645 22185 13679 22219
rect 17325 22185 17359 22219
rect 10425 22117 10459 22151
rect 13461 22117 13495 22151
rect 13553 22117 13587 22151
rect 1409 22049 1443 22083
rect 3801 22049 3835 22083
rect 13001 22049 13035 22083
rect 19257 22049 19291 22083
rect 1676 21981 1710 22015
rect 4057 21981 4091 22015
rect 7113 21981 7147 22015
rect 7389 21981 7423 22015
rect 8033 21981 8067 22015
rect 8401 21981 8435 22015
rect 8493 21981 8527 22015
rect 9873 21981 9907 22015
rect 10241 21981 10275 22015
rect 11437 21981 11471 22015
rect 11621 21981 11655 22015
rect 11897 21981 11931 22015
rect 11989 21981 12023 22015
rect 13369 21981 13403 22015
rect 13829 21981 13863 22015
rect 14105 21981 14139 22015
rect 14381 21981 14415 22015
rect 15577 21981 15611 22015
rect 15761 21981 15795 22015
rect 16773 21981 16807 22015
rect 17049 21981 17083 22015
rect 17187 21981 17221 22015
rect 17601 21981 17635 22015
rect 17877 21981 17911 22015
rect 18245 21981 18279 22015
rect 18337 21981 18371 22015
rect 18521 21981 18555 22015
rect 18705 21981 18739 22015
rect 20821 21981 20855 22015
rect 7021 21913 7055 21947
rect 7757 21913 7791 21947
rect 7941 21913 7975 21947
rect 10057 21913 10091 21947
rect 11713 21913 11747 21947
rect 12265 21913 12299 21947
rect 12465 21913 12499 21947
rect 12817 21913 12851 21947
rect 14473 21913 14507 21947
rect 16957 21913 16991 21947
rect 18613 21913 18647 21947
rect 19502 21913 19536 21947
rect 5181 21845 5215 21879
rect 7205 21845 7239 21879
rect 10149 21845 10183 21879
rect 11529 21845 11563 21879
rect 11811 21845 11845 21879
rect 12633 21845 12667 21879
rect 13093 21845 13127 21879
rect 14289 21845 14323 21879
rect 14657 21845 14691 21879
rect 15669 21845 15703 21879
rect 17417 21845 17451 21879
rect 17785 21845 17819 21879
rect 18061 21845 18095 21879
rect 18889 21845 18923 21879
rect 20637 21845 20671 21879
rect 20913 21845 20947 21879
rect 5457 21641 5491 21675
rect 7205 21641 7239 21675
rect 8861 21641 8895 21675
rect 13921 21641 13955 21675
rect 15853 21641 15887 21675
rect 16681 21641 16715 21675
rect 18429 21641 18463 21675
rect 19625 21641 19659 21675
rect 21833 21641 21867 21675
rect 22661 21641 22695 21675
rect 7748 21573 7782 21607
rect 12173 21573 12207 21607
rect 12786 21573 12820 21607
rect 14565 21573 14599 21607
rect 14781 21573 14815 21607
rect 15301 21573 15335 21607
rect 16957 21573 16991 21607
rect 1409 21505 1443 21539
rect 2329 21505 2363 21539
rect 2596 21505 2630 21539
rect 4997 21505 5031 21539
rect 5090 21505 5124 21539
rect 5825 21505 5859 21539
rect 6653 21505 6687 21539
rect 7113 21505 7147 21539
rect 7297 21505 7331 21539
rect 7481 21505 7515 21539
rect 8953 21505 8987 21539
rect 11897 21505 11931 21539
rect 12081 21505 12115 21539
rect 12265 21505 12299 21539
rect 12541 21505 12575 21539
rect 15025 21505 15059 21539
rect 15117 21505 15151 21539
rect 15393 21505 15427 21539
rect 15531 21505 15565 21539
rect 15853 21505 15887 21539
rect 16129 21505 16163 21539
rect 16865 21505 16899 21539
rect 17049 21505 17083 21539
rect 17187 21505 17221 21539
rect 17417 21505 17451 21539
rect 17969 21505 18003 21539
rect 18705 21505 18739 21539
rect 20177 21505 20211 21539
rect 22109 21505 22143 21539
rect 22569 21505 22603 21539
rect 22753 21505 22787 21539
rect 23397 21505 23431 21539
rect 23673 21505 23707 21539
rect 3985 21437 4019 21471
rect 5365 21437 5399 21471
rect 5641 21437 5675 21471
rect 5733 21437 5767 21471
rect 5917 21437 5951 21471
rect 6469 21437 6503 21471
rect 6745 21437 6779 21471
rect 6837 21437 6871 21471
rect 6929 21437 6963 21471
rect 16313 21437 16347 21471
rect 17325 21437 17359 21471
rect 18061 21437 18095 21471
rect 18429 21437 18463 21471
rect 22017 21437 22051 21471
rect 22385 21437 22419 21471
rect 22477 21437 22511 21471
rect 23305 21437 23339 21471
rect 23765 21437 23799 21471
rect 3709 21369 3743 21403
rect 12449 21369 12483 21403
rect 15301 21369 15335 21403
rect 17509 21369 17543 21403
rect 18337 21369 18371 21403
rect 23029 21369 23063 21403
rect 1593 21301 1627 21335
rect 4537 21301 4571 21335
rect 9045 21301 9079 21335
rect 14749 21301 14783 21335
rect 14933 21301 14967 21335
rect 15669 21301 15703 21335
rect 15945 21301 15979 21335
rect 18153 21301 18187 21335
rect 18613 21301 18647 21335
rect 2881 21097 2915 21131
rect 5825 21097 5859 21131
rect 10793 21097 10827 21131
rect 15025 21097 15059 21131
rect 15945 21097 15979 21131
rect 17601 21097 17635 21131
rect 18521 21097 18555 21131
rect 19257 21097 19291 21131
rect 21557 21097 21591 21131
rect 22661 21097 22695 21131
rect 2789 21029 2823 21063
rect 6653 21029 6687 21063
rect 6745 21029 6779 21063
rect 15761 21029 15795 21063
rect 21281 21029 21315 21063
rect 22569 21029 22603 21063
rect 5457 20961 5491 20995
rect 9413 20961 9447 20995
rect 17325 20961 17359 20995
rect 17417 20961 17451 20995
rect 18337 20961 18371 20995
rect 18889 20961 18923 20995
rect 22017 20961 22051 20995
rect 1409 20893 1443 20927
rect 1676 20893 1710 20927
rect 3433 20893 3467 20927
rect 3801 20893 3835 20927
rect 5273 20893 5307 20927
rect 5365 20893 5399 20927
rect 5641 20893 5675 20927
rect 5733 20893 5767 20927
rect 5917 20893 5951 20927
rect 6561 20893 6595 20927
rect 6837 20893 6871 20927
rect 7389 20893 7423 20927
rect 7573 20893 7607 20927
rect 7849 20893 7883 20927
rect 8953 20893 8987 20927
rect 9137 20893 9171 20927
rect 18245 20893 18279 20927
rect 18705 20893 18739 20927
rect 18797 20893 18831 20927
rect 18981 20893 19015 20927
rect 19441 20893 19475 20927
rect 19533 20893 19567 20927
rect 20177 20893 20211 20927
rect 20269 20893 20303 20927
rect 20545 20893 20579 20927
rect 20637 20893 20671 20927
rect 20729 20893 20763 20927
rect 20913 20893 20947 20927
rect 21189 20893 21223 20927
rect 21373 20893 21407 20927
rect 21465 20893 21499 20927
rect 21649 20893 21683 20927
rect 22201 20893 22235 20927
rect 22845 20893 22879 20927
rect 23121 20893 23155 20927
rect 23213 20893 23247 20927
rect 23489 20893 23523 20927
rect 4068 20825 4102 20859
rect 6377 20825 6411 20859
rect 7757 20825 7791 20859
rect 9680 20825 9714 20859
rect 14841 20825 14875 20859
rect 15057 20825 15091 20859
rect 16129 20825 16163 20859
rect 19257 20825 19291 20859
rect 20361 20825 20395 20859
rect 22293 20825 22327 20859
rect 23029 20825 23063 20859
rect 23305 20825 23339 20859
rect 5181 20757 5215 20791
rect 5549 20757 5583 20791
rect 9045 20757 9079 20791
rect 15209 20757 15243 20791
rect 15929 20757 15963 20791
rect 16957 20757 16991 20791
rect 19993 20757 20027 20791
rect 21097 20757 21131 20791
rect 22385 20757 22419 20791
rect 23213 20757 23247 20791
rect 5273 20553 5307 20587
rect 9321 20553 9355 20587
rect 12909 20553 12943 20587
rect 20361 20553 20395 20587
rect 5641 20485 5675 20519
rect 6929 20485 6963 20519
rect 10793 20485 10827 20519
rect 20545 20485 20579 20519
rect 4629 20417 4663 20451
rect 5181 20417 5215 20451
rect 5825 20417 5859 20451
rect 8953 20417 8987 20451
rect 9965 20417 9999 20451
rect 10609 20417 10643 20451
rect 10701 20417 10735 20451
rect 10977 20417 11011 20451
rect 11529 20417 11563 20451
rect 11785 20417 11819 20451
rect 13737 20417 13771 20451
rect 13826 20417 13860 20451
rect 13921 20417 13955 20451
rect 14105 20417 14139 20451
rect 14565 20417 14599 20451
rect 16037 20417 16071 20451
rect 20269 20417 20303 20451
rect 3249 20349 3283 20383
rect 4537 20349 4571 20383
rect 9045 20349 9079 20383
rect 24317 20349 24351 20383
rect 6653 20281 6687 20315
rect 10977 20281 11011 20315
rect 20545 20281 20579 20315
rect 24041 20281 24075 20315
rect 2697 20213 2731 20247
rect 3893 20213 3927 20247
rect 5457 20213 5491 20247
rect 6469 20213 6503 20247
rect 13461 20213 13495 20247
rect 14381 20213 14415 20247
rect 15761 20213 15795 20247
rect 23857 20213 23891 20247
rect 11897 20009 11931 20043
rect 15209 20009 15243 20043
rect 15669 20009 15703 20043
rect 17693 20009 17727 20043
rect 18797 20009 18831 20043
rect 20729 20009 20763 20043
rect 22661 20009 22695 20043
rect 24041 20009 24075 20043
rect 24225 20009 24259 20043
rect 24501 20009 24535 20043
rect 3617 19941 3651 19975
rect 6377 19941 6411 19975
rect 6561 19941 6595 19975
rect 8033 19941 8067 19975
rect 8401 19941 8435 19975
rect 9045 19941 9079 19975
rect 20913 19941 20947 19975
rect 24961 19941 24995 19975
rect 8125 19873 8159 19907
rect 16221 19873 16255 19907
rect 18337 19873 18371 19907
rect 19257 19873 19291 19907
rect 19717 19873 19751 19907
rect 19993 19873 20027 19907
rect 21281 19873 21315 19907
rect 22201 19873 22235 19907
rect 1409 19805 1443 19839
rect 2237 19805 2271 19839
rect 6653 19805 6687 19839
rect 9229 19805 9263 19839
rect 9965 19805 9999 19839
rect 10149 19805 10183 19839
rect 10609 19805 10643 19839
rect 12541 19805 12575 19839
rect 14105 19805 14139 19839
rect 15945 19805 15979 19839
rect 16037 19805 16071 19839
rect 16313 19805 16347 19839
rect 18521 19805 18555 19839
rect 19625 19805 19659 19839
rect 19901 19805 19935 19839
rect 20085 19805 20119 19839
rect 20453 19805 20487 19839
rect 20821 19805 20855 19839
rect 21925 19805 21959 19839
rect 22569 19805 22603 19839
rect 22937 19805 22971 19839
rect 23213 19805 23247 19839
rect 23489 19805 23523 19839
rect 23765 19805 23799 19839
rect 24409 19805 24443 19839
rect 24777 19805 24811 19839
rect 2504 19737 2538 19771
rect 4261 19737 4295 19771
rect 6009 19737 6043 19771
rect 6101 19737 6135 19771
rect 6920 19737 6954 19771
rect 12808 19737 12842 19771
rect 14565 19737 14599 19771
rect 15193 19737 15227 19771
rect 15393 19737 15427 19771
rect 15637 19737 15671 19771
rect 15853 19737 15887 19771
rect 16580 19737 16614 19771
rect 18705 19737 18739 19771
rect 23305 19737 23339 19771
rect 23857 19737 23891 19771
rect 1593 19669 1627 19703
rect 8585 19669 8619 19703
rect 10057 19669 10091 19703
rect 13921 19669 13955 19703
rect 14289 19669 14323 19703
rect 14657 19669 14691 19703
rect 15025 19669 15059 19703
rect 15485 19669 15519 19703
rect 16221 19669 16255 19703
rect 17785 19669 17819 19703
rect 20545 19669 20579 19703
rect 21189 19669 21223 19703
rect 23673 19669 23707 19703
rect 24057 19669 24091 19703
rect 5181 19465 5215 19499
rect 7021 19465 7055 19499
rect 10793 19465 10827 19499
rect 12265 19465 12299 19499
rect 13829 19465 13863 19499
rect 15577 19465 15611 19499
rect 16681 19465 16715 19499
rect 19993 19465 20027 19499
rect 20821 19465 20855 19499
rect 23857 19465 23891 19499
rect 24409 19465 24443 19499
rect 5825 19397 5859 19431
rect 7849 19397 7883 19431
rect 8125 19397 8159 19431
rect 8462 19397 8496 19431
rect 10241 19397 10275 19431
rect 10977 19397 11011 19431
rect 14105 19397 14139 19431
rect 14315 19397 14349 19431
rect 14841 19397 14875 19431
rect 15301 19397 15335 19431
rect 16957 19397 16991 19431
rect 18613 19397 18647 19431
rect 22937 19397 22971 19431
rect 23153 19397 23187 19431
rect 1409 19329 1443 19363
rect 1676 19329 1710 19363
rect 3801 19329 3835 19363
rect 4068 19329 4102 19363
rect 5641 19329 5675 19363
rect 5917 19329 5951 19363
rect 6009 19329 6043 19363
rect 6377 19329 6411 19363
rect 6470 19329 6504 19363
rect 6653 19329 6687 19363
rect 6745 19329 6779 19363
rect 6842 19329 6876 19363
rect 7619 19329 7653 19363
rect 7757 19329 7791 19363
rect 7941 19329 7975 19363
rect 11805 19329 11839 19363
rect 12633 19329 12667 19363
rect 12909 19329 12943 19363
rect 13093 19329 13127 19363
rect 13185 19329 13219 19363
rect 13277 19329 13311 19363
rect 14013 19329 14047 19363
rect 14197 19329 14231 19363
rect 15025 19329 15059 19363
rect 15117 19329 15151 19363
rect 15209 19329 15243 19363
rect 15393 19329 15427 19363
rect 15485 19329 15519 19363
rect 15669 19329 15703 19363
rect 16865 19329 16899 19363
rect 17049 19329 17083 19363
rect 17167 19329 17201 19363
rect 17325 19329 17359 19363
rect 18521 19329 18555 19363
rect 18705 19329 18739 19363
rect 18981 19329 19015 19363
rect 19809 19329 19843 19363
rect 20085 19329 20119 19363
rect 20177 19329 20211 19363
rect 20361 19329 20395 19363
rect 20453 19329 20487 19363
rect 20637 19329 20671 19363
rect 20913 19329 20947 19363
rect 23765 19329 23799 19363
rect 24041 19329 24075 19363
rect 24317 19329 24351 19363
rect 25053 19329 25087 19363
rect 7481 19261 7515 19295
rect 8217 19261 8251 19295
rect 10701 19261 10735 19295
rect 11688 19261 11722 19295
rect 11897 19261 11931 19295
rect 12173 19261 12207 19295
rect 12725 19261 12759 19295
rect 14473 19261 14507 19295
rect 14841 19261 14875 19295
rect 24225 19261 24259 19295
rect 24961 19261 24995 19295
rect 2789 19193 2823 19227
rect 6193 19193 6227 19227
rect 10241 19193 10275 19227
rect 19625 19193 19659 19227
rect 24685 19193 24719 19227
rect 9597 19125 9631 19159
rect 11529 19125 11563 19159
rect 13553 19125 13587 19159
rect 18889 19125 18923 19159
rect 20269 19125 20303 19159
rect 23121 19125 23155 19159
rect 23305 19125 23339 19159
rect 9781 18921 9815 18955
rect 10425 18921 10459 18955
rect 11253 18921 11287 18955
rect 12357 18921 12391 18955
rect 13185 18921 13219 18955
rect 14841 18921 14875 18955
rect 21649 18921 21683 18955
rect 23029 18921 23063 18955
rect 10977 18853 11011 18887
rect 11897 18853 11931 18887
rect 3893 18785 3927 18819
rect 10241 18785 10275 18819
rect 11529 18785 11563 18819
rect 13001 18785 13035 18819
rect 5457 18717 5491 18751
rect 9229 18717 9263 18751
rect 9965 18717 9999 18751
rect 10057 18717 10091 18751
rect 10149 18717 10183 18751
rect 10606 18717 10640 18751
rect 11069 18717 11103 18751
rect 11621 18717 11655 18751
rect 12081 18717 12115 18751
rect 12173 18717 12207 18751
rect 13277 18717 13311 18751
rect 15301 18717 15335 18751
rect 17969 18717 18003 18751
rect 18061 18717 18095 18751
rect 18245 18717 18279 18751
rect 18337 18717 18371 18751
rect 18429 18717 18463 18751
rect 18613 18717 18647 18751
rect 18705 18717 18739 18751
rect 18889 18717 18923 18751
rect 21465 18717 21499 18751
rect 21741 18717 21775 18751
rect 4160 18649 4194 18683
rect 11161 18649 11195 18683
rect 12541 18649 12575 18683
rect 14657 18649 14691 18683
rect 14873 18649 14907 18683
rect 18521 18649 18555 18683
rect 20085 18649 20119 18683
rect 20269 18649 20303 18683
rect 22661 18649 22695 18683
rect 22845 18649 22879 18683
rect 5273 18581 5307 18615
rect 6745 18581 6779 18615
rect 9045 18581 9079 18615
rect 10609 18581 10643 18615
rect 11805 18581 11839 18615
rect 12725 18581 12759 18615
rect 15025 18581 15059 18615
rect 17785 18581 17819 18615
rect 18889 18581 18923 18615
rect 21281 18581 21315 18615
rect 4813 18377 4847 18411
rect 6545 18377 6579 18411
rect 9965 18377 9999 18411
rect 10333 18377 10367 18411
rect 19533 18377 19567 18411
rect 20269 18377 20303 18411
rect 24501 18377 24535 18411
rect 24685 18377 24719 18411
rect 6745 18309 6779 18343
rect 7021 18309 7055 18343
rect 9413 18309 9447 18343
rect 14105 18309 14139 18343
rect 14749 18309 14783 18343
rect 19073 18309 19107 18343
rect 20453 18309 20487 18343
rect 21649 18309 21683 18343
rect 23397 18309 23431 18343
rect 25145 18309 25179 18343
rect 2237 18241 2271 18275
rect 2504 18241 2538 18275
rect 3709 18241 3743 18275
rect 3893 18241 3927 18275
rect 4077 18241 4111 18275
rect 4169 18241 4203 18275
rect 4353 18241 4387 18275
rect 4997 18241 5031 18275
rect 5089 18241 5123 18275
rect 5181 18241 5215 18275
rect 5299 18241 5333 18275
rect 5549 18241 5583 18275
rect 6837 18241 6871 18275
rect 7113 18241 7147 18275
rect 7472 18241 7506 18275
rect 9597 18241 9631 18275
rect 9873 18241 9907 18275
rect 10057 18241 10091 18275
rect 10241 18241 10275 18275
rect 10425 18241 10459 18275
rect 11897 18241 11931 18275
rect 11989 18241 12023 18275
rect 12173 18241 12207 18275
rect 12275 18241 12309 18275
rect 16937 18241 16971 18275
rect 18889 18241 18923 18275
rect 19165 18241 19199 18275
rect 19257 18241 19291 18275
rect 20085 18241 20119 18275
rect 20177 18241 20211 18275
rect 22385 18241 22419 18275
rect 23581 18241 23615 18275
rect 23764 18241 23798 18275
rect 23857 18241 23891 18275
rect 24409 18241 24443 18275
rect 24593 18241 24627 18275
rect 24869 18241 24903 18275
rect 25421 18241 25455 18275
rect 25605 18241 25639 18275
rect 5457 18173 5491 18207
rect 7205 18173 7239 18207
rect 9229 18173 9263 18207
rect 9781 18173 9815 18207
rect 16681 18173 16715 18207
rect 18153 18173 18187 18207
rect 18705 18173 18739 18207
rect 19809 18173 19843 18207
rect 20821 18173 20855 18207
rect 23673 18173 23707 18207
rect 25053 18173 25087 18207
rect 6377 18105 6411 18139
rect 8585 18105 8619 18139
rect 25237 18105 25271 18139
rect 3617 18037 3651 18071
rect 4261 18037 4295 18071
rect 6561 18037 6595 18071
rect 6837 18037 6871 18071
rect 8677 18037 8711 18071
rect 11713 18037 11747 18071
rect 12633 18037 12667 18071
rect 16037 18037 16071 18071
rect 18061 18037 18095 18071
rect 19441 18037 19475 18071
rect 19993 18037 20027 18071
rect 20453 18037 20487 18071
rect 24041 18037 24075 18071
rect 25145 18037 25179 18071
rect 2789 17833 2823 17867
rect 5549 17833 5583 17867
rect 6101 17833 6135 17867
rect 7389 17833 7423 17867
rect 9689 17833 9723 17867
rect 10333 17833 10367 17867
rect 11161 17833 11195 17867
rect 11805 17833 11839 17867
rect 13001 17833 13035 17867
rect 13461 17833 13495 17867
rect 16773 17833 16807 17867
rect 18061 17833 18095 17867
rect 18337 17833 18371 17867
rect 20177 17833 20211 17867
rect 22845 17833 22879 17867
rect 23029 17833 23063 17867
rect 24409 17833 24443 17867
rect 24593 17833 24627 17867
rect 25237 17833 25271 17867
rect 4905 17765 4939 17799
rect 9413 17765 9447 17799
rect 10793 17765 10827 17799
rect 15485 17765 15519 17799
rect 6745 17697 6779 17731
rect 8033 17697 8067 17731
rect 9597 17697 9631 17731
rect 9781 17697 9815 17731
rect 9965 17697 9999 17731
rect 11069 17697 11103 17731
rect 15853 17697 15887 17731
rect 17417 17697 17451 17731
rect 18153 17697 18187 17731
rect 2973 17629 3007 17663
rect 3065 17629 3099 17663
rect 3433 17629 3467 17663
rect 4721 17629 4755 17663
rect 4905 17629 4939 17663
rect 6009 17629 6043 17663
rect 6193 17629 6227 17663
rect 6653 17629 6687 17663
rect 6837 17629 6871 17663
rect 7573 17629 7607 17663
rect 7665 17629 7699 17663
rect 9229 17629 9263 17663
rect 9413 17629 9447 17663
rect 9873 17629 9907 17663
rect 10241 17629 10275 17663
rect 10425 17629 10459 17663
rect 10638 17629 10672 17663
rect 11161 17629 11195 17663
rect 11989 17629 12023 17663
rect 12725 17629 12759 17663
rect 13185 17629 13219 17663
rect 13553 17629 13587 17663
rect 14105 17629 14139 17663
rect 14381 17629 14415 17663
rect 16129 17629 16163 17663
rect 16957 17629 16991 17663
rect 17049 17629 17083 17663
rect 17141 17629 17175 17663
rect 17259 17629 17293 17663
rect 17785 17629 17819 17663
rect 17877 17629 17911 17663
rect 17969 17629 18003 17663
rect 18245 17629 18279 17663
rect 18429 17629 18463 17663
rect 19901 17629 19935 17663
rect 20177 17629 20211 17663
rect 22661 17629 22695 17663
rect 22845 17629 22879 17663
rect 24961 17629 24995 17663
rect 25053 17629 25087 17663
rect 25513 17629 25547 17663
rect 3157 17561 3191 17595
rect 3295 17561 3329 17595
rect 5733 17561 5767 17595
rect 5917 17561 5951 17595
rect 7757 17561 7791 17595
rect 7875 17561 7909 17595
rect 11713 17561 11747 17595
rect 11897 17561 11931 17595
rect 20085 17561 20119 17595
rect 25421 17561 25455 17595
rect 10609 17493 10643 17527
rect 17601 17493 17635 17527
rect 24593 17493 24627 17527
rect 3985 17289 4019 17323
rect 4905 17289 4939 17323
rect 6745 17289 6779 17323
rect 10517 17289 10551 17323
rect 11529 17289 11563 17323
rect 14749 17289 14783 17323
rect 16405 17289 16439 17323
rect 17877 17289 17911 17323
rect 19349 17289 19383 17323
rect 21189 17289 21223 17323
rect 21833 17289 21867 17323
rect 22017 17289 22051 17323
rect 22937 17289 22971 17323
rect 23213 17289 23247 17323
rect 25053 17289 25087 17323
rect 25221 17289 25255 17323
rect 8033 17221 8067 17255
rect 8585 17221 8619 17255
rect 11897 17221 11931 17255
rect 15485 17221 15519 17255
rect 16681 17221 16715 17255
rect 18214 17221 18248 17255
rect 21557 17221 21591 17255
rect 23381 17221 23415 17255
rect 23581 17221 23615 17255
rect 25421 17221 25455 17255
rect 1676 17153 1710 17187
rect 3801 17153 3835 17187
rect 4077 17153 4111 17187
rect 4445 17153 4479 17187
rect 4721 17153 4755 17187
rect 4997 17153 5031 17187
rect 5089 17153 5123 17187
rect 5273 17153 5307 17187
rect 5549 17153 5583 17187
rect 5733 17153 5767 17187
rect 6377 17153 6411 17187
rect 7205 17153 7239 17187
rect 7297 17153 7331 17187
rect 7481 17153 7515 17187
rect 7573 17153 7607 17187
rect 7849 17153 7883 17187
rect 8125 17153 8159 17187
rect 8493 17153 8527 17187
rect 8677 17153 8711 17187
rect 10057 17153 10091 17187
rect 10149 17153 10183 17187
rect 11713 17153 11747 17187
rect 11805 17153 11839 17187
rect 13665 17153 13699 17187
rect 14933 17153 14967 17187
rect 15025 17153 15059 17187
rect 15117 17153 15151 17187
rect 15255 17153 15289 17187
rect 15761 17153 15795 17187
rect 15853 17153 15887 17187
rect 16037 17153 16071 17187
rect 16313 17153 16347 17187
rect 16497 17153 16531 17187
rect 16865 17153 16899 17187
rect 17325 17153 17359 17187
rect 17509 17153 17543 17187
rect 17601 17153 17635 17187
rect 17693 17153 17727 17187
rect 17969 17153 18003 17187
rect 20453 17153 20487 17187
rect 20611 17153 20645 17187
rect 20729 17153 20763 17187
rect 20821 17153 20855 17187
rect 20913 17153 20947 17187
rect 21189 17153 21223 17187
rect 21373 17153 21407 17187
rect 21465 17153 21499 17187
rect 21649 17153 21683 17187
rect 22014 17153 22048 17187
rect 22385 17153 22419 17187
rect 22477 17153 22511 17187
rect 22569 17153 22603 17187
rect 22937 17153 22971 17187
rect 24777 17153 24811 17187
rect 24961 17153 24995 17187
rect 25513 17153 25547 17187
rect 25697 17153 25731 17187
rect 25789 17153 25823 17187
rect 26065 17153 26099 17187
rect 1409 17085 1443 17119
rect 3433 17085 3467 17119
rect 4537 17085 4571 17119
rect 6469 17085 6503 17119
rect 10241 17085 10275 17119
rect 13921 17085 13955 17119
rect 15393 17085 15427 17119
rect 15485 17085 15519 17119
rect 17049 17085 17083 17119
rect 23121 17085 23155 17119
rect 2789 17017 2823 17051
rect 12081 17017 12115 17051
rect 21097 17017 21131 17051
rect 24869 17017 24903 17051
rect 25881 17017 25915 17051
rect 2881 16949 2915 16983
rect 3617 16949 3651 16983
rect 4445 16949 4479 16983
rect 5457 16949 5491 16983
rect 5641 16949 5675 16983
rect 6377 16949 6411 16983
rect 7021 16949 7055 16983
rect 7665 16949 7699 16983
rect 9965 16949 9999 16983
rect 10241 16949 10275 16983
rect 12541 16949 12575 16983
rect 15669 16949 15703 16983
rect 15853 16949 15887 16983
rect 23397 16949 23431 16983
rect 25237 16949 25271 16983
rect 25513 16949 25547 16983
rect 1961 16745 1995 16779
rect 6561 16745 6595 16779
rect 9597 16745 9631 16779
rect 11069 16745 11103 16779
rect 12173 16745 12207 16779
rect 18061 16745 18095 16779
rect 20085 16745 20119 16779
rect 20545 16745 20579 16779
rect 21005 16745 21039 16779
rect 21189 16745 21223 16779
rect 23397 16745 23431 16779
rect 2973 16677 3007 16711
rect 10425 16677 10459 16711
rect 12357 16677 12391 16711
rect 19901 16677 19935 16711
rect 21557 16677 21591 16711
rect 3341 16609 3375 16643
rect 6653 16609 6687 16643
rect 9045 16609 9079 16643
rect 9781 16609 9815 16643
rect 10241 16609 10275 16643
rect 11621 16609 11655 16643
rect 11989 16609 12023 16643
rect 14473 16609 14507 16643
rect 17233 16609 17267 16643
rect 17693 16609 17727 16643
rect 18521 16609 18555 16643
rect 18705 16609 18739 16643
rect 19671 16609 19705 16643
rect 20269 16609 20303 16643
rect 21281 16609 21315 16643
rect 21465 16609 21499 16643
rect 23213 16609 23247 16643
rect 23581 16609 23615 16643
rect 2145 16541 2179 16575
rect 2605 16541 2639 16575
rect 2789 16541 2823 16575
rect 2881 16541 2915 16575
rect 3157 16541 3191 16575
rect 3985 16541 4019 16575
rect 4077 16541 4111 16575
rect 4445 16541 4479 16575
rect 4629 16541 4663 16575
rect 5825 16541 5859 16575
rect 5917 16541 5951 16575
rect 6561 16541 6595 16575
rect 6837 16541 6871 16575
rect 8953 16541 8987 16575
rect 9137 16541 9171 16575
rect 9873 16541 9907 16575
rect 10609 16541 10643 16575
rect 11437 16541 11471 16575
rect 12173 16541 12207 16575
rect 12449 16541 12483 16575
rect 13001 16541 13035 16575
rect 14105 16541 14139 16575
rect 17325 16541 17359 16575
rect 19533 16541 19567 16575
rect 19809 16541 19843 16575
rect 19993 16541 20027 16575
rect 20361 16541 20395 16575
rect 21373 16541 21407 16575
rect 21649 16541 21683 16575
rect 21741 16541 21775 16575
rect 23121 16541 23155 16575
rect 23765 16541 23799 16575
rect 24041 16541 24075 16575
rect 2237 16473 2271 16507
rect 2329 16473 2363 16507
rect 2467 16473 2501 16507
rect 6193 16473 6227 16507
rect 6285 16473 6319 16507
rect 10149 16473 10183 16507
rect 10793 16473 10827 16507
rect 11253 16473 11287 16507
rect 11713 16473 11747 16507
rect 14740 16473 14774 16507
rect 20085 16473 20119 16507
rect 4261 16405 4295 16439
rect 4537 16405 4571 16439
rect 5641 16405 5675 16439
rect 6377 16405 6411 16439
rect 11345 16405 11379 16439
rect 12541 16405 12575 16439
rect 13645 16405 13679 16439
rect 14289 16405 14323 16439
rect 15853 16405 15887 16439
rect 18429 16405 18463 16439
rect 23949 16405 23983 16439
rect 9965 16201 9999 16235
rect 12541 16201 12575 16235
rect 13185 16201 13219 16235
rect 13921 16201 13955 16235
rect 15025 16201 15059 16235
rect 15209 16201 15243 16235
rect 10241 16133 10275 16167
rect 10333 16133 10367 16167
rect 10885 16133 10919 16167
rect 12173 16133 12207 16167
rect 12389 16133 12423 16167
rect 13435 16133 13469 16167
rect 15393 16133 15427 16167
rect 4261 16065 4295 16099
rect 4445 16065 4479 16099
rect 4905 16065 4939 16099
rect 5273 16065 5307 16099
rect 5825 16065 5859 16099
rect 6009 16065 6043 16099
rect 6193 16065 6227 16099
rect 7481 16065 7515 16099
rect 7665 16065 7699 16099
rect 7757 16065 7791 16099
rect 8033 16065 8067 16099
rect 8217 16065 8251 16099
rect 8677 16065 8711 16099
rect 8769 16065 8803 16099
rect 8953 16065 8987 16099
rect 10144 16065 10178 16099
rect 10461 16065 10495 16099
rect 10609 16065 10643 16099
rect 11805 16065 11839 16099
rect 11989 16065 12023 16099
rect 12817 16065 12851 16099
rect 13277 16065 13311 16099
rect 13553 16065 13587 16099
rect 13645 16065 13679 16099
rect 13737 16065 13771 16099
rect 14013 16065 14047 16099
rect 14197 16065 14231 16099
rect 15117 16065 15151 16099
rect 16865 16065 16899 16099
rect 16957 16065 16991 16099
rect 24777 16065 24811 16099
rect 24869 16065 24903 16099
rect 25053 16065 25087 16099
rect 25329 16065 25363 16099
rect 25513 16065 25547 16099
rect 8585 15997 8619 16031
rect 9137 15997 9171 16031
rect 12909 15997 12943 16031
rect 14105 15997 14139 16031
rect 14841 15997 14875 16031
rect 17141 15997 17175 16031
rect 25421 15997 25455 16031
rect 4077 15929 4111 15963
rect 10701 15929 10735 15963
rect 11253 15929 11287 15963
rect 6193 15861 6227 15895
rect 7297 15861 7331 15895
rect 8033 15861 8067 15895
rect 8309 15861 8343 15895
rect 8493 15861 8527 15895
rect 10885 15861 10919 15895
rect 11805 15861 11839 15895
rect 12357 15861 12391 15895
rect 17049 15861 17083 15895
rect 25237 15861 25271 15895
rect 8125 15657 8159 15691
rect 17141 15657 17175 15691
rect 20361 15657 20395 15691
rect 21925 15657 21959 15691
rect 24961 15657 24995 15691
rect 4169 15589 4203 15623
rect 15301 15589 15335 15623
rect 18981 15589 19015 15623
rect 19257 15589 19291 15623
rect 19901 15589 19935 15623
rect 25605 15589 25639 15623
rect 4353 15521 4387 15555
rect 6193 15521 6227 15555
rect 18521 15521 18555 15555
rect 19717 15521 19751 15555
rect 24685 15521 24719 15555
rect 26065 15521 26099 15555
rect 26341 15521 26375 15555
rect 1961 15453 1995 15487
rect 4445 15453 4479 15487
rect 4813 15453 4847 15487
rect 5089 15453 5123 15487
rect 6101 15453 6135 15487
rect 8033 15453 8067 15487
rect 8217 15453 8251 15487
rect 8309 15453 8343 15487
rect 8493 15453 8527 15487
rect 13093 15453 13127 15487
rect 15025 15453 15059 15487
rect 15301 15453 15335 15487
rect 15761 15453 15795 15487
rect 17417 15453 17451 15487
rect 17509 15453 17543 15487
rect 17601 15453 17635 15487
rect 17877 15453 17911 15487
rect 17969 15453 18003 15487
rect 18889 15453 18923 15487
rect 19073 15453 19107 15487
rect 19625 15453 19659 15487
rect 20177 15453 20211 15487
rect 20453 15453 20487 15487
rect 20820 15453 20854 15487
rect 20913 15453 20947 15487
rect 21281 15453 21315 15487
rect 21465 15453 21499 15487
rect 21557 15453 21591 15487
rect 21741 15453 21775 15487
rect 22477 15453 22511 15487
rect 23706 15453 23740 15487
rect 24133 15453 24167 15487
rect 24225 15453 24259 15487
rect 24593 15453 24627 15487
rect 25237 15453 25271 15487
rect 25973 15453 26007 15487
rect 26249 15453 26283 15487
rect 26433 15453 26467 15487
rect 2228 15385 2262 15419
rect 15117 15385 15151 15419
rect 16028 15385 16062 15419
rect 17233 15385 17267 15419
rect 17739 15385 17773 15419
rect 23489 15385 23523 15419
rect 3341 15317 3375 15351
rect 4629 15317 4663 15351
rect 4721 15317 4755 15351
rect 4997 15317 5031 15351
rect 5457 15317 5491 15351
rect 8401 15317 8435 15351
rect 13185 15317 13219 15351
rect 20545 15317 20579 15351
rect 23581 15317 23615 15351
rect 23765 15317 23799 15351
rect 25053 15317 25087 15351
rect 2513 15113 2547 15147
rect 4337 15113 4371 15147
rect 8953 15113 8987 15147
rect 11345 15113 11379 15147
rect 14105 15113 14139 15147
rect 14749 15113 14783 15147
rect 16773 15113 16807 15147
rect 17049 15113 17083 15147
rect 17785 15113 17819 15147
rect 19993 15113 20027 15147
rect 21005 15113 21039 15147
rect 22477 15113 22511 15147
rect 23857 15113 23891 15147
rect 24685 15113 24719 15147
rect 24869 15113 24903 15147
rect 25145 15113 25179 15147
rect 2237 15045 2271 15079
rect 4537 15045 4571 15079
rect 9045 15045 9079 15079
rect 11774 15045 11808 15079
rect 13461 15045 13495 15079
rect 13829 15045 13863 15079
rect 15117 15045 15151 15079
rect 15235 15045 15269 15079
rect 16221 15045 16255 15079
rect 17141 15045 17175 15079
rect 18061 15045 18095 15079
rect 20729 15045 20763 15079
rect 24961 15045 24995 15079
rect 1961 14977 1995 15011
rect 2145 14977 2179 15011
rect 2329 14977 2363 15011
rect 3249 14977 3283 15011
rect 3433 14977 3467 15011
rect 3893 14977 3927 15011
rect 4813 14977 4847 15011
rect 4997 14977 5031 15011
rect 5089 14977 5123 15011
rect 5733 14977 5767 15011
rect 5917 14977 5951 15011
rect 7205 14977 7239 15011
rect 7297 14977 7331 15011
rect 9413 14977 9447 15011
rect 9689 14977 9723 15011
rect 10241 14977 10275 15011
rect 10425 14977 10459 15011
rect 10609 14977 10643 15011
rect 10793 14977 10827 15011
rect 10977 14977 11011 15011
rect 11069 14977 11103 15011
rect 11161 14977 11195 15011
rect 13093 14977 13127 15011
rect 13277 14977 13311 15011
rect 13369 14977 13403 15011
rect 13599 14977 13633 15011
rect 14013 14977 14047 15011
rect 14197 14977 14231 15011
rect 14933 14977 14967 15011
rect 15025 14977 15059 15011
rect 15669 14977 15703 15011
rect 15945 14977 15979 15011
rect 16681 14977 16715 15011
rect 16865 14977 16899 15011
rect 17969 14977 18003 15011
rect 18153 14977 18187 15011
rect 18337 14977 18371 15011
rect 19809 14977 19843 15011
rect 20085 14977 20119 15011
rect 20637 14977 20671 15011
rect 20913 14977 20947 15011
rect 21189 14977 21223 15011
rect 21281 14977 21315 15011
rect 21649 14977 21683 15011
rect 21833 14977 21867 15011
rect 21925 14977 21959 15011
rect 22109 14977 22143 15011
rect 22201 14977 22235 15011
rect 22293 14977 22327 15011
rect 23765 14977 23799 15011
rect 23949 14977 23983 15011
rect 24688 14977 24722 15011
rect 25237 14977 25271 15011
rect 3065 14909 3099 14943
rect 3709 14909 3743 14943
rect 8861 14909 8895 14943
rect 9781 14909 9815 14943
rect 9873 14909 9907 14943
rect 9965 14909 9999 14943
rect 11529 14909 11563 14943
rect 13737 14909 13771 14943
rect 15393 14909 15427 14943
rect 15485 14909 15519 14943
rect 16221 14909 16255 14943
rect 24225 14909 24259 14943
rect 4169 14841 4203 14875
rect 8493 14841 8527 14875
rect 9505 14841 9539 14875
rect 19809 14841 19843 14875
rect 20913 14841 20947 14875
rect 24961 14841 24995 14875
rect 4077 14773 4111 14807
rect 4353 14773 4387 14807
rect 4629 14773 4663 14807
rect 5917 14773 5951 14807
rect 6101 14773 6135 14807
rect 6561 14773 6595 14807
rect 9321 14773 9355 14807
rect 12909 14773 12943 14807
rect 14381 14773 14415 14807
rect 15853 14773 15887 14807
rect 16037 14773 16071 14807
rect 21189 14773 21223 14807
rect 24317 14773 24351 14807
rect 1961 14569 1995 14603
rect 10241 14569 10275 14603
rect 13185 14569 13219 14603
rect 14841 14569 14875 14603
rect 18521 14569 18555 14603
rect 21649 14569 21683 14603
rect 22385 14569 22419 14603
rect 24501 14569 24535 14603
rect 10793 14501 10827 14535
rect 17877 14501 17911 14535
rect 23305 14501 23339 14535
rect 1685 14433 1719 14467
rect 4445 14433 4479 14467
rect 6745 14433 6779 14467
rect 7021 14433 7055 14467
rect 8401 14433 8435 14467
rect 8493 14433 8527 14467
rect 8677 14433 8711 14467
rect 23489 14433 23523 14467
rect 1593 14365 1627 14399
rect 2053 14365 2087 14399
rect 2237 14365 2271 14399
rect 3617 14365 3651 14399
rect 3985 14365 4019 14399
rect 4077 14365 4111 14399
rect 4353 14365 4387 14399
rect 6653 14365 6687 14399
rect 8585 14365 8619 14399
rect 9505 14365 9539 14399
rect 9689 14365 9723 14399
rect 10517 14365 10551 14399
rect 10609 14365 10643 14399
rect 10793 14365 10827 14399
rect 12725 14365 12759 14399
rect 12817 14365 12851 14399
rect 13001 14365 13035 14399
rect 13277 14365 13311 14399
rect 15025 14365 15059 14399
rect 15209 14365 15243 14399
rect 16221 14365 16255 14399
rect 16313 14365 16347 14399
rect 18061 14365 18095 14399
rect 18337 14365 18371 14399
rect 18429 14365 18463 14399
rect 18613 14365 18647 14399
rect 21741 14365 21775 14399
rect 21833 14365 21867 14399
rect 22293 14365 22327 14399
rect 22477 14365 22511 14399
rect 24409 14365 24443 14399
rect 24593 14365 24627 14399
rect 26617 14365 26651 14399
rect 26709 14365 26743 14399
rect 10057 14297 10091 14331
rect 10257 14297 10291 14331
rect 23029 14297 23063 14331
rect 2145 14229 2179 14263
rect 2973 14229 3007 14263
rect 3801 14229 3835 14263
rect 8217 14229 8251 14263
rect 9505 14229 9539 14263
rect 10425 14229 10459 14263
rect 13921 14229 13955 14263
rect 16037 14229 16071 14263
rect 16681 14229 16715 14263
rect 18245 14229 18279 14263
rect 21465 14229 21499 14263
rect 26065 14229 26099 14263
rect 1586 14025 1620 14059
rect 2329 14025 2363 14059
rect 3985 14025 4019 14059
rect 4997 14025 5031 14059
rect 6377 14025 6411 14059
rect 7757 14025 7791 14059
rect 11897 14025 11931 14059
rect 16155 14025 16189 14059
rect 17969 14025 18003 14059
rect 19625 14025 19659 14059
rect 21373 14025 21407 14059
rect 22569 14025 22603 14059
rect 26249 14025 26283 14059
rect 26709 14025 26743 14059
rect 2053 13957 2087 13991
rect 2666 13957 2700 13991
rect 4813 13957 4847 13991
rect 7021 13957 7055 13991
rect 8185 13957 8219 13991
rect 8401 13957 8435 13991
rect 13308 13957 13342 13991
rect 13645 13957 13679 13991
rect 14013 13957 14047 13991
rect 14131 13957 14165 13991
rect 15945 13957 15979 13991
rect 19717 13957 19751 13991
rect 22937 13957 22971 13991
rect 23213 13957 23247 13991
rect 25145 13957 25179 13991
rect 19441 13923 19475 13957
rect 1409 13889 1443 13923
rect 1501 13889 1535 13923
rect 1685 13889 1719 13923
rect 1777 13889 1811 13923
rect 1961 13889 1995 13923
rect 2145 13889 2179 13923
rect 4260 13889 4294 13923
rect 4353 13889 4387 13923
rect 4445 13889 4479 13923
rect 7665 13889 7699 13923
rect 7941 13889 7975 13923
rect 10057 13889 10091 13923
rect 10333 13889 10367 13923
rect 10517 13889 10551 13923
rect 11989 13889 12023 13923
rect 13553 13889 13587 13923
rect 13829 13889 13863 13923
rect 13921 13889 13955 13923
rect 14289 13889 14323 13923
rect 14565 13889 14599 13923
rect 14657 13889 14691 13923
rect 17233 13889 17267 13923
rect 17509 13889 17543 13923
rect 17601 13889 17635 13923
rect 17693 13889 17727 13923
rect 17877 13889 17911 13923
rect 17969 13889 18003 13923
rect 18061 13889 18095 13923
rect 18245 13889 18279 13923
rect 19073 13889 19107 13923
rect 19165 13889 19199 13923
rect 19533 13889 19567 13923
rect 19793 13879 19827 13913
rect 20085 13889 20119 13923
rect 20369 13889 20403 13923
rect 21189 13889 21223 13923
rect 21465 13889 21499 13923
rect 22753 13889 22787 13923
rect 23029 13889 23063 13923
rect 23121 13889 23155 13923
rect 23397 13889 23431 13923
rect 25053 13889 25087 13923
rect 25237 13889 25271 13923
rect 26065 13889 26099 13923
rect 26525 13889 26559 13923
rect 2421 13821 2455 13855
rect 5365 13821 5399 13855
rect 6101 13821 6135 13855
rect 6699 13821 6733 13855
rect 6837 13821 6871 13855
rect 9781 13821 9815 13855
rect 19257 13821 19291 13855
rect 25605 13821 25639 13855
rect 25973 13821 26007 13855
rect 26341 13821 26375 13855
rect 12173 13753 12207 13787
rect 16957 13753 16991 13787
rect 19993 13753 20027 13787
rect 20269 13753 20303 13787
rect 23121 13753 23155 13787
rect 3801 13685 3835 13719
rect 4813 13685 4847 13719
rect 7941 13685 7975 13719
rect 8033 13685 8067 13719
rect 8217 13685 8251 13719
rect 9505 13685 9539 13719
rect 9965 13685 9999 13719
rect 10333 13685 10367 13719
rect 14381 13685 14415 13719
rect 16129 13685 16163 13719
rect 16313 13685 16347 13719
rect 17417 13685 17451 13719
rect 17877 13685 17911 13719
rect 19441 13685 19475 13719
rect 21005 13685 21039 13719
rect 2053 13481 2087 13515
rect 4169 13481 4203 13515
rect 8125 13481 8159 13515
rect 8217 13481 8251 13515
rect 11069 13481 11103 13515
rect 14197 13481 14231 13515
rect 14289 13481 14323 13515
rect 19809 13481 19843 13515
rect 21005 13481 21039 13515
rect 21097 13481 21131 13515
rect 22937 13481 22971 13515
rect 24593 13481 24627 13515
rect 25697 13481 25731 13515
rect 1869 13413 1903 13447
rect 7205 13413 7239 13447
rect 8309 13413 8343 13447
rect 20085 13413 20119 13447
rect 24409 13413 24443 13447
rect 10885 13345 10919 13379
rect 11345 13345 11379 13379
rect 14105 13345 14139 13379
rect 15209 13345 15243 13379
rect 16129 13345 16163 13379
rect 19257 13345 19291 13379
rect 20269 13345 20303 13379
rect 20361 13345 20395 13379
rect 20729 13345 20763 13379
rect 21189 13345 21223 13379
rect 25881 13345 25915 13379
rect 25973 13345 26007 13379
rect 3985 13277 4019 13311
rect 5456 13277 5490 13311
rect 5549 13277 5583 13311
rect 7297 13277 7331 13311
rect 7573 13277 7607 13311
rect 7757 13277 7791 13311
rect 8401 13277 8435 13311
rect 8585 13277 8619 13311
rect 8953 13277 8987 13311
rect 9137 13277 9171 13311
rect 10149 13277 10183 13311
rect 10333 13277 10367 13311
rect 11161 13277 11195 13311
rect 11437 13277 11471 13311
rect 14381 13277 14415 13311
rect 14749 13277 14783 13311
rect 14933 13277 14967 13311
rect 15301 13277 15335 13311
rect 15485 13277 15519 13311
rect 16313 13277 16347 13311
rect 19625 13277 19659 13311
rect 20453 13277 20487 13311
rect 20545 13277 20579 13311
rect 21281 13277 21315 13311
rect 21465 13277 21499 13311
rect 21741 13277 21775 13311
rect 24593 13277 24627 13311
rect 24685 13277 24719 13311
rect 26065 13277 26099 13311
rect 26157 13277 26191 13311
rect 2021 13209 2055 13243
rect 2237 13209 2271 13243
rect 3801 13209 3835 13243
rect 7021 13209 7055 13243
rect 14841 13209 14875 13243
rect 15071 13209 15105 13243
rect 15393 13209 15427 13243
rect 21557 13209 21591 13243
rect 23121 13209 23155 13243
rect 25053 13209 25087 13243
rect 5181 13141 5215 13175
rect 7297 13141 7331 13175
rect 7665 13141 7699 13175
rect 7849 13141 7883 13175
rect 9045 13141 9079 13175
rect 10149 13141 10183 13175
rect 10885 13141 10919 13175
rect 11805 13141 11839 13175
rect 14565 13141 14599 13175
rect 16497 13141 16531 13175
rect 19441 13141 19475 13175
rect 21925 13141 21959 13175
rect 22753 13141 22787 13175
rect 22921 13141 22955 13175
rect 14841 12937 14875 12971
rect 16681 12937 16715 12971
rect 18337 12937 18371 12971
rect 20453 12937 20487 12971
rect 26157 12937 26191 12971
rect 10977 12869 11011 12903
rect 13461 12869 13495 12903
rect 14105 12869 14139 12903
rect 15209 12869 15243 12903
rect 15577 12869 15611 12903
rect 15669 12869 15703 12903
rect 16497 12869 16531 12903
rect 18797 12869 18831 12903
rect 23949 12869 23983 12903
rect 24041 12869 24075 12903
rect 24133 12869 24167 12903
rect 25973 12869 26007 12903
rect 26617 12869 26651 12903
rect 3709 12801 3743 12835
rect 3801 12801 3835 12835
rect 3985 12801 4019 12835
rect 7021 12801 7055 12835
rect 8125 12801 8159 12835
rect 8401 12801 8435 12835
rect 9873 12801 9907 12835
rect 10057 12801 10091 12835
rect 10149 12801 10183 12835
rect 10333 12801 10367 12835
rect 10425 12801 10459 12835
rect 10701 12801 10735 12835
rect 11161 12801 11195 12835
rect 13369 12801 13403 12835
rect 13553 12801 13587 12835
rect 13737 12801 13771 12835
rect 15025 12801 15059 12835
rect 15485 12801 15519 12835
rect 15853 12801 15887 12835
rect 16221 12801 16255 12835
rect 16313 12801 16347 12835
rect 16865 12801 16899 12835
rect 16957 12801 16991 12835
rect 17233 12801 17267 12835
rect 18429 12801 18463 12835
rect 18613 12801 18647 12835
rect 18889 12801 18923 12835
rect 19165 12801 19199 12835
rect 20361 12801 20395 12835
rect 20729 12801 20763 12835
rect 23673 12801 23707 12835
rect 23765 12801 23799 12835
rect 24409 12801 24443 12835
rect 25053 12801 25087 12835
rect 25604 12801 25638 12835
rect 25697 12801 25731 12835
rect 25789 12801 25823 12835
rect 26433 12801 26467 12835
rect 3893 12733 3927 12767
rect 6377 12733 6411 12767
rect 6929 12733 6963 12767
rect 8309 12733 8343 12767
rect 10517 12733 10551 12767
rect 14657 12733 14691 12767
rect 16497 12733 16531 12767
rect 17325 12733 17359 12767
rect 17877 12733 17911 12767
rect 17969 12733 18003 12767
rect 19349 12733 19383 12767
rect 20545 12733 20579 12767
rect 23949 12733 23983 12767
rect 24593 12733 24627 12767
rect 24961 12733 24995 12767
rect 25329 12733 25363 12767
rect 26249 12733 26283 12767
rect 17693 12665 17727 12699
rect 18981 12665 19015 12699
rect 3525 12597 3559 12631
rect 7941 12597 7975 12631
rect 8125 12597 8159 12631
rect 10885 12597 10919 12631
rect 11253 12597 11287 12631
rect 13185 12597 13219 12631
rect 15301 12597 15335 12631
rect 20729 12597 20763 12631
rect 24777 12597 24811 12631
rect 4261 12393 4295 12427
rect 7297 12393 7331 12427
rect 8217 12393 8251 12427
rect 9413 12393 9447 12427
rect 16865 12393 16899 12427
rect 17601 12393 17635 12427
rect 19625 12393 19659 12427
rect 20361 12393 20395 12427
rect 21649 12393 21683 12427
rect 25697 12393 25731 12427
rect 9229 12325 9263 12359
rect 9965 12325 9999 12359
rect 22845 12325 22879 12359
rect 3065 12257 3099 12291
rect 5273 12257 5307 12291
rect 5733 12257 5767 12291
rect 7665 12257 7699 12291
rect 7757 12257 7791 12291
rect 15485 12257 15519 12291
rect 20085 12257 20119 12291
rect 20545 12257 20579 12291
rect 22017 12257 22051 12291
rect 22477 12257 22511 12291
rect 22753 12257 22787 12291
rect 25053 12257 25087 12291
rect 25237 12257 25271 12291
rect 1961 12189 1995 12223
rect 2145 12189 2179 12223
rect 2283 12189 2317 12223
rect 2421 12189 2455 12223
rect 2697 12189 2731 12223
rect 2881 12189 2915 12223
rect 2973 12189 3007 12223
rect 3157 12189 3191 12223
rect 3801 12189 3835 12223
rect 3985 12189 4019 12223
rect 4537 12189 4571 12223
rect 5365 12189 5399 12223
rect 5825 12189 5859 12223
rect 6653 12189 6687 12223
rect 6837 12189 6871 12223
rect 7021 12189 7055 12223
rect 7113 12189 7147 12223
rect 7389 12189 7423 12223
rect 7573 12189 7607 12223
rect 7941 12189 7975 12223
rect 8401 12189 8435 12223
rect 8493 12189 8527 12223
rect 8677 12189 8711 12223
rect 8769 12189 8803 12223
rect 9689 12189 9723 12223
rect 9781 12189 9815 12223
rect 9965 12189 9999 12223
rect 11621 12189 11655 12223
rect 11805 12189 11839 12223
rect 11989 12189 12023 12223
rect 12173 12189 12207 12223
rect 12449 12189 12483 12223
rect 12633 12189 12667 12223
rect 15741 12189 15775 12223
rect 17601 12189 17635 12223
rect 17785 12189 17819 12223
rect 17877 12189 17911 12223
rect 19993 12189 20027 12223
rect 20637 12189 20671 12223
rect 21925 12189 21959 12223
rect 22385 12189 22419 12223
rect 23029 12189 23063 12223
rect 23213 12189 23247 12223
rect 23397 12189 23431 12223
rect 25513 12189 25547 12223
rect 25881 12189 25915 12223
rect 2053 12121 2087 12155
rect 4077 12121 4111 12155
rect 4282 12121 4316 12155
rect 9397 12121 9431 12155
rect 9597 12121 9631 12155
rect 23121 12121 23155 12155
rect 1777 12053 1811 12087
rect 2513 12053 2547 12087
rect 3893 12053 3927 12087
rect 4445 12053 4479 12087
rect 4813 12053 4847 12087
rect 6745 12053 6779 12087
rect 8125 12053 8159 12087
rect 11713 12053 11747 12087
rect 12357 12053 12391 12087
rect 12541 12053 12575 12087
rect 25421 12053 25455 12087
rect 2789 11849 2823 11883
rect 10701 11849 10735 11883
rect 14657 11849 14691 11883
rect 18981 11849 19015 11883
rect 24149 11849 24183 11883
rect 24317 11849 24351 11883
rect 24777 11849 24811 11883
rect 3801 11781 3835 11815
rect 13522 11781 13556 11815
rect 18797 11781 18831 11815
rect 23765 11781 23799 11815
rect 23949 11781 23983 11815
rect 25421 11781 25455 11815
rect 1409 11713 1443 11747
rect 1676 11713 1710 11747
rect 3157 11713 3191 11747
rect 3709 11713 3743 11747
rect 3893 11713 3927 11747
rect 5089 11713 5123 11747
rect 5273 11713 5307 11747
rect 5549 11713 5583 11747
rect 5733 11713 5767 11747
rect 6561 11713 6595 11747
rect 6929 11713 6963 11747
rect 7205 11713 7239 11747
rect 7849 11713 7883 11747
rect 8953 11713 8987 11747
rect 9137 11713 9171 11747
rect 10241 11713 10275 11747
rect 10333 11713 10367 11747
rect 10517 11713 10551 11747
rect 11621 11713 11655 11747
rect 11805 11713 11839 11747
rect 12173 11713 12207 11747
rect 12449 11713 12483 11747
rect 12633 11713 12667 11747
rect 13277 11713 13311 11747
rect 18613 11713 18647 11747
rect 20821 11713 20855 11747
rect 23489 11713 23523 11747
rect 24409 11713 24443 11747
rect 24593 11713 24627 11747
rect 26157 11713 26191 11747
rect 26249 11713 26283 11747
rect 26985 11713 27019 11747
rect 27169 11713 27203 11747
rect 27261 11713 27295 11747
rect 3249 11645 3283 11679
rect 4721 11645 4755 11679
rect 7113 11645 7147 11679
rect 7573 11645 7607 11679
rect 11897 11645 11931 11679
rect 11989 11645 12023 11679
rect 20913 11645 20947 11679
rect 21189 11645 21223 11679
rect 23305 11645 23339 11679
rect 23857 11645 23891 11679
rect 26065 11645 26099 11679
rect 26341 11645 26375 11679
rect 3525 11577 3559 11611
rect 25697 11577 25731 11611
rect 25881 11577 25915 11611
rect 6101 11509 6135 11543
rect 9137 11509 9171 11543
rect 12357 11509 12391 11543
rect 12449 11509 12483 11543
rect 24133 11509 24167 11543
rect 26525 11509 26559 11543
rect 4813 11305 4847 11339
rect 8309 11305 8343 11339
rect 9137 11305 9171 11339
rect 10885 11305 10919 11339
rect 19257 11305 19291 11339
rect 22109 11305 22143 11339
rect 24593 11305 24627 11339
rect 26157 11305 26191 11339
rect 11345 11237 11379 11271
rect 14841 11237 14875 11271
rect 7389 11169 7423 11203
rect 7757 11169 7791 11203
rect 8125 11169 8159 11203
rect 9045 11169 9079 11203
rect 10701 11169 10735 11203
rect 13001 11169 13035 11203
rect 14565 11169 14599 11203
rect 16037 11169 16071 11203
rect 26065 11169 26099 11203
rect 26249 11169 26283 11203
rect 4721 11101 4755 11135
rect 4905 11101 4939 11135
rect 5089 11101 5123 11135
rect 5549 11101 5583 11135
rect 5733 11101 5767 11135
rect 7849 11101 7883 11135
rect 8401 11101 8435 11135
rect 8953 11101 8987 11135
rect 9965 11101 9999 11135
rect 10057 11101 10091 11135
rect 10241 11101 10275 11135
rect 10333 11101 10367 11135
rect 10609 11101 10643 11135
rect 11069 11101 11103 11135
rect 11345 11101 11379 11135
rect 12541 11101 12575 11135
rect 12725 11101 12759 11135
rect 13093 11101 13127 11135
rect 14473 11101 14507 11135
rect 15025 11101 15059 11135
rect 17233 11101 17267 11135
rect 17417 11101 17451 11135
rect 17764 11101 17798 11135
rect 18061 11101 18095 11135
rect 18245 11101 18279 11135
rect 19257 11101 19291 11135
rect 19441 11101 19475 11135
rect 22385 11101 22419 11135
rect 24501 11101 24535 11135
rect 24685 11101 24719 11135
rect 25973 11101 26007 11135
rect 5273 11033 5307 11067
rect 5641 11033 5675 11067
rect 8033 11033 8067 11067
rect 9781 11033 9815 11067
rect 19073 11033 19107 11067
rect 22109 11033 22143 11067
rect 5457 10965 5491 10999
rect 8125 10965 8159 10999
rect 9321 10965 9355 10999
rect 11161 10965 11195 10999
rect 12633 10965 12667 10999
rect 13921 10965 13955 10999
rect 17693 10965 17727 10999
rect 19625 10965 19659 10999
rect 22293 10965 22327 10999
rect 12909 10761 12943 10795
rect 18153 10761 18187 10795
rect 20653 10761 20687 10795
rect 20821 10761 20855 10795
rect 22201 10761 22235 10795
rect 9413 10693 9447 10727
rect 13093 10693 13127 10727
rect 17233 10693 17267 10727
rect 17811 10693 17845 10727
rect 17985 10693 18019 10727
rect 19993 10693 20027 10727
rect 20193 10693 20227 10727
rect 20453 10693 20487 10727
rect 22937 10693 22971 10727
rect 25697 10693 25731 10727
rect 4537 10625 4571 10659
rect 4629 10625 4663 10659
rect 4905 10625 4939 10659
rect 5089 10625 5123 10659
rect 6653 10625 6687 10659
rect 7665 10625 7699 10659
rect 9137 10625 9171 10659
rect 9321 10625 9355 10659
rect 9505 10625 9539 10659
rect 12357 10625 12391 10659
rect 12449 10625 12483 10659
rect 12633 10625 12667 10659
rect 12725 10625 12759 10659
rect 12817 10625 12851 10659
rect 16129 10625 16163 10659
rect 16313 10625 16347 10659
rect 16865 10625 16899 10659
rect 17049 10625 17083 10659
rect 17325 10625 17359 10659
rect 17693 10625 17727 10659
rect 19625 10625 19659 10659
rect 20913 10625 20947 10659
rect 21005 10625 21039 10659
rect 22017 10625 22051 10659
rect 22293 10625 22327 10659
rect 22477 10625 22511 10659
rect 22753 10625 22787 10659
rect 24317 10625 24351 10659
rect 24501 10625 24535 10659
rect 24685 10625 24719 10659
rect 3341 10557 3375 10591
rect 4169 10557 4203 10591
rect 4261 10557 4295 10591
rect 4445 10557 4479 10591
rect 4721 10557 4755 10591
rect 6561 10557 6595 10591
rect 7389 10557 7423 10591
rect 19441 10557 19475 10591
rect 21189 10557 21223 10591
rect 21833 10557 21867 10591
rect 22661 10557 22695 10591
rect 24409 10557 24443 10591
rect 4997 10489 5031 10523
rect 13093 10489 13127 10523
rect 16129 10489 16163 10523
rect 21097 10489 21131 10523
rect 22569 10489 22603 10523
rect 7757 10421 7791 10455
rect 9689 10421 9723 10455
rect 12173 10421 12207 10455
rect 17929 10421 17963 10455
rect 19809 10421 19843 10455
rect 20177 10421 20211 10455
rect 20361 10421 20395 10455
rect 20637 10421 20671 10455
rect 6285 10217 6319 10251
rect 11897 10217 11931 10251
rect 15025 10217 15059 10251
rect 15485 10217 15519 10251
rect 16037 10217 16071 10251
rect 16773 10217 16807 10251
rect 16865 10217 16899 10251
rect 21373 10217 21407 10251
rect 21833 10217 21867 10251
rect 22569 10217 22603 10251
rect 25973 10217 26007 10251
rect 26341 10217 26375 10251
rect 26433 10217 26467 10251
rect 17509 10149 17543 10183
rect 18521 10149 18555 10183
rect 20959 10149 20993 10183
rect 21189 10149 21223 10183
rect 23857 10149 23891 10183
rect 9321 10081 9355 10115
rect 15577 10081 15611 10115
rect 16129 10081 16163 10115
rect 18061 10081 18095 10115
rect 19993 10081 20027 10115
rect 21465 10081 21499 10115
rect 23581 10081 23615 10115
rect 5457 10013 5491 10047
rect 5641 10013 5675 10047
rect 5733 10013 5767 10047
rect 6469 10013 6503 10047
rect 6837 10013 6871 10047
rect 8033 10013 8067 10047
rect 8217 10013 8251 10047
rect 9229 10013 9263 10047
rect 10425 10013 10459 10047
rect 10793 10013 10827 10047
rect 14289 10013 14323 10047
rect 14565 10013 14599 10047
rect 15209 10013 15243 10047
rect 15393 10013 15427 10047
rect 15761 10013 15795 10047
rect 16037 10013 16071 10047
rect 16589 10013 16623 10047
rect 16773 10013 16807 10047
rect 17049 10013 17083 10047
rect 17141 10013 17175 10047
rect 17325 10013 17359 10047
rect 17417 10013 17451 10047
rect 17785 10013 17819 10047
rect 18153 10013 18187 10047
rect 19717 10013 19751 10047
rect 20177 10013 20211 10047
rect 20361 10013 20395 10047
rect 20821 10013 20855 10047
rect 21097 10013 21131 10047
rect 21281 10013 21315 10047
rect 21649 10013 21683 10047
rect 21932 10013 21966 10047
rect 22018 10013 22052 10047
rect 22201 10013 22235 10047
rect 22293 10013 22327 10047
rect 22390 10013 22424 10047
rect 23489 10013 23523 10047
rect 23949 10013 23983 10047
rect 24133 10013 24167 10047
rect 25513 10013 25547 10047
rect 25789 10013 25823 10047
rect 26065 10013 26099 10047
rect 26341 10013 26375 10047
rect 26617 10013 26651 10047
rect 26709 10013 26743 10047
rect 6561 9945 6595 9979
rect 6653 9945 6687 9979
rect 14749 9945 14783 9979
rect 15301 9945 15335 9979
rect 15485 9945 15519 9979
rect 17509 9945 17543 9979
rect 19809 9945 19843 9979
rect 21373 9945 21407 9979
rect 26433 9945 26467 9979
rect 5273 9877 5307 9911
rect 5825 9877 5859 9911
rect 7849 9877 7883 9911
rect 10057 9877 10091 9911
rect 14105 9877 14139 9911
rect 14473 9877 14507 9911
rect 15945 9877 15979 9911
rect 16405 9877 16439 9911
rect 17693 9877 17727 9911
rect 24041 9877 24075 9911
rect 25605 9877 25639 9911
rect 26157 9877 26191 9911
rect 9321 9673 9355 9707
rect 23489 9673 23523 9707
rect 3601 9605 3635 9639
rect 3801 9605 3835 9639
rect 6745 9605 6779 9639
rect 7481 9605 7515 9639
rect 8769 9605 8803 9639
rect 3893 9537 3927 9571
rect 4077 9537 4111 9571
rect 4169 9537 4203 9571
rect 4445 9537 4479 9571
rect 5181 9537 5215 9571
rect 5457 9537 5491 9571
rect 5651 9537 5685 9571
rect 6377 9537 6411 9571
rect 6837 9537 6871 9571
rect 7205 9537 7239 9571
rect 7297 9537 7331 9571
rect 7941 9537 7975 9571
rect 9321 9537 9355 9571
rect 11713 9537 11747 9571
rect 12817 9537 12851 9571
rect 13001 9537 13035 9571
rect 14841 9537 14875 9571
rect 15485 9537 15519 9571
rect 17049 9537 17083 9571
rect 17325 9537 17359 9571
rect 19533 9537 19567 9571
rect 19625 9537 19659 9571
rect 19809 9537 19843 9571
rect 23673 9537 23707 9571
rect 23765 9537 23799 9571
rect 23949 9537 23983 9571
rect 24041 9537 24075 9571
rect 4629 9469 4663 9503
rect 4721 9469 4755 9503
rect 4813 9469 4847 9503
rect 4997 9469 5031 9503
rect 5089 9469 5123 9503
rect 5273 9469 5307 9503
rect 7757 9469 7791 9503
rect 8585 9469 8619 9503
rect 9413 9469 9447 9503
rect 11805 9469 11839 9503
rect 14473 9469 14507 9503
rect 15117 9469 15151 9503
rect 15393 9469 15427 9503
rect 17141 9469 17175 9503
rect 19717 9469 19751 9503
rect 7481 9401 7515 9435
rect 12081 9401 12115 9435
rect 14565 9401 14599 9435
rect 17233 9401 17267 9435
rect 3433 9333 3467 9367
rect 3617 9333 3651 9367
rect 3893 9333 3927 9367
rect 4261 9333 4295 9367
rect 5549 9333 5583 9367
rect 6561 9333 6595 9367
rect 16865 9333 16899 9367
rect 19993 9333 20027 9367
rect 8125 9129 8159 9163
rect 12817 9129 12851 9163
rect 16221 9129 16255 9163
rect 19717 9129 19751 9163
rect 21833 9129 21867 9163
rect 11345 9061 11379 9095
rect 19901 9061 19935 9095
rect 21557 9061 21591 9095
rect 22201 9061 22235 9095
rect 5365 8993 5399 9027
rect 5825 8993 5859 9027
rect 6561 8993 6595 9027
rect 10057 8993 10091 9027
rect 13645 8993 13679 9027
rect 15301 8993 15335 9027
rect 16865 8993 16899 9027
rect 17601 8993 17635 9027
rect 20177 8993 20211 9027
rect 24777 8993 24811 9027
rect 3801 8925 3835 8959
rect 3985 8925 4019 8959
rect 5273 8925 5307 8959
rect 5733 8925 5767 8959
rect 5917 8925 5951 8959
rect 6745 8925 6779 8959
rect 7941 8925 7975 8959
rect 8125 8925 8159 8959
rect 11069 8925 11103 8959
rect 11345 8925 11379 8959
rect 12357 8925 12391 8959
rect 12633 8925 12667 8959
rect 13553 8925 13587 8959
rect 13921 8925 13955 8959
rect 14289 8925 14323 8959
rect 14473 8925 14507 8959
rect 16773 8925 16807 8959
rect 17693 8925 17727 8959
rect 17877 8925 17911 8959
rect 17969 8925 18003 8959
rect 18153 8925 18187 8959
rect 20269 8925 20303 8959
rect 21557 8925 21591 8959
rect 21741 8925 21775 8959
rect 21833 8925 21867 8959
rect 22017 8925 22051 8959
rect 22385 8925 22419 8959
rect 22845 8925 22879 8959
rect 24041 8925 24075 8959
rect 24225 8925 24259 8959
rect 24409 8925 24443 8959
rect 24685 8925 24719 8959
rect 24961 8925 24995 8959
rect 25145 8925 25179 8959
rect 25513 8925 25547 8959
rect 25697 8925 25731 8959
rect 25881 8925 25915 8959
rect 10885 8857 10919 8891
rect 13829 8857 13863 8891
rect 16037 8857 16071 8891
rect 16237 8857 16271 8891
rect 19533 8857 19567 8891
rect 21097 8857 21131 8891
rect 25605 8857 25639 8891
rect 4169 8789 4203 8823
rect 5641 8789 5675 8823
rect 7481 8789 7515 8823
rect 7757 8789 7791 8823
rect 11161 8789 11195 8823
rect 12449 8789 12483 8823
rect 16405 8789 16439 8823
rect 17693 8789 17727 8823
rect 18061 8789 18095 8823
rect 19733 8789 19767 8823
rect 22661 8789 22695 8823
rect 22753 8789 22787 8823
rect 24133 8789 24167 8823
rect 25329 8789 25363 8823
rect 4721 8585 4755 8619
rect 10149 8585 10183 8619
rect 20269 8585 20303 8619
rect 22569 8585 22603 8619
rect 6745 8517 6779 8551
rect 15945 8517 15979 8551
rect 21557 8517 21591 8551
rect 3525 8449 3559 8483
rect 4629 8449 4663 8483
rect 4905 8449 4939 8483
rect 6561 8449 6595 8483
rect 9505 8449 9539 8483
rect 11069 8449 11103 8483
rect 11253 8449 11287 8483
rect 12081 8449 12115 8483
rect 12633 8449 12667 8483
rect 14013 8449 14047 8483
rect 14197 8449 14231 8483
rect 14933 8449 14967 8483
rect 16957 8449 16991 8483
rect 17049 8449 17083 8483
rect 17509 8449 17543 8483
rect 17693 8449 17727 8483
rect 17969 8449 18003 8483
rect 18245 8449 18279 8483
rect 18613 8449 18647 8483
rect 20177 8449 20211 8483
rect 20453 8449 20487 8483
rect 20729 8449 20763 8483
rect 20821 8449 20855 8483
rect 21005 8449 21039 8483
rect 21373 8449 21407 8483
rect 21833 8449 21867 8483
rect 22017 8449 22051 8483
rect 22109 8449 22143 8483
rect 22293 8449 22327 8483
rect 22753 8449 22787 8483
rect 23305 8449 23339 8483
rect 25053 8449 25087 8483
rect 3433 8381 3467 8415
rect 6377 8381 6411 8415
rect 9597 8381 9631 8415
rect 10517 8381 10551 8415
rect 13921 8381 13955 8415
rect 16865 8381 16899 8415
rect 17141 8381 17175 8415
rect 18061 8381 18095 8415
rect 21189 8381 21223 8415
rect 25145 8381 25179 8415
rect 3893 8313 3927 8347
rect 9965 8313 9999 8347
rect 16681 8313 16715 8347
rect 20637 8313 20671 8347
rect 22201 8313 22235 8347
rect 24685 8313 24719 8347
rect 4905 8245 4939 8279
rect 9781 8245 9815 8279
rect 10149 8245 10183 8279
rect 11069 8245 11103 8279
rect 14013 8245 14047 8279
rect 20085 8245 20119 8279
rect 4997 8041 5031 8075
rect 12725 8041 12759 8075
rect 15209 8041 15243 8075
rect 19441 8041 19475 8075
rect 22753 8041 22787 8075
rect 24041 8041 24075 8075
rect 5457 7973 5491 8007
rect 13737 7973 13771 8007
rect 4353 7905 4387 7939
rect 4813 7905 4847 7939
rect 5089 7905 5123 7939
rect 11437 7905 11471 7939
rect 13093 7905 13127 7939
rect 13829 7905 13863 7939
rect 24133 7905 24167 7939
rect 4721 7837 4755 7871
rect 5273 7837 5307 7871
rect 6009 7837 6043 7871
rect 7665 7837 7699 7871
rect 7757 7837 7791 7871
rect 7849 7837 7883 7871
rect 8401 7837 8435 7871
rect 8493 7837 8527 7871
rect 8585 7837 8619 7871
rect 8953 7837 8987 7871
rect 9137 7837 9171 7871
rect 9781 7837 9815 7871
rect 9873 7837 9907 7871
rect 9965 7837 9999 7871
rect 10149 7837 10183 7871
rect 11345 7837 11379 7871
rect 13185 7837 13219 7871
rect 13369 7837 13403 7871
rect 14197 7837 14231 7871
rect 14565 7837 14599 7871
rect 14657 7837 14691 7871
rect 14933 7837 14967 7871
rect 15030 7837 15064 7871
rect 17601 7837 17635 7871
rect 17877 7837 17911 7871
rect 19625 7837 19659 7871
rect 19809 7837 19843 7871
rect 22109 7837 22143 7871
rect 22293 7837 22327 7871
rect 22569 7837 22603 7871
rect 23673 7837 23707 7871
rect 5641 7769 5675 7803
rect 7941 7769 7975 7803
rect 8217 7769 8251 7803
rect 12541 7769 12575 7803
rect 12741 7769 12775 7803
rect 14381 7769 14415 7803
rect 14841 7769 14875 7803
rect 17693 7769 17727 7803
rect 20085 7769 20119 7803
rect 23397 7769 23431 7803
rect 5825 7701 5859 7735
rect 8125 7701 8159 7735
rect 8953 7701 8987 7735
rect 9505 7701 9539 7735
rect 12081 7701 12115 7735
rect 12909 7701 12943 7735
rect 18061 7701 18095 7735
rect 19993 7701 20027 7735
rect 23765 7701 23799 7735
rect 23857 7701 23891 7735
rect 4537 7497 4571 7531
rect 4905 7497 4939 7531
rect 6745 7497 6779 7531
rect 11069 7497 11103 7531
rect 13645 7497 13679 7531
rect 18797 7497 18831 7531
rect 21189 7497 21223 7531
rect 23029 7497 23063 7531
rect 24961 7497 24995 7531
rect 25697 7497 25731 7531
rect 5825 7429 5859 7463
rect 5917 7429 5951 7463
rect 7205 7429 7239 7463
rect 7849 7429 7883 7463
rect 8493 7429 8527 7463
rect 8585 7429 8619 7463
rect 11253 7429 11287 7463
rect 20821 7429 20855 7463
rect 22845 7429 22879 7463
rect 23121 7429 23155 7463
rect 25881 7429 25915 7463
rect 4445 7361 4479 7395
rect 4629 7361 4663 7395
rect 4721 7361 4755 7395
rect 5549 7361 5583 7395
rect 5641 7361 5675 7395
rect 6009 7361 6043 7395
rect 6377 7361 6411 7395
rect 6561 7361 6595 7395
rect 6653 7361 6687 7395
rect 7389 7361 7423 7395
rect 7757 7361 7791 7395
rect 7941 7361 7975 7395
rect 8309 7361 8343 7395
rect 8677 7361 8711 7395
rect 9965 7361 9999 7395
rect 10701 7361 10735 7395
rect 10885 7361 10919 7395
rect 10977 7361 11011 7395
rect 11805 7361 11839 7395
rect 12725 7361 12759 7395
rect 13185 7361 13219 7395
rect 13277 7361 13311 7395
rect 13369 7361 13403 7395
rect 14289 7361 14323 7395
rect 14473 7361 14507 7395
rect 14749 7361 14783 7395
rect 15209 7361 15243 7395
rect 15393 7361 15427 7395
rect 17233 7361 17267 7395
rect 17325 7361 17359 7395
rect 17509 7361 17543 7395
rect 17601 7361 17635 7395
rect 17969 7361 18003 7395
rect 19809 7361 19843 7395
rect 19993 7361 20027 7395
rect 21127 7361 21161 7395
rect 21511 7361 21545 7395
rect 23213 7361 23247 7395
rect 24133 7361 24167 7395
rect 24317 7361 24351 7395
rect 25329 7361 25363 7395
rect 25605 7361 25639 7395
rect 7665 7293 7699 7327
rect 11713 7293 11747 7327
rect 12633 7293 12667 7327
rect 13461 7293 13495 7327
rect 14841 7293 14875 7327
rect 16221 7293 16255 7327
rect 18061 7293 18095 7327
rect 21649 7293 21683 7327
rect 24041 7293 24075 7327
rect 25421 7293 25455 7327
rect 6193 7225 6227 7259
rect 6469 7225 6503 7259
rect 7573 7225 7607 7259
rect 11253 7225 11287 7259
rect 21005 7225 21039 7259
rect 25881 7225 25915 7259
rect 8861 7157 8895 7191
rect 10057 7157 10091 7191
rect 10885 7157 10919 7191
rect 12817 7157 12851 7191
rect 17049 7157 17083 7191
rect 23397 7157 23431 7191
rect 24501 7157 24535 7191
rect 21097 6953 21131 6987
rect 21557 6953 21591 6987
rect 23765 6953 23799 6987
rect 17141 6885 17175 6919
rect 21741 6885 21775 6919
rect 22385 6885 22419 6919
rect 21373 6817 21407 6851
rect 21925 6817 21959 6851
rect 26249 6817 26283 6851
rect 6009 6749 6043 6783
rect 6193 6749 6227 6783
rect 6285 6749 6319 6783
rect 6469 6749 6503 6783
rect 9045 6749 9079 6783
rect 9229 6749 9263 6783
rect 10333 6749 10367 6783
rect 10425 6749 10459 6783
rect 10609 6749 10643 6783
rect 10701 6749 10735 6783
rect 10793 6749 10827 6783
rect 11069 6749 11103 6783
rect 15945 6749 15979 6783
rect 16129 6749 16163 6783
rect 16313 6749 16347 6783
rect 16405 6749 16439 6783
rect 16773 6749 16807 6783
rect 17049 6749 17083 6783
rect 17233 6749 17267 6783
rect 17417 6749 17451 6783
rect 19257 6749 19291 6783
rect 19717 6749 19751 6783
rect 19901 6749 19935 6783
rect 20177 6749 20211 6783
rect 21557 6749 21591 6783
rect 22017 6749 22051 6783
rect 23305 6749 23339 6783
rect 23581 6749 23615 6783
rect 23765 6749 23799 6783
rect 25053 6749 25087 6783
rect 25145 6749 25179 6783
rect 25329 6749 25363 6783
rect 25421 6749 25455 6783
rect 25513 6749 25547 6783
rect 25881 6749 25915 6783
rect 26157 6749 26191 6783
rect 10149 6681 10183 6715
rect 16037 6681 16071 6715
rect 16589 6681 16623 6715
rect 20729 6681 20763 6715
rect 20913 6681 20947 6715
rect 21281 6681 21315 6715
rect 24869 6681 24903 6715
rect 25697 6681 25731 6715
rect 25789 6681 25823 6715
rect 6193 6613 6227 6647
rect 6377 6613 6411 6647
rect 10057 6613 10091 6647
rect 10891 6613 10925 6647
rect 10977 6613 11011 6647
rect 19349 6613 19383 6647
rect 20361 6613 20395 6647
rect 23949 6613 23983 6647
rect 26065 6613 26099 6647
rect 4997 6409 5031 6443
rect 5641 6409 5675 6443
rect 8309 6409 8343 6443
rect 14749 6409 14783 6443
rect 14933 6409 14967 6443
rect 15577 6409 15611 6443
rect 16037 6409 16071 6443
rect 21005 6409 21039 6443
rect 23673 6409 23707 6443
rect 25421 6409 25455 6443
rect 5825 6341 5859 6375
rect 6653 6341 6687 6375
rect 13553 6341 13587 6375
rect 14013 6341 14047 6375
rect 18705 6341 18739 6375
rect 23305 6341 23339 6375
rect 4994 6273 5028 6307
rect 5365 6273 5399 6307
rect 5549 6273 5583 6307
rect 6377 6273 6411 6307
rect 6561 6273 6595 6307
rect 6745 6273 6779 6307
rect 7573 6273 7607 6307
rect 7757 6273 7791 6307
rect 10333 6273 10367 6307
rect 11805 6273 11839 6307
rect 12265 6273 12299 6307
rect 12449 6273 12483 6307
rect 12725 6273 12759 6307
rect 13001 6273 13035 6307
rect 13093 6273 13127 6307
rect 13277 6273 13311 6307
rect 13369 6273 13403 6307
rect 13829 6273 13863 6307
rect 14752 6273 14786 6307
rect 15209 6273 15243 6307
rect 15853 6273 15887 6307
rect 16129 6273 16163 6307
rect 18475 6273 18509 6307
rect 18613 6273 18647 6307
rect 18797 6273 18831 6307
rect 20637 6273 20671 6307
rect 20821 6273 20855 6307
rect 21097 6273 21131 6307
rect 21373 6273 21407 6307
rect 23213 6273 23247 6307
rect 23489 6273 23523 6307
rect 23765 6273 23799 6307
rect 23949 6273 23983 6307
rect 25329 6273 25363 6307
rect 5457 6205 5491 6239
rect 10425 6205 10459 6239
rect 11897 6205 11931 6239
rect 14289 6205 14323 6239
rect 14381 6205 14415 6239
rect 15117 6205 15151 6239
rect 18337 6205 18371 6239
rect 23857 6205 23891 6239
rect 5825 6137 5859 6171
rect 6929 6137 6963 6171
rect 10701 6137 10735 6171
rect 12173 6137 12207 6171
rect 12541 6137 12575 6171
rect 12633 6137 12667 6171
rect 13277 6137 13311 6171
rect 14197 6137 14231 6171
rect 18981 6137 19015 6171
rect 21189 6137 21223 6171
rect 4813 6069 4847 6103
rect 11805 6069 11839 6103
rect 12909 6069 12943 6103
rect 13737 6069 13771 6103
rect 15669 6069 15703 6103
rect 21097 6069 21131 6103
rect 11253 5865 11287 5899
rect 12633 5865 12667 5899
rect 12725 5865 12759 5899
rect 13093 5865 13127 5899
rect 14841 5865 14875 5899
rect 18429 5865 18463 5899
rect 20913 5865 20947 5899
rect 22017 5865 22051 5899
rect 25421 5865 25455 5899
rect 9965 5797 9999 5831
rect 11069 5797 11103 5831
rect 12173 5797 12207 5831
rect 12265 5797 12299 5831
rect 18889 5797 18923 5831
rect 21557 5797 21591 5831
rect 23857 5797 23891 5831
rect 23949 5797 23983 5831
rect 7481 5729 7515 5763
rect 7757 5729 7791 5763
rect 9505 5729 9539 5763
rect 12541 5729 12575 5763
rect 16957 5729 16991 5763
rect 20269 5729 20303 5763
rect 21097 5729 21131 5763
rect 25513 5729 25547 5763
rect 5917 5661 5951 5695
rect 6101 5661 6135 5695
rect 7389 5661 7423 5695
rect 9597 5661 9631 5695
rect 12081 5661 12115 5695
rect 12357 5661 12391 5695
rect 12817 5661 12851 5695
rect 13277 5661 13311 5695
rect 14473 5661 14507 5695
rect 16681 5661 16715 5695
rect 16865 5661 16899 5695
rect 17049 5661 17083 5695
rect 17420 5661 17454 5695
rect 17693 5661 17727 5695
rect 17877 5661 17911 5695
rect 17969 5661 18003 5695
rect 18245 5661 18279 5695
rect 18705 5661 18739 5695
rect 18981 5661 19015 5695
rect 19809 5661 19843 5695
rect 20361 5661 20395 5695
rect 20453 5661 20487 5695
rect 20920 5661 20954 5695
rect 21281 5661 21315 5695
rect 21557 5661 21591 5695
rect 21649 5661 21683 5695
rect 21925 5661 21959 5695
rect 22109 5661 22143 5695
rect 22201 5661 22235 5695
rect 22385 5661 22419 5695
rect 23765 5661 23799 5695
rect 24041 5661 24075 5695
rect 24994 5661 25028 5695
rect 10793 5593 10827 5627
rect 13461 5593 13495 5627
rect 14657 5593 14691 5627
rect 17785 5593 17819 5627
rect 18797 5593 18831 5627
rect 21189 5593 21223 5627
rect 21373 5593 21407 5627
rect 21741 5593 21775 5627
rect 6009 5525 6043 5559
rect 11897 5525 11931 5559
rect 16773 5525 16807 5559
rect 17417 5525 17451 5559
rect 17601 5525 17635 5559
rect 18061 5525 18095 5559
rect 20729 5525 20763 5559
rect 22293 5525 22327 5559
rect 23581 5525 23615 5559
rect 24869 5525 24903 5559
rect 25053 5525 25087 5559
rect 5825 5321 5859 5355
rect 6929 5321 6963 5355
rect 11897 5321 11931 5355
rect 17693 5321 17727 5355
rect 19901 5321 19935 5355
rect 22937 5321 22971 5355
rect 23673 5321 23707 5355
rect 25329 5321 25363 5355
rect 4445 5253 4479 5287
rect 13829 5253 13863 5287
rect 15945 5253 15979 5287
rect 18797 5253 18831 5287
rect 4997 5185 5031 5219
rect 5733 5185 5767 5219
rect 6009 5185 6043 5219
rect 6193 5185 6227 5219
rect 6469 5185 6503 5219
rect 6653 5185 6687 5219
rect 6745 5185 6779 5219
rect 7941 5185 7975 5219
rect 8217 5185 8251 5219
rect 8309 5185 8343 5219
rect 8769 5185 8803 5219
rect 9137 5185 9171 5219
rect 9597 5185 9631 5219
rect 11713 5185 11747 5219
rect 11989 5185 12023 5219
rect 12081 5185 12115 5219
rect 12265 5185 12299 5219
rect 13737 5185 13771 5219
rect 14013 5185 14047 5219
rect 14289 5185 14323 5219
rect 15117 5185 15151 5219
rect 16313 5185 16347 5219
rect 16497 5185 16531 5219
rect 16681 5185 16715 5219
rect 16773 5185 16807 5219
rect 16957 5185 16991 5219
rect 17049 5185 17083 5219
rect 17325 5185 17359 5219
rect 17693 5185 17727 5219
rect 18061 5185 18095 5219
rect 19809 5185 19843 5219
rect 19993 5185 20027 5219
rect 21465 5185 21499 5219
rect 21557 5185 21591 5219
rect 22109 5185 22143 5219
rect 22569 5185 22603 5219
rect 22661 5185 22695 5219
rect 23305 5185 23339 5219
rect 24685 5185 24719 5219
rect 24869 5185 24903 5219
rect 25145 5185 25179 5219
rect 6561 5117 6595 5151
rect 8033 5117 8067 5151
rect 8677 5117 8711 5151
rect 9965 5117 9999 5151
rect 14749 5117 14783 5151
rect 15025 5117 15059 5151
rect 16405 5117 16439 5151
rect 17877 5117 17911 5151
rect 22201 5117 22235 5151
rect 23213 5117 23247 5151
rect 4721 5049 4755 5083
rect 5273 5049 5307 5083
rect 14565 5049 14599 5083
rect 17233 5049 17267 5083
rect 4905 4981 4939 5015
rect 5457 4981 5491 5015
rect 8493 4981 8527 5015
rect 11529 4981 11563 5015
rect 12173 4981 12207 5015
rect 14013 4981 14047 5015
rect 22385 4981 22419 5015
rect 22569 4981 22603 5015
rect 14657 4777 14691 4811
rect 18429 4777 18463 4811
rect 20453 4777 20487 4811
rect 24593 4777 24627 4811
rect 6561 4709 6595 4743
rect 22109 4709 22143 4743
rect 25329 4709 25363 4743
rect 4721 4641 4755 4675
rect 6101 4641 6135 4675
rect 8493 4641 8527 4675
rect 8677 4641 8711 4675
rect 9045 4641 9079 4675
rect 9137 4641 9171 4675
rect 9229 4641 9263 4675
rect 9321 4641 9355 4675
rect 12633 4641 12667 4675
rect 13001 4641 13035 4675
rect 13369 4641 13403 4675
rect 14381 4641 14415 4675
rect 16405 4641 16439 4675
rect 18245 4641 18279 4675
rect 20545 4641 20579 4675
rect 25053 4641 25087 4675
rect 4813 4573 4847 4607
rect 5273 4573 5307 4607
rect 5457 4573 5491 4607
rect 6193 4573 6227 4607
rect 7481 4573 7515 4607
rect 8585 4573 8619 4607
rect 8769 4573 8803 4607
rect 10517 4573 10551 4607
rect 10701 4573 10735 4607
rect 12541 4573 12575 4607
rect 13185 4573 13219 4607
rect 14289 4573 14323 4607
rect 15577 4573 15611 4607
rect 15669 4573 15703 4607
rect 16313 4573 16347 4607
rect 16497 4573 16531 4607
rect 18153 4573 18187 4607
rect 20269 4573 20303 4607
rect 21925 4573 21959 4607
rect 22293 4573 22327 4607
rect 24409 4573 24443 4607
rect 24961 4573 24995 4607
rect 5641 4505 5675 4539
rect 5181 4437 5215 4471
rect 9505 4437 9539 4471
rect 10609 4437 10643 4471
rect 12909 4437 12943 4471
rect 15853 4437 15887 4471
rect 20085 4437 20119 4471
rect 22385 4437 22419 4471
rect 11529 4233 11563 4267
rect 24961 4233 24995 4267
rect 12173 4165 12207 4199
rect 15761 4165 15795 4199
rect 15945 4165 15979 4199
rect 24501 4165 24535 4199
rect 9781 4097 9815 4131
rect 9965 4097 9999 4131
rect 10057 4097 10091 4131
rect 10425 4097 10459 4131
rect 10885 4097 10919 4131
rect 10977 4097 11011 4131
rect 11069 4097 11103 4131
rect 11161 4097 11195 4131
rect 11713 4097 11747 4131
rect 14841 4097 14875 4131
rect 15209 4097 15243 4131
rect 15301 4097 15335 4131
rect 15485 4097 15519 4131
rect 15577 4097 15611 4131
rect 16313 4097 16347 4131
rect 17141 4097 17175 4131
rect 17325 4097 17359 4131
rect 19809 4097 19843 4131
rect 20085 4097 20119 4131
rect 20269 4097 20303 4131
rect 20545 4097 20579 4131
rect 21005 4097 21039 4131
rect 21373 4097 21407 4131
rect 22293 4097 22327 4131
rect 22753 4097 22787 4131
rect 23213 4097 23247 4131
rect 23397 4097 23431 4131
rect 23489 4097 23523 4131
rect 23857 4097 23891 4131
rect 24317 4097 24351 4131
rect 24593 4097 24627 4131
rect 24685 4097 24719 4131
rect 25421 4097 25455 4131
rect 25513 4097 25547 4131
rect 10609 4029 10643 4063
rect 10701 4029 10735 4063
rect 11805 4029 11839 4063
rect 21833 4029 21867 4063
rect 22201 4029 22235 4063
rect 22477 4029 22511 4063
rect 22569 4029 22603 4063
rect 23673 4029 23707 4063
rect 24041 4029 24075 4063
rect 10425 3961 10459 3995
rect 22937 3961 22971 3995
rect 25053 3961 25087 3995
rect 25697 3961 25731 3995
rect 9965 3893 9999 3927
rect 11805 3893 11839 3927
rect 15025 3893 15059 3927
rect 16957 3893 16991 3927
rect 23029 3893 23063 3927
rect 24869 3893 24903 3927
rect 19809 3689 19843 3723
rect 20453 3689 20487 3723
rect 21925 3689 21959 3723
rect 23489 3689 23523 3723
rect 23857 3689 23891 3723
rect 13921 3621 13955 3655
rect 15669 3621 15703 3655
rect 17693 3621 17727 3655
rect 18521 3621 18555 3655
rect 22109 3621 22143 3655
rect 22753 3621 22787 3655
rect 23121 3621 23155 3655
rect 25237 3621 25271 3655
rect 16681 3553 16715 3587
rect 17877 3553 17911 3587
rect 18061 3553 18095 3587
rect 20637 3553 20671 3587
rect 23305 3553 23339 3587
rect 24961 3553 24995 3587
rect 9045 3485 9079 3519
rect 11253 3485 11287 3519
rect 11437 3485 11471 3519
rect 11897 3485 11931 3519
rect 13553 3485 13587 3519
rect 13646 3485 13680 3519
rect 14105 3485 14139 3519
rect 14565 3485 14599 3519
rect 15025 3485 15059 3519
rect 15393 3485 15427 3519
rect 15761 3485 15795 3519
rect 16405 3485 16439 3519
rect 16497 3485 16531 3519
rect 16773 3485 16807 3519
rect 17049 3485 17083 3519
rect 17325 3485 17359 3519
rect 17417 3485 17451 3519
rect 18153 3485 18187 3519
rect 20085 3485 20119 3519
rect 20177 3485 20211 3519
rect 20545 3485 20579 3519
rect 20821 3485 20855 3519
rect 21085 3485 21119 3519
rect 21281 3485 21315 3519
rect 21741 3485 21775 3519
rect 21925 3485 21959 3519
rect 22201 3485 22235 3519
rect 22385 3485 22419 3519
rect 22569 3485 22603 3519
rect 23397 3485 23431 3519
rect 23581 3485 23615 3519
rect 23673 3485 23707 3519
rect 23857 3485 23891 3519
rect 24869 3485 24903 3519
rect 10057 3417 10091 3451
rect 11621 3417 11655 3451
rect 16865 3417 16899 3451
rect 17233 3417 17267 3451
rect 21005 3417 21039 3451
rect 21465 3417 21499 3451
rect 22477 3417 22511 3451
rect 22845 3417 22879 3451
rect 11805 3349 11839 3383
rect 16221 3349 16255 3383
rect 20269 3349 20303 3383
rect 21189 3349 21223 3383
rect 10149 3145 10183 3179
rect 10885 3145 10919 3179
rect 15945 3145 15979 3179
rect 16405 3145 16439 3179
rect 16973 3145 17007 3179
rect 17233 3145 17267 3179
rect 19717 3145 19751 3179
rect 20453 3145 20487 3179
rect 21373 3145 21407 3179
rect 22201 3145 22235 3179
rect 22569 3145 22603 3179
rect 10425 3077 10459 3111
rect 10517 3077 10551 3111
rect 12541 3077 12575 3111
rect 16037 3077 16071 3111
rect 16221 3077 16255 3111
rect 16773 3077 16807 3111
rect 20637 3077 20671 3111
rect 9781 3009 9815 3043
rect 10241 3009 10275 3043
rect 10609 3009 10643 3043
rect 11069 3009 11103 3043
rect 11253 3009 11287 3043
rect 11989 3009 12023 3043
rect 12449 3009 12483 3043
rect 12633 3009 12667 3043
rect 13277 3009 13311 3043
rect 13461 3009 13495 3043
rect 15209 3009 15243 3043
rect 15577 3009 15611 3043
rect 17417 3009 17451 3043
rect 18153 3009 18187 3043
rect 18337 3009 18371 3043
rect 18429 3009 18463 3043
rect 18705 3009 18739 3043
rect 18889 3009 18923 3043
rect 19993 3009 20027 3043
rect 20821 3009 20855 3043
rect 21281 3009 21315 3043
rect 21465 3009 21499 3043
rect 22109 3009 22143 3043
rect 1409 2941 1443 2975
rect 9873 2941 9907 2975
rect 12081 2941 12115 2975
rect 17509 2941 17543 2975
rect 17877 2941 17911 2975
rect 17969 2941 18003 2975
rect 19901 2941 19935 2975
rect 20361 2941 20395 2975
rect 21925 2941 21959 2975
rect 27537 2941 27571 2975
rect 10793 2873 10827 2907
rect 12357 2873 12391 2907
rect 17141 2873 17175 2907
rect 11069 2805 11103 2839
rect 16957 2805 16991 2839
rect 10425 2601 10459 2635
rect 12081 2601 12115 2635
rect 13553 2601 13587 2635
rect 15577 2601 15611 2635
rect 17877 2601 17911 2635
rect 15393 2533 15427 2567
rect 15761 2533 15795 2567
rect 10241 2397 10275 2431
rect 10425 2397 10459 2431
rect 11621 2397 11655 2431
rect 11897 2397 11931 2431
rect 13461 2397 13495 2431
rect 13645 2397 13679 2431
rect 15117 2397 15151 2431
rect 15669 2397 15703 2431
rect 15853 2397 15887 2431
rect 17693 2397 17727 2431
rect 17877 2397 17911 2431
rect 11713 2261 11747 2295
<< metal1 >>
rect 1104 28858 27876 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 27876 28858
rect 1104 28784 27876 28806
rect 5810 28704 5816 28756
rect 5868 28744 5874 28756
rect 6089 28747 6147 28753
rect 6089 28744 6101 28747
rect 5868 28716 6101 28744
rect 5868 28704 5874 28716
rect 6089 28713 6101 28716
rect 6135 28713 6147 28747
rect 6089 28707 6147 28713
rect 6454 28704 6460 28756
rect 6512 28744 6518 28756
rect 6549 28747 6607 28753
rect 6549 28744 6561 28747
rect 6512 28716 6561 28744
rect 6512 28704 6518 28716
rect 6549 28713 6561 28716
rect 6595 28713 6607 28747
rect 6549 28707 6607 28713
rect 9030 28704 9036 28756
rect 9088 28744 9094 28756
rect 9861 28747 9919 28753
rect 9861 28744 9873 28747
rect 9088 28716 9873 28744
rect 9088 28704 9094 28716
rect 9861 28713 9873 28716
rect 9907 28713 9919 28747
rect 9861 28707 9919 28713
rect 3234 28568 3240 28620
rect 3292 28608 3298 28620
rect 3329 28611 3387 28617
rect 3329 28608 3341 28611
rect 3292 28580 3341 28608
rect 3292 28568 3298 28580
rect 3329 28577 3341 28580
rect 3375 28577 3387 28611
rect 3329 28571 3387 28577
rect 4614 28500 4620 28552
rect 4672 28540 4678 28552
rect 4893 28543 4951 28549
rect 4893 28540 4905 28543
rect 4672 28512 4905 28540
rect 4672 28500 4678 28512
rect 4893 28509 4905 28512
rect 4939 28509 4951 28543
rect 4893 28503 4951 28509
rect 5534 28500 5540 28552
rect 5592 28540 5598 28552
rect 5905 28543 5963 28549
rect 5905 28540 5917 28543
rect 5592 28512 5917 28540
rect 5592 28500 5598 28512
rect 5905 28509 5917 28512
rect 5951 28509 5963 28543
rect 5905 28503 5963 28509
rect 6178 28500 6184 28552
rect 6236 28540 6242 28552
rect 6365 28543 6423 28549
rect 6365 28540 6377 28543
rect 6236 28512 6377 28540
rect 6236 28500 6242 28512
rect 6365 28509 6377 28512
rect 6411 28509 6423 28543
rect 8113 28543 8171 28549
rect 8113 28540 8125 28543
rect 6365 28503 6423 28509
rect 7760 28512 8125 28540
rect 7760 28484 7788 28512
rect 8113 28509 8125 28512
rect 8159 28509 8171 28543
rect 8113 28503 8171 28509
rect 8386 28500 8392 28552
rect 8444 28540 8450 28552
rect 8665 28543 8723 28549
rect 8665 28540 8677 28543
rect 8444 28512 8677 28540
rect 8444 28500 8450 28512
rect 8665 28509 8677 28512
rect 8711 28509 8723 28543
rect 8665 28503 8723 28509
rect 9122 28500 9128 28552
rect 9180 28540 9186 28552
rect 9493 28543 9551 28549
rect 9493 28540 9505 28543
rect 9180 28512 9505 28540
rect 9180 28500 9186 28512
rect 9493 28509 9505 28512
rect 9539 28509 9551 28543
rect 9493 28503 9551 28509
rect 9674 28500 9680 28552
rect 9732 28500 9738 28552
rect 12345 28543 12403 28549
rect 12345 28509 12357 28543
rect 12391 28509 12403 28543
rect 12345 28503 12403 28509
rect 4706 28432 4712 28484
rect 4764 28432 4770 28484
rect 7742 28432 7748 28484
rect 7800 28432 7806 28484
rect 7868 28475 7926 28481
rect 7868 28441 7880 28475
rect 7914 28472 7926 28475
rect 8941 28475 8999 28481
rect 8941 28472 8953 28475
rect 7914 28444 8953 28472
rect 7914 28441 7926 28444
rect 7868 28435 7926 28441
rect 8941 28441 8953 28444
rect 8987 28441 8999 28475
rect 12360 28472 12388 28503
rect 12526 28500 12532 28552
rect 12584 28500 12590 28552
rect 17034 28500 17040 28552
rect 17092 28500 17098 28552
rect 17221 28543 17279 28549
rect 17221 28509 17233 28543
rect 17267 28509 17279 28543
rect 17221 28503 17279 28509
rect 13170 28472 13176 28484
rect 12360 28444 13176 28472
rect 8941 28435 8999 28441
rect 13170 28432 13176 28444
rect 13228 28432 13234 28484
rect 16850 28432 16856 28484
rect 16908 28472 16914 28484
rect 17236 28472 17264 28503
rect 16908 28444 17264 28472
rect 16908 28432 16914 28444
rect 5077 28407 5135 28413
rect 5077 28373 5089 28407
rect 5123 28404 5135 28407
rect 6546 28404 6552 28416
rect 5123 28376 6552 28404
rect 5123 28373 5135 28376
rect 5077 28367 5135 28373
rect 6546 28364 6552 28376
rect 6604 28364 6610 28416
rect 6733 28407 6791 28413
rect 6733 28373 6745 28407
rect 6779 28404 6791 28407
rect 7282 28404 7288 28416
rect 6779 28376 7288 28404
rect 6779 28373 6791 28376
rect 6733 28367 6791 28373
rect 7282 28364 7288 28376
rect 7340 28364 7346 28416
rect 8478 28364 8484 28416
rect 8536 28364 8542 28416
rect 12437 28407 12495 28413
rect 12437 28373 12449 28407
rect 12483 28404 12495 28407
rect 12710 28404 12716 28416
rect 12483 28376 12716 28404
rect 12483 28373 12495 28376
rect 12437 28367 12495 28373
rect 12710 28364 12716 28376
rect 12768 28364 12774 28416
rect 17126 28364 17132 28416
rect 17184 28364 17190 28416
rect 1104 28314 27876 28336
rect 1104 28262 4874 28314
rect 4926 28262 4938 28314
rect 4990 28262 5002 28314
rect 5054 28262 5066 28314
rect 5118 28262 5130 28314
rect 5182 28262 27876 28314
rect 1104 28240 27876 28262
rect 4617 28203 4675 28209
rect 4617 28169 4629 28203
rect 4663 28200 4675 28203
rect 4706 28200 4712 28212
rect 4663 28172 4712 28200
rect 4663 28169 4675 28172
rect 4617 28163 4675 28169
rect 4706 28160 4712 28172
rect 4764 28160 4770 28212
rect 6178 28160 6184 28212
rect 6236 28160 6242 28212
rect 6917 28203 6975 28209
rect 6917 28169 6929 28203
rect 6963 28169 6975 28203
rect 6917 28163 6975 28169
rect 2768 28135 2826 28141
rect 2768 28101 2780 28135
rect 2814 28132 2826 28135
rect 2958 28132 2964 28144
rect 2814 28104 2964 28132
rect 2814 28101 2826 28104
rect 2768 28095 2826 28101
rect 2958 28092 2964 28104
rect 3016 28092 3022 28144
rect 4249 28135 4307 28141
rect 4249 28101 4261 28135
rect 4295 28132 4307 28135
rect 4798 28132 4804 28144
rect 4295 28104 4804 28132
rect 4295 28101 4307 28104
rect 4249 28095 4307 28101
rect 4798 28092 4804 28104
rect 4856 28092 4862 28144
rect 5552 28104 6500 28132
rect 1673 28067 1731 28073
rect 1673 28033 1685 28067
rect 1719 28064 1731 28067
rect 1762 28064 1768 28076
rect 1719 28036 1768 28064
rect 1719 28033 1731 28036
rect 1673 28027 1731 28033
rect 1762 28024 1768 28036
rect 1820 28024 1826 28076
rect 1854 28024 1860 28076
rect 1912 28024 1918 28076
rect 3326 28024 3332 28076
rect 3384 28064 3390 28076
rect 4458 28070 4516 28073
rect 4448 28067 4660 28070
rect 3384 28036 4384 28064
rect 4448 28036 4470 28067
rect 3384 28024 3390 28036
rect 1394 27956 1400 28008
rect 1452 27996 1458 28008
rect 4356 28005 4384 28036
rect 4458 28033 4470 28036
rect 4504 28064 4660 28067
rect 4709 28067 4767 28073
rect 4709 28064 4721 28067
rect 4504 28042 4721 28064
rect 4504 28033 4516 28042
rect 4632 28036 4721 28042
rect 4458 28027 4516 28033
rect 4709 28033 4721 28036
rect 4755 28064 4767 28067
rect 4890 28064 4896 28076
rect 4755 28036 4896 28064
rect 4755 28033 4767 28036
rect 4709 28027 4767 28033
rect 4890 28024 4896 28036
rect 4948 28024 4954 28076
rect 5552 28073 5580 28104
rect 4985 28067 5043 28073
rect 4985 28033 4997 28067
rect 5031 28033 5043 28067
rect 4985 28027 5043 28033
rect 5537 28067 5595 28073
rect 5537 28033 5549 28067
rect 5583 28033 5595 28067
rect 5537 28027 5595 28033
rect 2501 27999 2559 28005
rect 2501 27996 2513 27999
rect 1452 27968 2513 27996
rect 1452 27956 1458 27968
rect 2501 27965 2513 27968
rect 2547 27965 2559 27999
rect 3973 27999 4031 28005
rect 3973 27996 3985 27999
rect 2501 27959 2559 27965
rect 3896 27968 3985 27996
rect 3896 27928 3924 27968
rect 3973 27965 3985 27968
rect 4019 27965 4031 27999
rect 3973 27959 4031 27965
rect 4341 27999 4399 28005
rect 4341 27965 4353 27999
rect 4387 27996 4399 27999
rect 4801 27999 4859 28005
rect 4801 27996 4813 27999
rect 4387 27968 4813 27996
rect 4387 27965 4399 27968
rect 4341 27959 4399 27965
rect 4801 27965 4813 27968
rect 4847 27965 4859 27999
rect 4801 27959 4859 27965
rect 5000 27928 5028 28027
rect 5626 28024 5632 28076
rect 5684 28073 5690 28076
rect 5684 28067 5733 28073
rect 5684 28033 5687 28067
rect 5721 28033 5733 28067
rect 5684 28027 5733 28033
rect 5684 28024 5690 28027
rect 5810 28024 5816 28076
rect 5868 28024 5874 28076
rect 5902 28024 5908 28076
rect 5960 28024 5966 28076
rect 5997 28067 6055 28073
rect 5997 28033 6009 28067
rect 6043 28064 6055 28067
rect 6365 28067 6423 28073
rect 6043 28036 6132 28064
rect 6043 28033 6055 28036
rect 5997 28027 6055 28033
rect 3896 27900 5028 27928
rect 5169 27931 5227 27937
rect 3896 27872 3924 27900
rect 5169 27897 5181 27931
rect 5215 27928 5227 27931
rect 6104 27928 6132 28036
rect 6365 28033 6377 28067
rect 6411 28033 6423 28067
rect 6472 28064 6500 28104
rect 6546 28092 6552 28144
rect 6604 28092 6610 28144
rect 6638 28064 6644 28076
rect 6472 28036 6644 28064
rect 6365 28027 6423 28033
rect 6270 27956 6276 28008
rect 6328 27996 6334 28008
rect 6380 27996 6408 28027
rect 6638 28024 6644 28036
rect 6696 28024 6702 28076
rect 6730 28024 6736 28076
rect 6788 28024 6794 28076
rect 6932 28064 6960 28163
rect 7098 28160 7104 28212
rect 7156 28200 7162 28212
rect 7377 28203 7435 28209
rect 7377 28200 7389 28203
rect 7156 28172 7389 28200
rect 7156 28160 7162 28172
rect 7377 28169 7389 28172
rect 7423 28169 7435 28203
rect 7377 28163 7435 28169
rect 9122 28160 9128 28212
rect 9180 28160 9186 28212
rect 9309 28203 9367 28209
rect 9309 28169 9321 28203
rect 9355 28200 9367 28203
rect 9674 28200 9680 28212
rect 9355 28172 9680 28200
rect 9355 28169 9367 28172
rect 9309 28163 9367 28169
rect 8012 28135 8070 28141
rect 8012 28101 8024 28135
rect 8058 28132 8070 28135
rect 8478 28132 8484 28144
rect 8058 28104 8484 28132
rect 8058 28101 8070 28104
rect 8012 28095 8070 28101
rect 8478 28092 8484 28104
rect 8536 28092 8542 28144
rect 7193 28067 7251 28073
rect 7193 28064 7205 28067
rect 6932 28036 7205 28064
rect 7193 28033 7205 28036
rect 7239 28033 7251 28067
rect 9324 28064 9352 28163
rect 9674 28160 9680 28172
rect 9732 28160 9738 28212
rect 16574 28200 16580 28212
rect 16546 28160 16580 28200
rect 16632 28200 16638 28212
rect 17034 28200 17040 28212
rect 16632 28172 17040 28200
rect 16632 28160 16638 28172
rect 17034 28160 17040 28172
rect 17092 28200 17098 28212
rect 18049 28203 18107 28209
rect 18049 28200 18061 28203
rect 17092 28172 18061 28200
rect 17092 28160 17098 28172
rect 18049 28169 18061 28172
rect 18095 28169 18107 28203
rect 18049 28163 18107 28169
rect 14090 28132 14096 28144
rect 12636 28104 14096 28132
rect 7193 28027 7251 28033
rect 7300 28036 9352 28064
rect 7300 27996 7328 28036
rect 10410 28024 10416 28076
rect 10468 28073 10474 28076
rect 12636 28073 12664 28104
rect 14090 28092 14096 28104
rect 14148 28132 14154 28144
rect 16301 28135 16359 28141
rect 14148 28104 14504 28132
rect 14148 28092 14154 28104
rect 10468 28027 10480 28073
rect 10965 28067 11023 28073
rect 10965 28033 10977 28067
rect 11011 28064 11023 28067
rect 11793 28067 11851 28073
rect 11793 28064 11805 28067
rect 11011 28036 11805 28064
rect 11011 28033 11023 28036
rect 10965 28027 11023 28033
rect 11793 28033 11805 28036
rect 11839 28033 11851 28067
rect 11793 28027 11851 28033
rect 12621 28067 12679 28073
rect 12621 28033 12633 28067
rect 12667 28033 12679 28067
rect 12621 28027 12679 28033
rect 10468 28024 10474 28027
rect 12710 28024 12716 28076
rect 12768 28064 12774 28076
rect 14476 28073 14504 28104
rect 16301 28101 16313 28135
rect 16347 28132 16359 28135
rect 16546 28132 16574 28160
rect 18598 28132 18604 28144
rect 16347 28104 16574 28132
rect 16684 28104 18604 28132
rect 16347 28101 16359 28104
rect 16301 28095 16359 28101
rect 14734 28073 14740 28076
rect 12877 28067 12935 28073
rect 12877 28064 12889 28067
rect 12768 28036 12889 28064
rect 12768 28024 12774 28036
rect 12877 28033 12889 28036
rect 12923 28033 12935 28067
rect 12877 28027 12935 28033
rect 14461 28067 14519 28073
rect 14461 28033 14473 28067
rect 14507 28033 14519 28067
rect 14461 28027 14519 28033
rect 14728 28027 14740 28073
rect 14734 28024 14740 28027
rect 14792 28024 14798 28076
rect 16684 28073 16712 28104
rect 18598 28092 18604 28104
rect 18656 28132 18662 28144
rect 18656 28104 19564 28132
rect 18656 28092 18662 28104
rect 16485 28067 16543 28073
rect 16485 28033 16497 28067
rect 16531 28064 16543 28067
rect 16669 28067 16727 28073
rect 16531 28036 16620 28064
rect 16531 28033 16543 28036
rect 16485 28027 16543 28033
rect 6328 27968 7328 27996
rect 6328 27956 6334 27968
rect 7742 27956 7748 28008
rect 7800 27956 7806 28008
rect 10689 27999 10747 28005
rect 10689 27965 10701 27999
rect 10735 27996 10747 27999
rect 10870 27996 10876 28008
rect 10735 27968 10876 27996
rect 10735 27965 10747 27968
rect 10689 27959 10747 27965
rect 10870 27956 10876 27968
rect 10928 27956 10934 28008
rect 11057 27999 11115 28005
rect 11057 27996 11069 27999
rect 10980 27968 11069 27996
rect 10980 27940 11008 27968
rect 11057 27965 11069 27968
rect 11103 27965 11115 27999
rect 11057 27959 11115 27965
rect 12437 27999 12495 28005
rect 12437 27965 12449 27999
rect 12483 27965 12495 27999
rect 12437 27959 12495 27965
rect 5215 27900 6132 27928
rect 5215 27897 5227 27900
rect 5169 27891 5227 27897
rect 10962 27888 10968 27940
rect 11020 27888 11026 27940
rect 12452 27928 12480 27959
rect 12618 27928 12624 27940
rect 12452 27900 12624 27928
rect 12618 27888 12624 27900
rect 12676 27888 12682 27940
rect 1670 27820 1676 27872
rect 1728 27820 1734 27872
rect 3878 27820 3884 27872
rect 3936 27820 3942 27872
rect 4798 27820 4804 27872
rect 4856 27820 4862 27872
rect 5810 27820 5816 27872
rect 5868 27860 5874 27872
rect 6270 27860 6276 27872
rect 5868 27832 6276 27860
rect 5868 27820 5874 27832
rect 6270 27820 6276 27832
rect 6328 27820 6334 27872
rect 11330 27820 11336 27872
rect 11388 27820 11394 27872
rect 13998 27820 14004 27872
rect 14056 27820 14062 27872
rect 15746 27820 15752 27872
rect 15804 27860 15810 27872
rect 15841 27863 15899 27869
rect 15841 27860 15853 27863
rect 15804 27832 15853 27860
rect 15804 27820 15810 27832
rect 15841 27829 15853 27832
rect 15887 27829 15899 27863
rect 15841 27823 15899 27829
rect 16114 27820 16120 27872
rect 16172 27820 16178 27872
rect 16592 27860 16620 28036
rect 16669 28033 16681 28067
rect 16715 28033 16727 28067
rect 16669 28027 16727 28033
rect 16758 28024 16764 28076
rect 16816 28064 16822 28076
rect 19536 28073 19564 28104
rect 16925 28067 16983 28073
rect 16925 28064 16937 28067
rect 16816 28036 16937 28064
rect 16816 28024 16822 28036
rect 16925 28033 16937 28036
rect 16971 28033 16983 28067
rect 16925 28027 16983 28033
rect 19265 28067 19323 28073
rect 19265 28033 19277 28067
rect 19311 28064 19323 28067
rect 19521 28067 19579 28073
rect 19311 28036 19472 28064
rect 19311 28033 19323 28036
rect 19265 28027 19323 28033
rect 19444 27996 19472 28036
rect 19521 28033 19533 28067
rect 19567 28033 19579 28067
rect 19521 28027 19579 28033
rect 19613 27999 19671 28005
rect 19613 27996 19625 27999
rect 19444 27968 19625 27996
rect 19613 27965 19625 27968
rect 19659 27965 19671 27999
rect 19613 27959 19671 27965
rect 20165 27999 20223 28005
rect 20165 27965 20177 27999
rect 20211 27965 20223 27999
rect 20165 27959 20223 27965
rect 16850 27860 16856 27872
rect 16592 27832 16856 27860
rect 16850 27820 16856 27832
rect 16908 27820 16914 27872
rect 18138 27820 18144 27872
rect 18196 27820 18202 27872
rect 18230 27820 18236 27872
rect 18288 27860 18294 27872
rect 20180 27860 20208 27959
rect 18288 27832 20208 27860
rect 18288 27820 18294 27832
rect 1104 27770 27876 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 27876 27770
rect 1104 27696 27876 27718
rect 3142 27616 3148 27668
rect 3200 27656 3206 27668
rect 4525 27659 4583 27665
rect 3200 27628 3556 27656
rect 3200 27616 3206 27628
rect 3528 27588 3556 27628
rect 4525 27625 4537 27659
rect 4571 27656 4583 27659
rect 4706 27656 4712 27668
rect 4571 27628 4712 27656
rect 4571 27625 4583 27628
rect 4525 27619 4583 27625
rect 4706 27616 4712 27628
rect 4764 27616 4770 27668
rect 6181 27659 6239 27665
rect 6181 27625 6193 27659
rect 6227 27656 6239 27659
rect 6638 27656 6644 27668
rect 6227 27628 6644 27656
rect 6227 27625 6239 27628
rect 6181 27619 6239 27625
rect 6638 27616 6644 27628
rect 6696 27616 6702 27668
rect 12526 27616 12532 27668
rect 12584 27656 12590 27668
rect 12897 27659 12955 27665
rect 12897 27656 12909 27659
rect 12584 27628 12909 27656
rect 12584 27616 12590 27628
rect 12897 27625 12909 27628
rect 12943 27625 12955 27659
rect 12897 27619 12955 27625
rect 16209 27659 16267 27665
rect 16209 27625 16221 27659
rect 16255 27656 16267 27659
rect 17126 27656 17132 27668
rect 16255 27628 17132 27656
rect 16255 27625 16267 27628
rect 16209 27619 16267 27625
rect 17126 27616 17132 27628
rect 17184 27616 17190 27668
rect 4614 27588 4620 27600
rect 3528 27560 4620 27588
rect 4614 27548 4620 27560
rect 4672 27548 4678 27600
rect 4801 27591 4859 27597
rect 4801 27557 4813 27591
rect 4847 27588 4859 27591
rect 5902 27588 5908 27600
rect 4847 27560 5908 27588
rect 4847 27557 4859 27560
rect 4801 27551 4859 27557
rect 5902 27548 5908 27560
rect 5960 27548 5966 27600
rect 6270 27548 6276 27600
rect 6328 27548 6334 27600
rect 10410 27548 10416 27600
rect 10468 27548 10474 27600
rect 13909 27591 13967 27597
rect 13909 27588 13921 27591
rect 10612 27560 10824 27588
rect 1394 27480 1400 27532
rect 1452 27480 1458 27532
rect 2406 27480 2412 27532
rect 2464 27520 2470 27532
rect 3053 27523 3111 27529
rect 3053 27520 3065 27523
rect 2464 27492 3065 27520
rect 2464 27480 2470 27492
rect 3053 27489 3065 27492
rect 3099 27520 3111 27523
rect 3099 27492 4844 27520
rect 3099 27489 3111 27492
rect 3053 27483 3111 27489
rect 3712 27464 3740 27492
rect 4816 27464 4844 27492
rect 9674 27480 9680 27532
rect 9732 27480 9738 27532
rect 10321 27523 10379 27529
rect 10321 27489 10333 27523
rect 10367 27520 10379 27523
rect 10612 27520 10640 27560
rect 10367 27492 10640 27520
rect 10689 27523 10747 27529
rect 10367 27489 10379 27492
rect 10321 27483 10379 27489
rect 10689 27489 10701 27523
rect 10735 27489 10747 27523
rect 10689 27483 10747 27489
rect 1670 27461 1676 27464
rect 1664 27452 1676 27461
rect 1631 27424 1676 27452
rect 1664 27415 1676 27424
rect 1670 27412 1676 27415
rect 1728 27412 1734 27464
rect 2961 27455 3019 27461
rect 2961 27421 2973 27455
rect 3007 27452 3019 27455
rect 3326 27452 3332 27464
rect 3007 27424 3332 27452
rect 3007 27421 3019 27424
rect 2961 27415 3019 27421
rect 3326 27412 3332 27424
rect 3384 27412 3390 27464
rect 3418 27412 3424 27464
rect 3476 27412 3482 27464
rect 3605 27455 3663 27461
rect 3605 27421 3617 27455
rect 3651 27452 3663 27455
rect 3694 27452 3700 27464
rect 3651 27424 3700 27452
rect 3651 27421 3663 27424
rect 3605 27415 3663 27421
rect 3694 27412 3700 27424
rect 3752 27412 3758 27464
rect 4341 27455 4399 27461
rect 4341 27421 4353 27455
rect 4387 27421 4399 27455
rect 4341 27415 4399 27421
rect 2590 27344 2596 27396
rect 2648 27384 2654 27396
rect 3237 27387 3295 27393
rect 3237 27384 3249 27387
rect 2648 27356 3249 27384
rect 2648 27344 2654 27356
rect 3237 27353 3249 27356
rect 3283 27384 3295 27387
rect 3878 27384 3884 27396
rect 3283 27356 3884 27384
rect 3283 27353 3295 27356
rect 3237 27347 3295 27353
rect 3878 27344 3884 27356
rect 3936 27384 3942 27396
rect 4356 27384 4384 27415
rect 4798 27412 4804 27464
rect 4856 27412 4862 27464
rect 4985 27455 5043 27461
rect 4985 27421 4997 27455
rect 5031 27421 5043 27455
rect 4985 27415 5043 27421
rect 5000 27384 5028 27415
rect 6178 27412 6184 27464
rect 6236 27412 6242 27464
rect 7377 27455 7435 27461
rect 7377 27421 7389 27455
rect 7423 27452 7435 27455
rect 8846 27452 8852 27464
rect 7423 27424 8852 27452
rect 7423 27421 7435 27424
rect 7377 27415 7435 27421
rect 7760 27396 7788 27424
rect 8846 27412 8852 27424
rect 8904 27412 8910 27464
rect 3936 27356 5028 27384
rect 6549 27387 6607 27393
rect 3936 27344 3942 27356
rect 6549 27353 6561 27387
rect 6595 27384 6607 27387
rect 6822 27384 6828 27396
rect 6595 27356 6828 27384
rect 6595 27353 6607 27356
rect 6549 27347 6607 27353
rect 6822 27344 6828 27356
rect 6880 27384 6886 27396
rect 7466 27384 7472 27396
rect 6880 27356 7472 27384
rect 6880 27344 6886 27356
rect 7466 27344 7472 27356
rect 7524 27344 7530 27396
rect 7650 27393 7656 27396
rect 7644 27347 7656 27393
rect 7650 27344 7656 27347
rect 7708 27344 7714 27396
rect 7742 27344 7748 27396
rect 7800 27344 7806 27396
rect 10704 27384 10732 27483
rect 10796 27461 10824 27560
rect 13556 27560 13921 27588
rect 10870 27480 10876 27532
rect 10928 27520 10934 27532
rect 13556 27529 13584 27560
rect 13909 27557 13921 27560
rect 13955 27557 13967 27591
rect 13909 27551 13967 27557
rect 16393 27591 16451 27597
rect 16393 27557 16405 27591
rect 16439 27588 16451 27591
rect 16758 27588 16764 27600
rect 16439 27560 16764 27588
rect 16439 27557 16451 27560
rect 16393 27551 16451 27557
rect 16758 27548 16764 27560
rect 16816 27548 16822 27600
rect 17681 27591 17739 27597
rect 17681 27557 17693 27591
rect 17727 27588 17739 27591
rect 18230 27588 18236 27600
rect 17727 27560 18236 27588
rect 17727 27557 17739 27560
rect 17681 27551 17739 27557
rect 18230 27548 18236 27560
rect 18288 27548 18294 27600
rect 11241 27523 11299 27529
rect 11241 27520 11253 27523
rect 10928 27492 11253 27520
rect 10928 27480 10934 27492
rect 11241 27489 11253 27492
rect 11287 27489 11299 27523
rect 11241 27483 11299 27489
rect 13541 27523 13599 27529
rect 13541 27489 13553 27523
rect 13587 27489 13599 27523
rect 13541 27483 13599 27489
rect 13998 27480 14004 27532
rect 14056 27520 14062 27532
rect 14645 27523 14703 27529
rect 14645 27520 14657 27523
rect 14056 27492 14657 27520
rect 14056 27480 14062 27492
rect 14645 27489 14657 27492
rect 14691 27489 14703 27523
rect 14645 27483 14703 27489
rect 17126 27480 17132 27532
rect 17184 27520 17190 27532
rect 17221 27523 17279 27529
rect 17221 27520 17233 27523
rect 17184 27492 17233 27520
rect 17184 27480 17190 27492
rect 17221 27489 17233 27492
rect 17267 27489 17279 27523
rect 17221 27483 17279 27489
rect 18138 27480 18144 27532
rect 18196 27520 18202 27532
rect 18325 27523 18383 27529
rect 18325 27520 18337 27523
rect 18196 27492 18337 27520
rect 18196 27480 18202 27492
rect 18325 27489 18337 27492
rect 18371 27489 18383 27523
rect 18325 27483 18383 27489
rect 10781 27455 10839 27461
rect 10781 27421 10793 27455
rect 10827 27421 10839 27455
rect 10781 27415 10839 27421
rect 11330 27412 11336 27464
rect 11388 27452 11394 27464
rect 11497 27455 11555 27461
rect 11497 27452 11509 27455
rect 11388 27424 11509 27452
rect 11388 27412 11394 27424
rect 11497 27421 11509 27424
rect 11543 27421 11555 27455
rect 11497 27415 11555 27421
rect 13630 27412 13636 27464
rect 13688 27412 13694 27464
rect 13725 27455 13783 27461
rect 13725 27421 13737 27455
rect 13771 27452 13783 27455
rect 15746 27452 15752 27464
rect 13771 27424 15752 27452
rect 13771 27421 13783 27424
rect 13725 27415 13783 27421
rect 13354 27384 13360 27396
rect 10704 27356 12434 27384
rect 2777 27319 2835 27325
rect 2777 27285 2789 27319
rect 2823 27316 2835 27319
rect 3418 27316 3424 27328
rect 2823 27288 3424 27316
rect 2823 27285 2835 27288
rect 2777 27279 2835 27285
rect 3418 27276 3424 27288
rect 3476 27276 3482 27328
rect 3786 27276 3792 27328
rect 3844 27276 3850 27328
rect 6362 27276 6368 27328
rect 6420 27316 6426 27328
rect 6457 27319 6515 27325
rect 6457 27316 6469 27319
rect 6420 27288 6469 27316
rect 6420 27276 6426 27288
rect 6457 27285 6469 27288
rect 6503 27285 6515 27319
rect 6457 27279 6515 27285
rect 8754 27276 8760 27328
rect 8812 27276 8818 27328
rect 12406 27316 12434 27356
rect 12544 27356 13360 27384
rect 12544 27316 12572 27356
rect 13354 27344 13360 27356
rect 13412 27344 13418 27396
rect 13538 27344 13544 27396
rect 13596 27384 13602 27396
rect 13740 27384 13768 27415
rect 15746 27412 15752 27424
rect 15804 27412 15810 27464
rect 17313 27455 17371 27461
rect 17313 27421 17325 27455
rect 17359 27452 17371 27455
rect 17773 27455 17831 27461
rect 17773 27452 17785 27455
rect 17359 27424 17785 27452
rect 17359 27421 17371 27424
rect 17313 27415 17371 27421
rect 17773 27421 17785 27424
rect 17819 27421 17831 27455
rect 17773 27415 17831 27421
rect 13596 27356 13768 27384
rect 13909 27387 13967 27393
rect 13596 27344 13602 27356
rect 13909 27353 13921 27387
rect 13955 27384 13967 27387
rect 14093 27387 14151 27393
rect 14093 27384 14105 27387
rect 13955 27356 14105 27384
rect 13955 27353 13967 27356
rect 13909 27347 13967 27353
rect 14093 27353 14105 27356
rect 14139 27353 14151 27387
rect 15654 27384 15660 27396
rect 14093 27347 14151 27353
rect 14200 27356 15660 27384
rect 12406 27288 12572 27316
rect 12618 27276 12624 27328
rect 12676 27276 12682 27328
rect 13372 27316 13400 27344
rect 14200 27316 14228 27356
rect 15654 27344 15660 27356
rect 15712 27384 15718 27396
rect 16025 27387 16083 27393
rect 16025 27384 16037 27387
rect 15712 27356 16037 27384
rect 15712 27344 15718 27356
rect 16025 27353 16037 27356
rect 16071 27353 16083 27387
rect 16025 27347 16083 27353
rect 16114 27344 16120 27396
rect 16172 27384 16178 27396
rect 16225 27387 16283 27393
rect 16225 27384 16237 27387
rect 16172 27356 16237 27384
rect 16172 27344 16178 27356
rect 16225 27353 16237 27356
rect 16271 27353 16283 27387
rect 16225 27347 16283 27353
rect 13372 27288 14228 27316
rect 14274 27276 14280 27328
rect 14332 27316 14338 27328
rect 15105 27319 15163 27325
rect 15105 27316 15117 27319
rect 14332 27288 15117 27316
rect 14332 27276 14338 27288
rect 15105 27285 15117 27288
rect 15151 27285 15163 27319
rect 15105 27279 15163 27285
rect 1104 27226 27876 27248
rect 1104 27174 4874 27226
rect 4926 27174 4938 27226
rect 4990 27174 5002 27226
rect 5054 27174 5066 27226
rect 5118 27174 5130 27226
rect 5182 27174 27876 27226
rect 1104 27152 27876 27174
rect 1673 27115 1731 27121
rect 1673 27081 1685 27115
rect 1719 27112 1731 27115
rect 1762 27112 1768 27124
rect 1719 27084 1768 27112
rect 1719 27081 1731 27084
rect 1673 27075 1731 27081
rect 1762 27072 1768 27084
rect 1820 27072 1826 27124
rect 1854 27072 1860 27124
rect 1912 27112 1918 27124
rect 2041 27115 2099 27121
rect 2041 27112 2053 27115
rect 1912 27084 2053 27112
rect 1912 27072 1918 27084
rect 2041 27081 2053 27084
rect 2087 27081 2099 27115
rect 2041 27075 2099 27081
rect 3145 27115 3203 27121
rect 3145 27081 3157 27115
rect 3191 27112 3203 27115
rect 3786 27112 3792 27124
rect 3191 27084 3792 27112
rect 3191 27081 3203 27084
rect 3145 27075 3203 27081
rect 2056 27044 2084 27075
rect 3786 27072 3792 27084
rect 3844 27072 3850 27124
rect 7650 27072 7656 27124
rect 7708 27112 7714 27124
rect 7929 27115 7987 27121
rect 7929 27112 7941 27115
rect 7708 27084 7941 27112
rect 7708 27072 7714 27084
rect 7929 27081 7941 27084
rect 7975 27081 7987 27115
rect 13906 27112 13912 27124
rect 7929 27075 7987 27081
rect 12912 27084 13912 27112
rect 2056 27016 2728 27044
rect 1949 26979 2007 26985
rect 1949 26945 1961 26979
rect 1995 26945 2007 26979
rect 1949 26939 2007 26945
rect 1673 26911 1731 26917
rect 1673 26877 1685 26911
rect 1719 26877 1731 26911
rect 1964 26908 1992 26939
rect 2038 26936 2044 26988
rect 2096 26976 2102 26988
rect 2225 26979 2283 26985
rect 2225 26976 2237 26979
rect 2096 26948 2237 26976
rect 2096 26936 2102 26948
rect 2225 26945 2237 26948
rect 2271 26945 2283 26979
rect 2225 26939 2283 26945
rect 2406 26936 2412 26988
rect 2464 26936 2470 26988
rect 2590 26936 2596 26988
rect 2648 26936 2654 26988
rect 2700 26985 2728 27016
rect 2884 27016 3280 27044
rect 2685 26979 2743 26985
rect 2685 26945 2697 26979
rect 2731 26976 2743 26979
rect 2884 26976 2912 27016
rect 3252 26985 3280 27016
rect 4154 27004 4160 27056
rect 4212 27044 4218 27056
rect 4709 27047 4767 27053
rect 4709 27044 4721 27047
rect 4212 27016 4721 27044
rect 4212 27004 4218 27016
rect 4709 27013 4721 27016
rect 4755 27044 4767 27047
rect 4798 27044 4804 27056
rect 4755 27016 4804 27044
rect 4755 27013 4767 27016
rect 4709 27007 4767 27013
rect 4798 27004 4804 27016
rect 4856 27004 4862 27056
rect 8110 27053 8116 27056
rect 8097 27047 8116 27053
rect 8097 27013 8109 27047
rect 8097 27007 8116 27013
rect 8110 27004 8116 27007
rect 8168 27004 8174 27056
rect 8294 27004 8300 27056
rect 8352 27004 8358 27056
rect 2731 26948 2912 26976
rect 2961 26979 3019 26985
rect 2731 26945 2743 26948
rect 2685 26939 2743 26945
rect 2961 26945 2973 26979
rect 3007 26945 3019 26979
rect 2961 26939 3019 26945
rect 3237 26979 3295 26985
rect 3237 26945 3249 26979
rect 3283 26945 3295 26979
rect 3237 26939 3295 26945
rect 4525 26979 4583 26985
rect 4525 26945 4537 26979
rect 4571 26976 4583 26979
rect 4614 26976 4620 26988
rect 4571 26948 4620 26976
rect 4571 26945 4583 26948
rect 4525 26939 4583 26945
rect 2424 26908 2452 26936
rect 2866 26908 2872 26920
rect 1964 26880 2452 26908
rect 2516 26880 2872 26908
rect 1673 26871 1731 26877
rect 1688 26840 1716 26871
rect 2516 26840 2544 26880
rect 2866 26868 2872 26880
rect 2924 26868 2930 26920
rect 1688 26812 2544 26840
rect 2777 26843 2835 26849
rect 2777 26809 2789 26843
rect 2823 26840 2835 26843
rect 2976 26840 3004 26939
rect 4614 26936 4620 26948
rect 4672 26936 4678 26988
rect 5261 26979 5319 26985
rect 5261 26945 5273 26979
rect 5307 26976 5319 26979
rect 5810 26976 5816 26988
rect 5307 26948 5816 26976
rect 5307 26945 5319 26948
rect 5261 26939 5319 26945
rect 5810 26936 5816 26948
rect 5868 26936 5874 26988
rect 6638 26936 6644 26988
rect 6696 26976 6702 26988
rect 7193 26979 7251 26985
rect 7193 26976 7205 26979
rect 6696 26948 7205 26976
rect 6696 26936 6702 26948
rect 7193 26945 7205 26948
rect 7239 26945 7251 26979
rect 7193 26939 7251 26945
rect 9217 26979 9275 26985
rect 9217 26945 9229 26979
rect 9263 26945 9275 26979
rect 9217 26939 9275 26945
rect 9232 26908 9260 26939
rect 9306 26936 9312 26988
rect 9364 26936 9370 26988
rect 9490 26936 9496 26988
rect 9548 26936 9554 26988
rect 12434 26936 12440 26988
rect 12492 26936 12498 26988
rect 12912 26985 12940 27084
rect 13906 27072 13912 27084
rect 13964 27072 13970 27124
rect 14182 27112 14188 27124
rect 14016 27084 14188 27112
rect 13341 27047 13399 27053
rect 13341 27013 13353 27047
rect 13387 27044 13399 27047
rect 13387 27016 13492 27044
rect 13387 27013 13399 27016
rect 13341 27007 13399 27013
rect 12897 26979 12955 26985
rect 12897 26945 12909 26979
rect 12943 26945 12955 26979
rect 13464 26976 13492 27016
rect 13538 27004 13544 27056
rect 13596 27004 13602 27056
rect 13814 27053 13820 27056
rect 13801 27047 13820 27053
rect 13801 27013 13813 27047
rect 13801 27007 13820 27013
rect 13814 27004 13820 27007
rect 13872 27004 13878 27056
rect 14016 27053 14044 27084
rect 14182 27072 14188 27084
rect 14240 27072 14246 27124
rect 15654 27072 15660 27124
rect 15712 27112 15718 27124
rect 15749 27115 15807 27121
rect 15749 27112 15761 27115
rect 15712 27084 15761 27112
rect 15712 27072 15718 27084
rect 15749 27081 15761 27084
rect 15795 27081 15807 27115
rect 20809 27115 20867 27121
rect 20809 27112 20821 27115
rect 15749 27075 15807 27081
rect 18340 27084 20821 27112
rect 14001 27047 14059 27053
rect 14001 27013 14013 27047
rect 14047 27013 14059 27047
rect 14001 27007 14059 27013
rect 13630 26976 13636 26988
rect 13464 26948 13636 26976
rect 12897 26939 12955 26945
rect 13630 26936 13636 26948
rect 13688 26976 13694 26988
rect 13688 26948 14228 26976
rect 13688 26936 13694 26948
rect 9398 26908 9404 26920
rect 9232 26880 9404 26908
rect 9398 26868 9404 26880
rect 9456 26868 9462 26920
rect 9953 26911 10011 26917
rect 9953 26877 9965 26911
rect 9999 26877 10011 26911
rect 9953 26871 10011 26877
rect 12805 26911 12863 26917
rect 12805 26877 12817 26911
rect 12851 26908 12863 26911
rect 12986 26908 12992 26920
rect 12851 26880 12992 26908
rect 12851 26877 12863 26880
rect 12805 26871 12863 26877
rect 2823 26812 3004 26840
rect 9493 26843 9551 26849
rect 2823 26809 2835 26812
rect 2777 26803 2835 26809
rect 9493 26809 9505 26843
rect 9539 26840 9551 26843
rect 9968 26840 9996 26871
rect 12986 26868 12992 26880
rect 13044 26868 13050 26920
rect 14200 26917 14228 26948
rect 14274 26936 14280 26988
rect 14332 26936 14338 26988
rect 14366 26936 14372 26988
rect 14424 26976 14430 26988
rect 15470 26976 15476 26988
rect 14424 26948 15476 26976
rect 14424 26936 14430 26948
rect 15470 26936 15476 26948
rect 15528 26936 15534 26988
rect 15933 26979 15991 26985
rect 15933 26945 15945 26979
rect 15979 26976 15991 26979
rect 16022 26976 16028 26988
rect 15979 26948 16028 26976
rect 15979 26945 15991 26948
rect 15933 26939 15991 26945
rect 16022 26936 16028 26948
rect 16080 26936 16086 26988
rect 16209 26979 16267 26985
rect 16209 26945 16221 26979
rect 16255 26976 16267 26979
rect 16482 26976 16488 26988
rect 16255 26948 16488 26976
rect 16255 26945 16267 26948
rect 16209 26939 16267 26945
rect 16482 26936 16488 26948
rect 16540 26936 16546 26988
rect 16850 26936 16856 26988
rect 16908 26976 16914 26988
rect 17310 26976 17316 26988
rect 16908 26948 17316 26976
rect 16908 26936 16914 26948
rect 17310 26936 17316 26948
rect 17368 26976 17374 26988
rect 18340 26985 18368 27084
rect 20809 27081 20821 27084
rect 20855 27081 20867 27115
rect 20809 27075 20867 27081
rect 18417 27047 18475 27053
rect 18417 27013 18429 27047
rect 18463 27044 18475 27047
rect 18846 27047 18904 27053
rect 18846 27044 18858 27047
rect 18463 27016 18858 27044
rect 18463 27013 18475 27016
rect 18417 27007 18475 27013
rect 18846 27013 18858 27016
rect 18892 27013 18904 27047
rect 18846 27007 18904 27013
rect 18325 26979 18383 26985
rect 18325 26976 18337 26979
rect 17368 26948 18337 26976
rect 17368 26936 17374 26948
rect 18325 26945 18337 26948
rect 18371 26945 18383 26979
rect 18325 26939 18383 26945
rect 18506 26936 18512 26988
rect 18564 26936 18570 26988
rect 18598 26936 18604 26988
rect 18656 26936 18662 26988
rect 20990 26936 20996 26988
rect 21048 26936 21054 26988
rect 14185 26911 14243 26917
rect 13096 26880 14136 26908
rect 13096 26849 13124 26880
rect 9539 26812 9996 26840
rect 13081 26843 13139 26849
rect 9539 26809 9551 26812
rect 9493 26803 9551 26809
rect 13081 26809 13093 26843
rect 13127 26809 13139 26843
rect 13998 26840 14004 26852
rect 13081 26803 13139 26809
rect 13556 26812 14004 26840
rect 1857 26775 1915 26781
rect 1857 26741 1869 26775
rect 1903 26772 1915 26775
rect 1946 26772 1952 26784
rect 1903 26744 1952 26772
rect 1903 26741 1915 26744
rect 1857 26735 1915 26741
rect 1946 26732 1952 26744
rect 2004 26732 2010 26784
rect 2958 26732 2964 26784
rect 3016 26732 3022 26784
rect 4798 26732 4804 26784
rect 4856 26772 4862 26784
rect 4893 26775 4951 26781
rect 4893 26772 4905 26775
rect 4856 26744 4905 26772
rect 4856 26732 4862 26744
rect 4893 26741 4905 26744
rect 4939 26741 4951 26775
rect 4893 26735 4951 26741
rect 5166 26732 5172 26784
rect 5224 26732 5230 26784
rect 7101 26775 7159 26781
rect 7101 26741 7113 26775
rect 7147 26772 7159 26775
rect 7190 26772 7196 26784
rect 7147 26744 7196 26772
rect 7147 26741 7159 26744
rect 7101 26735 7159 26741
rect 7190 26732 7196 26744
rect 7248 26772 7254 26784
rect 7374 26772 7380 26784
rect 7248 26744 7380 26772
rect 7248 26732 7254 26744
rect 7374 26732 7380 26744
rect 7432 26732 7438 26784
rect 7834 26732 7840 26784
rect 7892 26772 7898 26784
rect 8113 26775 8171 26781
rect 8113 26772 8125 26775
rect 7892 26744 8125 26772
rect 7892 26732 7898 26744
rect 8113 26741 8125 26744
rect 8159 26741 8171 26775
rect 8113 26735 8171 26741
rect 10594 26732 10600 26784
rect 10652 26732 10658 26784
rect 12618 26732 12624 26784
rect 12676 26732 12682 26784
rect 13170 26732 13176 26784
rect 13228 26732 13234 26784
rect 13357 26775 13415 26781
rect 13357 26741 13369 26775
rect 13403 26772 13415 26775
rect 13556 26772 13584 26812
rect 13998 26800 14004 26812
rect 14056 26800 14062 26852
rect 14108 26840 14136 26880
rect 14185 26877 14197 26911
rect 14231 26877 14243 26911
rect 14185 26871 14243 26877
rect 14645 26911 14703 26917
rect 14645 26877 14657 26911
rect 14691 26908 14703 26911
rect 14734 26908 14740 26920
rect 14691 26880 14740 26908
rect 14691 26877 14703 26880
rect 14645 26871 14703 26877
rect 14734 26868 14740 26880
rect 14792 26868 14798 26920
rect 16114 26868 16120 26920
rect 16172 26868 16178 26920
rect 17126 26868 17132 26920
rect 17184 26868 17190 26920
rect 20625 26911 20683 26917
rect 20625 26877 20637 26911
rect 20671 26908 20683 26911
rect 21177 26911 21235 26917
rect 21177 26908 21189 26911
rect 20671 26880 21189 26908
rect 20671 26877 20683 26880
rect 20625 26871 20683 26877
rect 21177 26877 21189 26880
rect 21223 26877 21235 26911
rect 21177 26871 21235 26877
rect 14108 26812 15976 26840
rect 13403 26744 13584 26772
rect 13403 26741 13415 26744
rect 13357 26735 13415 26741
rect 13630 26732 13636 26784
rect 13688 26732 13694 26784
rect 13817 26775 13875 26781
rect 13817 26741 13829 26775
rect 13863 26772 13875 26775
rect 14274 26772 14280 26784
rect 13863 26744 14280 26772
rect 13863 26741 13875 26744
rect 13817 26735 13875 26741
rect 14274 26732 14280 26744
rect 14332 26732 14338 26784
rect 14366 26732 14372 26784
rect 14424 26772 14430 26784
rect 15948 26781 15976 26812
rect 17494 26800 17500 26852
rect 17552 26800 17558 26852
rect 19981 26843 20039 26849
rect 19981 26809 19993 26843
rect 20027 26840 20039 26843
rect 20640 26840 20668 26871
rect 20027 26812 20668 26840
rect 20027 26809 20039 26812
rect 19981 26803 20039 26809
rect 14921 26775 14979 26781
rect 14921 26772 14933 26775
rect 14424 26744 14933 26772
rect 14424 26732 14430 26744
rect 14921 26741 14933 26744
rect 14967 26741 14979 26775
rect 14921 26735 14979 26741
rect 15933 26775 15991 26781
rect 15933 26741 15945 26775
rect 15979 26741 15991 26775
rect 15933 26735 15991 26741
rect 17586 26732 17592 26784
rect 17644 26732 17650 26784
rect 20070 26732 20076 26784
rect 20128 26732 20134 26784
rect 1104 26682 27876 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 27876 26682
rect 1104 26608 27876 26630
rect 1210 26528 1216 26580
rect 1268 26568 1274 26580
rect 1857 26571 1915 26577
rect 1857 26568 1869 26571
rect 1268 26540 1869 26568
rect 1268 26528 1274 26540
rect 1857 26537 1869 26540
rect 1903 26537 1915 26571
rect 1857 26531 1915 26537
rect 3786 26528 3792 26580
rect 3844 26568 3850 26580
rect 4065 26571 4123 26577
rect 4065 26568 4077 26571
rect 3844 26540 4077 26568
rect 3844 26528 3850 26540
rect 4065 26537 4077 26540
rect 4111 26537 4123 26571
rect 4065 26531 4123 26537
rect 4525 26571 4583 26577
rect 4525 26537 4537 26571
rect 4571 26568 4583 26571
rect 4614 26568 4620 26580
rect 4571 26540 4620 26568
rect 4571 26537 4583 26540
rect 4525 26531 4583 26537
rect 4614 26528 4620 26540
rect 4672 26528 4678 26580
rect 5537 26571 5595 26577
rect 5537 26537 5549 26571
rect 5583 26568 5595 26571
rect 5626 26568 5632 26580
rect 5583 26540 5632 26568
rect 5583 26537 5595 26540
rect 5537 26531 5595 26537
rect 5166 26500 5172 26512
rect 2746 26472 5172 26500
rect 1673 26367 1731 26373
rect 1673 26333 1685 26367
rect 1719 26333 1731 26367
rect 1673 26327 1731 26333
rect 1688 26296 1716 26327
rect 1854 26324 1860 26376
rect 1912 26364 1918 26376
rect 2041 26367 2099 26373
rect 2041 26364 2053 26367
rect 1912 26336 2053 26364
rect 1912 26324 1918 26336
rect 2041 26333 2053 26336
rect 2087 26364 2099 26367
rect 2746 26364 2774 26472
rect 3878 26392 3884 26444
rect 3936 26432 3942 26444
rect 4249 26435 4307 26441
rect 4249 26432 4261 26435
rect 3936 26404 4261 26432
rect 3936 26392 3942 26404
rect 4249 26401 4261 26404
rect 4295 26401 4307 26435
rect 4249 26395 4307 26401
rect 2087 26336 2774 26364
rect 2869 26367 2927 26373
rect 2087 26333 2099 26336
rect 2041 26327 2099 26333
rect 2869 26333 2881 26367
rect 2915 26364 2927 26367
rect 2958 26364 2964 26376
rect 2915 26336 2964 26364
rect 2915 26333 2927 26336
rect 2869 26327 2927 26333
rect 2958 26324 2964 26336
rect 3016 26324 3022 26376
rect 3053 26367 3111 26373
rect 3053 26333 3065 26367
rect 3099 26364 3111 26367
rect 3142 26364 3148 26376
rect 3099 26336 3148 26364
rect 3099 26333 3111 26336
rect 3053 26327 3111 26333
rect 3142 26324 3148 26336
rect 3200 26324 3206 26376
rect 3326 26324 3332 26376
rect 3384 26364 3390 26376
rect 3694 26364 3700 26376
rect 3384 26336 3700 26364
rect 3384 26324 3390 26336
rect 3694 26324 3700 26336
rect 3752 26364 3758 26376
rect 3973 26367 4031 26373
rect 3973 26364 3985 26367
rect 3752 26336 3985 26364
rect 3752 26324 3758 26336
rect 3973 26333 3985 26336
rect 4019 26333 4031 26367
rect 3973 26327 4031 26333
rect 4430 26324 4436 26376
rect 4488 26364 4494 26376
rect 4798 26373 4804 26376
rect 4617 26367 4675 26373
rect 4617 26364 4629 26367
rect 4488 26336 4629 26364
rect 4488 26324 4494 26336
rect 4617 26333 4629 26336
rect 4663 26333 4675 26367
rect 4617 26327 4675 26333
rect 4775 26367 4804 26373
rect 4775 26333 4787 26367
rect 4775 26327 4804 26333
rect 4798 26324 4804 26327
rect 4856 26324 4862 26376
rect 4908 26373 4936 26472
rect 5166 26460 5172 26472
rect 5224 26500 5230 26512
rect 5350 26500 5356 26512
rect 5224 26472 5356 26500
rect 5224 26460 5230 26472
rect 5350 26460 5356 26472
rect 5408 26460 5414 26512
rect 5258 26392 5264 26444
rect 5316 26392 5322 26444
rect 4893 26367 4951 26373
rect 4893 26333 4905 26367
rect 4939 26333 4951 26367
rect 4893 26327 4951 26333
rect 4982 26324 4988 26376
rect 5040 26324 5046 26376
rect 5077 26367 5135 26373
rect 5077 26333 5089 26367
rect 5123 26364 5135 26367
rect 5552 26364 5580 26531
rect 5626 26528 5632 26540
rect 5684 26528 5690 26580
rect 6454 26528 6460 26580
rect 6512 26528 6518 26580
rect 6549 26571 6607 26577
rect 6549 26537 6561 26571
rect 6595 26568 6607 26571
rect 6730 26568 6736 26580
rect 6595 26540 6736 26568
rect 6595 26537 6607 26540
rect 6549 26531 6607 26537
rect 6730 26528 6736 26540
rect 6788 26528 6794 26580
rect 7374 26528 7380 26580
rect 7432 26528 7438 26580
rect 7466 26528 7472 26580
rect 7524 26568 7530 26580
rect 7837 26571 7895 26577
rect 7837 26568 7849 26571
rect 7524 26540 7849 26568
rect 7524 26528 7530 26540
rect 7837 26537 7849 26540
rect 7883 26537 7895 26571
rect 7837 26531 7895 26537
rect 8110 26528 8116 26580
rect 8168 26568 8174 26580
rect 8205 26571 8263 26577
rect 8205 26568 8217 26571
rect 8168 26540 8217 26568
rect 8168 26528 8174 26540
rect 8205 26537 8217 26540
rect 8251 26537 8263 26571
rect 8205 26531 8263 26537
rect 13725 26571 13783 26577
rect 13725 26537 13737 26571
rect 13771 26568 13783 26571
rect 13998 26568 14004 26580
rect 13771 26540 14004 26568
rect 13771 26537 13783 26540
rect 13725 26531 13783 26537
rect 13998 26528 14004 26540
rect 14056 26528 14062 26580
rect 15470 26528 15476 26580
rect 15528 26528 15534 26580
rect 16301 26571 16359 26577
rect 16301 26568 16313 26571
rect 16132 26540 16313 26568
rect 7006 26500 7012 26512
rect 6840 26472 7012 26500
rect 6362 26432 6368 26444
rect 5736 26404 6368 26432
rect 5736 26376 5764 26404
rect 6362 26392 6368 26404
rect 6420 26432 6426 26444
rect 6840 26441 6868 26472
rect 7006 26460 7012 26472
rect 7064 26460 7070 26512
rect 7098 26460 7104 26512
rect 7156 26500 7162 26512
rect 7193 26503 7251 26509
rect 7193 26500 7205 26503
rect 7156 26472 7205 26500
rect 7156 26460 7162 26472
rect 7193 26469 7205 26472
rect 7239 26469 7251 26503
rect 7193 26463 7251 26469
rect 12710 26460 12716 26512
rect 12768 26500 12774 26512
rect 13173 26503 13231 26509
rect 13173 26500 13185 26503
rect 12768 26472 13185 26500
rect 12768 26460 12774 26472
rect 13173 26469 13185 26472
rect 13219 26469 13231 26503
rect 13173 26463 13231 26469
rect 6825 26435 6883 26441
rect 6825 26432 6837 26435
rect 6420 26404 6837 26432
rect 6420 26392 6426 26404
rect 6825 26401 6837 26404
rect 6871 26401 6883 26435
rect 6825 26395 6883 26401
rect 6914 26392 6920 26444
rect 6972 26392 6978 26444
rect 8386 26432 8392 26444
rect 7852 26404 8392 26432
rect 5123 26336 5580 26364
rect 5123 26333 5135 26336
rect 5077 26327 5135 26333
rect 5718 26324 5724 26376
rect 5776 26324 5782 26376
rect 6181 26367 6239 26373
rect 6181 26333 6193 26367
rect 6227 26333 6239 26367
rect 6181 26327 6239 26333
rect 4062 26296 4068 26308
rect 1688 26268 4068 26296
rect 4062 26256 4068 26268
rect 4120 26256 4126 26308
rect 5902 26256 5908 26308
rect 5960 26256 5966 26308
rect 1486 26188 1492 26240
rect 1544 26188 1550 26240
rect 2774 26188 2780 26240
rect 2832 26228 2838 26240
rect 2869 26231 2927 26237
rect 2869 26228 2881 26231
rect 2832 26200 2881 26228
rect 2832 26188 2838 26200
rect 2869 26197 2881 26200
rect 2915 26197 2927 26231
rect 2869 26191 2927 26197
rect 5994 26188 6000 26240
rect 6052 26188 6058 26240
rect 6196 26228 6224 26327
rect 6270 26324 6276 26376
rect 6328 26324 6334 26376
rect 6546 26324 6552 26376
rect 6604 26364 6610 26376
rect 6707 26367 6765 26373
rect 6707 26364 6719 26367
rect 6604 26336 6719 26364
rect 6604 26324 6610 26336
rect 6707 26333 6719 26336
rect 6753 26333 6765 26367
rect 6707 26327 6765 26333
rect 7009 26367 7067 26373
rect 7009 26333 7021 26367
rect 7055 26333 7067 26367
rect 7009 26327 7067 26333
rect 6362 26256 6368 26308
rect 6420 26296 6426 26308
rect 6457 26299 6515 26305
rect 6457 26296 6469 26299
rect 6420 26268 6469 26296
rect 6420 26256 6426 26268
rect 6457 26265 6469 26268
rect 6503 26265 6515 26299
rect 7024 26296 7052 26327
rect 7466 26324 7472 26376
rect 7524 26324 7530 26376
rect 7852 26373 7880 26404
rect 8386 26392 8392 26404
rect 8444 26432 8450 26444
rect 9398 26432 9404 26444
rect 8444 26404 9404 26432
rect 8444 26392 8450 26404
rect 9398 26392 9404 26404
rect 9456 26392 9462 26444
rect 14090 26432 14096 26444
rect 12406 26404 14096 26432
rect 7561 26367 7619 26373
rect 7561 26333 7573 26367
rect 7607 26364 7619 26367
rect 7837 26367 7895 26373
rect 7837 26364 7849 26367
rect 7607 26336 7849 26364
rect 7607 26333 7619 26336
rect 7561 26327 7619 26333
rect 7837 26333 7849 26336
rect 7883 26333 7895 26367
rect 7837 26327 7895 26333
rect 7929 26367 7987 26373
rect 7929 26333 7941 26367
rect 7975 26364 7987 26367
rect 8481 26367 8539 26373
rect 8481 26364 8493 26367
rect 7975 26336 8493 26364
rect 7975 26333 7987 26336
rect 7929 26327 7987 26333
rect 8481 26333 8493 26336
rect 8527 26333 8539 26367
rect 8481 26327 8539 26333
rect 7190 26296 7196 26308
rect 6457 26259 6515 26265
rect 6564 26268 7196 26296
rect 6564 26228 6592 26268
rect 7190 26256 7196 26268
rect 7248 26256 7254 26308
rect 7944 26296 7972 26327
rect 8570 26324 8576 26376
rect 8628 26324 8634 26376
rect 8665 26367 8723 26373
rect 8665 26333 8677 26367
rect 8711 26333 8723 26367
rect 8665 26327 8723 26333
rect 10433 26367 10491 26373
rect 10433 26333 10445 26367
rect 10479 26364 10491 26367
rect 10594 26364 10600 26376
rect 10479 26336 10600 26364
rect 10479 26333 10491 26336
rect 10433 26327 10491 26333
rect 7883 26268 7972 26296
rect 6196 26200 6592 26228
rect 6638 26188 6644 26240
rect 6696 26228 6702 26240
rect 7883 26228 7911 26268
rect 8202 26256 8208 26308
rect 8260 26296 8266 26308
rect 8680 26296 8708 26327
rect 10594 26324 10600 26336
rect 10652 26324 10658 26376
rect 10689 26367 10747 26373
rect 10689 26333 10701 26367
rect 10735 26364 10747 26367
rect 10781 26367 10839 26373
rect 10781 26364 10793 26367
rect 10735 26336 10793 26364
rect 10735 26333 10747 26336
rect 10689 26327 10747 26333
rect 10781 26333 10793 26336
rect 10827 26364 10839 26367
rect 10870 26364 10876 26376
rect 10827 26336 10876 26364
rect 10827 26333 10839 26336
rect 10781 26327 10839 26333
rect 10870 26324 10876 26336
rect 10928 26364 10934 26376
rect 11606 26364 11612 26376
rect 10928 26336 11612 26364
rect 10928 26324 10934 26336
rect 11606 26324 11612 26336
rect 11664 26364 11670 26376
rect 12406 26364 12434 26404
rect 14090 26392 14096 26404
rect 14148 26392 14154 26444
rect 16132 26432 16160 26540
rect 16301 26537 16313 26540
rect 16347 26537 16359 26571
rect 16301 26531 16359 26537
rect 16482 26528 16488 26580
rect 16540 26528 16546 26580
rect 16666 26528 16672 26580
rect 16724 26568 16730 26580
rect 17126 26568 17132 26580
rect 16724 26540 17132 26568
rect 16724 26528 16730 26540
rect 17126 26528 17132 26540
rect 17184 26528 17190 26580
rect 18506 26528 18512 26580
rect 18564 26568 18570 26580
rect 19613 26571 19671 26577
rect 19613 26568 19625 26571
rect 18564 26540 19625 26568
rect 18564 26528 18570 26540
rect 19613 26537 19625 26540
rect 19659 26537 19671 26571
rect 19613 26531 19671 26537
rect 16574 26500 16580 26512
rect 16546 26460 16580 26500
rect 16632 26460 16638 26512
rect 16546 26432 16574 26460
rect 20990 26432 20996 26444
rect 16132 26404 16574 26432
rect 19628 26404 20996 26432
rect 11664 26336 12434 26364
rect 12529 26367 12587 26373
rect 11664 26324 11670 26336
rect 12529 26333 12541 26367
rect 12575 26364 12587 26367
rect 12575 26336 12609 26364
rect 12575 26333 12587 26336
rect 12529 26327 12587 26333
rect 8260 26268 8708 26296
rect 11048 26299 11106 26305
rect 8260 26256 8266 26268
rect 11048 26265 11060 26299
rect 11094 26296 11106 26299
rect 11238 26296 11244 26308
rect 11094 26268 11244 26296
rect 11094 26265 11106 26268
rect 11048 26259 11106 26265
rect 11238 26256 11244 26268
rect 11296 26256 11302 26308
rect 12544 26296 12572 26327
rect 13262 26324 13268 26376
rect 13320 26364 13326 26376
rect 13449 26367 13507 26373
rect 13449 26364 13461 26367
rect 13320 26336 13461 26364
rect 13320 26324 13326 26336
rect 13449 26333 13461 26336
rect 13495 26333 13507 26367
rect 13449 26327 13507 26333
rect 14182 26324 14188 26376
rect 14240 26364 14246 26376
rect 15102 26364 15108 26376
rect 14240 26336 15108 26364
rect 14240 26324 14246 26336
rect 15102 26324 15108 26336
rect 15160 26364 15166 26376
rect 15841 26367 15899 26373
rect 15841 26364 15853 26367
rect 15160 26336 15853 26364
rect 15160 26324 15166 26336
rect 15841 26333 15853 26336
rect 15887 26333 15899 26367
rect 15841 26327 15899 26333
rect 15930 26324 15936 26376
rect 15988 26324 15994 26376
rect 16301 26367 16359 26373
rect 16301 26333 16313 26367
rect 16347 26364 16359 26367
rect 16347 26336 17264 26364
rect 16347 26333 16359 26336
rect 16301 26327 16359 26333
rect 17236 26308 17264 26336
rect 17586 26324 17592 26376
rect 17644 26364 17650 26376
rect 18426 26367 18484 26373
rect 18426 26364 18438 26367
rect 17644 26336 18438 26364
rect 17644 26324 17650 26336
rect 18426 26333 18438 26336
rect 18472 26333 18484 26367
rect 18426 26327 18484 26333
rect 18598 26324 18604 26376
rect 18656 26364 18662 26376
rect 19628 26373 19656 26404
rect 20990 26392 20996 26404
rect 21048 26392 21054 26444
rect 18693 26367 18751 26373
rect 18693 26364 18705 26367
rect 18656 26336 18705 26364
rect 18656 26324 18662 26336
rect 18693 26333 18705 26336
rect 18739 26333 18751 26367
rect 18693 26327 18751 26333
rect 19613 26367 19671 26373
rect 19613 26333 19625 26367
rect 19659 26333 19671 26367
rect 19613 26327 19671 26333
rect 19797 26367 19855 26373
rect 19797 26333 19809 26367
rect 19843 26364 19855 26367
rect 20070 26364 20076 26376
rect 19843 26336 20076 26364
rect 19843 26333 19855 26336
rect 19797 26327 19855 26333
rect 20070 26324 20076 26336
rect 20128 26324 20134 26376
rect 12986 26296 12992 26308
rect 12176 26268 12992 26296
rect 6696 26200 7911 26228
rect 9309 26231 9367 26237
rect 6696 26188 6702 26200
rect 9309 26197 9321 26231
rect 9355 26228 9367 26231
rect 9398 26228 9404 26240
rect 9355 26200 9404 26228
rect 9355 26197 9367 26200
rect 9309 26191 9367 26197
rect 9398 26188 9404 26200
rect 9456 26188 9462 26240
rect 12176 26237 12204 26268
rect 12986 26256 12992 26268
rect 13044 26256 13050 26308
rect 13081 26299 13139 26305
rect 13081 26265 13093 26299
rect 13127 26296 13139 26299
rect 13173 26299 13231 26305
rect 13173 26296 13185 26299
rect 13127 26268 13185 26296
rect 13127 26265 13139 26268
rect 13081 26259 13139 26265
rect 13173 26265 13185 26268
rect 13219 26265 13231 26299
rect 13173 26259 13231 26265
rect 13538 26256 13544 26308
rect 13596 26256 13602 26308
rect 14338 26299 14396 26305
rect 14338 26296 14350 26299
rect 13924 26268 14350 26296
rect 12161 26231 12219 26237
rect 12161 26197 12173 26231
rect 12207 26197 12219 26231
rect 12161 26191 12219 26197
rect 12434 26188 12440 26240
rect 12492 26228 12498 26240
rect 13262 26228 13268 26240
rect 12492 26200 13268 26228
rect 12492 26188 12498 26200
rect 13262 26188 13268 26200
rect 13320 26228 13326 26240
rect 13357 26231 13415 26237
rect 13357 26228 13369 26231
rect 13320 26200 13369 26228
rect 13320 26188 13326 26200
rect 13357 26197 13369 26200
rect 13403 26197 13415 26231
rect 13357 26191 13415 26197
rect 13722 26188 13728 26240
rect 13780 26237 13786 26240
rect 13924 26237 13952 26268
rect 14338 26265 14350 26268
rect 14384 26265 14396 26299
rect 14338 26259 14396 26265
rect 16850 26256 16856 26308
rect 16908 26256 16914 26308
rect 16942 26256 16948 26308
rect 17000 26296 17006 26308
rect 17000 26268 17172 26296
rect 17000 26256 17006 26268
rect 13780 26231 13799 26237
rect 13787 26197 13799 26231
rect 13780 26191 13799 26197
rect 13909 26231 13967 26237
rect 13909 26197 13921 26231
rect 13955 26228 13967 26231
rect 13955 26200 13989 26228
rect 13955 26197 13967 26200
rect 13909 26191 13967 26197
rect 13780 26188 13786 26191
rect 16574 26188 16580 26240
rect 16632 26228 16638 26240
rect 17034 26228 17040 26240
rect 16632 26200 17040 26228
rect 16632 26188 16638 26200
rect 17034 26188 17040 26200
rect 17092 26188 17098 26240
rect 17144 26228 17172 26268
rect 17218 26256 17224 26308
rect 17276 26296 17282 26308
rect 18138 26296 18144 26308
rect 17276 26268 18144 26296
rect 17276 26256 17282 26268
rect 18138 26256 18144 26268
rect 18196 26256 18202 26308
rect 17313 26231 17371 26237
rect 17313 26228 17325 26231
rect 17144 26200 17325 26228
rect 17313 26197 17325 26200
rect 17359 26197 17371 26231
rect 17313 26191 17371 26197
rect 1104 26138 27876 26160
rect 1104 26086 4874 26138
rect 4926 26086 4938 26138
rect 4990 26086 5002 26138
rect 5054 26086 5066 26138
rect 5118 26086 5130 26138
rect 5182 26086 27876 26138
rect 1104 26064 27876 26086
rect 2041 26027 2099 26033
rect 2041 25993 2053 26027
rect 2087 26024 2099 26027
rect 2225 26027 2283 26033
rect 2225 26024 2237 26027
rect 2087 25996 2237 26024
rect 2087 25993 2099 25996
rect 2041 25987 2099 25993
rect 2225 25993 2237 25996
rect 2271 25993 2283 26027
rect 2225 25987 2283 25993
rect 2590 25984 2596 26036
rect 2648 26024 2654 26036
rect 3878 26024 3884 26036
rect 2648 25996 3884 26024
rect 2648 25984 2654 25996
rect 2774 25956 2780 25968
rect 2148 25928 2780 25956
rect 1854 25848 1860 25900
rect 1912 25848 1918 25900
rect 2148 25897 2176 25928
rect 2774 25916 2780 25928
rect 2832 25916 2838 25968
rect 2869 25959 2927 25965
rect 2869 25925 2881 25959
rect 2915 25956 2927 25959
rect 3602 25956 3608 25968
rect 2915 25928 3608 25956
rect 2915 25925 2927 25928
rect 2869 25919 2927 25925
rect 3602 25916 3608 25928
rect 3660 25916 3666 25968
rect 2133 25891 2191 25897
rect 2133 25857 2145 25891
rect 2179 25857 2191 25891
rect 2133 25851 2191 25857
rect 2409 25891 2467 25897
rect 2409 25857 2421 25891
rect 2455 25888 2467 25891
rect 2498 25888 2504 25900
rect 2455 25860 2504 25888
rect 2455 25857 2467 25860
rect 2409 25851 2467 25857
rect 2498 25848 2504 25860
rect 2556 25848 2562 25900
rect 2958 25848 2964 25900
rect 3016 25888 3022 25900
rect 3329 25891 3387 25897
rect 3329 25888 3341 25891
rect 3016 25860 3341 25888
rect 3016 25848 3022 25860
rect 3329 25857 3341 25860
rect 3375 25857 3387 25891
rect 3329 25851 3387 25857
rect 2593 25823 2651 25829
rect 2593 25789 2605 25823
rect 2639 25820 2651 25823
rect 3234 25820 3240 25832
rect 2639 25792 3240 25820
rect 2639 25789 2651 25792
rect 2593 25783 2651 25789
rect 3234 25780 3240 25792
rect 3292 25780 3298 25832
rect 3344 25820 3372 25851
rect 3418 25848 3424 25900
rect 3476 25848 3482 25900
rect 3804 25897 3832 25996
rect 3878 25984 3884 25996
rect 3936 25984 3942 26036
rect 4062 25984 4068 26036
rect 4120 25984 4126 26036
rect 4982 26024 4988 26036
rect 4172 25996 4988 26024
rect 3970 25916 3976 25968
rect 4028 25956 4034 25968
rect 4172 25956 4200 25996
rect 4982 25984 4988 25996
rect 5040 25984 5046 26036
rect 5534 25984 5540 26036
rect 5592 25984 5598 26036
rect 5902 25984 5908 26036
rect 5960 26024 5966 26036
rect 6730 26024 6736 26036
rect 5960 25996 6736 26024
rect 5960 25984 5966 25996
rect 6730 25984 6736 25996
rect 6788 25984 6794 26036
rect 7190 25984 7196 26036
rect 7248 25984 7254 26036
rect 8941 26027 8999 26033
rect 8941 26024 8953 26027
rect 8220 25996 8953 26024
rect 4430 25956 4436 25968
rect 4028 25928 4200 25956
rect 4264 25928 4436 25956
rect 4028 25916 4034 25928
rect 3789 25891 3847 25897
rect 3789 25857 3801 25891
rect 3835 25888 3847 25891
rect 4062 25888 4068 25900
rect 3835 25860 4068 25888
rect 3835 25857 3847 25860
rect 3789 25851 3847 25857
rect 4062 25848 4068 25860
rect 4120 25848 4126 25900
rect 4264 25897 4292 25928
rect 4430 25916 4436 25928
rect 4488 25956 4494 25968
rect 4706 25956 4712 25968
rect 4488 25928 4712 25956
rect 4488 25916 4494 25928
rect 4706 25916 4712 25928
rect 4764 25916 4770 25968
rect 5350 25956 5356 25968
rect 5276 25928 5356 25956
rect 4249 25891 4307 25897
rect 4249 25857 4261 25891
rect 4295 25857 4307 25891
rect 4249 25851 4307 25857
rect 4341 25891 4399 25897
rect 4341 25857 4353 25891
rect 4387 25888 4399 25891
rect 4614 25888 4620 25900
rect 4387 25860 4620 25888
rect 4387 25857 4399 25860
rect 4341 25851 4399 25857
rect 4614 25848 4620 25860
rect 4672 25848 4678 25900
rect 5276 25897 5304 25928
rect 5350 25916 5356 25928
rect 5408 25916 5414 25968
rect 6365 25959 6423 25965
rect 6365 25925 6377 25959
rect 6411 25956 6423 25959
rect 6454 25956 6460 25968
rect 6411 25928 6460 25956
rect 6411 25925 6423 25928
rect 6365 25919 6423 25925
rect 6454 25916 6460 25928
rect 6512 25956 6518 25968
rect 6512 25928 6684 25956
rect 6512 25916 6518 25928
rect 5261 25891 5319 25897
rect 5261 25857 5273 25891
rect 5307 25857 5319 25891
rect 5261 25851 5319 25857
rect 6270 25848 6276 25900
rect 6328 25888 6334 25900
rect 6546 25888 6552 25900
rect 6328 25860 6552 25888
rect 6328 25848 6334 25860
rect 6546 25848 6552 25860
rect 6604 25848 6610 25900
rect 6656 25888 6684 25928
rect 7006 25916 7012 25968
rect 7064 25956 7070 25968
rect 7377 25959 7435 25965
rect 7377 25956 7389 25959
rect 7064 25928 7389 25956
rect 7064 25916 7070 25928
rect 7377 25925 7389 25928
rect 7423 25956 7435 25959
rect 8220 25956 8248 25996
rect 8941 25993 8953 25996
rect 8987 25993 8999 26027
rect 8941 25987 8999 25993
rect 9309 26027 9367 26033
rect 9309 25993 9321 26027
rect 9355 26024 9367 26027
rect 9490 26024 9496 26036
rect 9355 25996 9496 26024
rect 9355 25993 9367 25996
rect 9309 25987 9367 25993
rect 9490 25984 9496 25996
rect 9548 25984 9554 26036
rect 11238 25984 11244 26036
rect 11296 25984 11302 26036
rect 12973 26027 13031 26033
rect 12973 25993 12985 26027
rect 13019 26024 13031 26027
rect 13078 26024 13084 26036
rect 13019 25996 13084 26024
rect 13019 25993 13031 25996
rect 12973 25987 13031 25993
rect 13078 25984 13084 25996
rect 13136 26024 13142 26036
rect 13446 26024 13452 26036
rect 13136 25996 13452 26024
rect 13136 25984 13142 25996
rect 13446 25984 13452 25996
rect 13504 25984 13510 26036
rect 13722 25984 13728 26036
rect 13780 25984 13786 26036
rect 14090 25984 14096 26036
rect 14148 25984 14154 26036
rect 14182 25984 14188 26036
rect 14240 26024 14246 26036
rect 14461 26027 14519 26033
rect 14461 26024 14473 26027
rect 14240 25996 14473 26024
rect 14240 25984 14246 25996
rect 14461 25993 14473 25996
rect 14507 25993 14519 26027
rect 14461 25987 14519 25993
rect 16114 25984 16120 26036
rect 16172 25984 16178 26036
rect 17494 25984 17500 26036
rect 17552 25984 17558 26036
rect 21082 25984 21088 26036
rect 21140 25984 21146 26036
rect 13173 25959 13231 25965
rect 7423 25928 8248 25956
rect 7423 25925 7435 25928
rect 7377 25919 7435 25925
rect 8220 25900 8248 25928
rect 8588 25928 9628 25956
rect 8588 25900 8616 25928
rect 9600 25900 9628 25928
rect 13173 25925 13185 25959
rect 13219 25956 13231 25959
rect 13262 25956 13268 25968
rect 13219 25928 13268 25956
rect 13219 25925 13231 25928
rect 13173 25919 13231 25925
rect 13262 25916 13268 25928
rect 13320 25916 13326 25968
rect 13814 25916 13820 25968
rect 13872 25956 13878 25968
rect 13872 25928 14596 25956
rect 13872 25916 13878 25928
rect 14568 25900 14596 25928
rect 15470 25916 15476 25968
rect 15528 25916 15534 25968
rect 16022 25916 16028 25968
rect 16080 25956 16086 25968
rect 16301 25959 16359 25965
rect 16301 25956 16313 25959
rect 16080 25928 16313 25956
rect 16080 25916 16086 25928
rect 16301 25925 16313 25928
rect 16347 25925 16359 25959
rect 16301 25919 16359 25925
rect 17218 25916 17224 25968
rect 17276 25916 17282 25968
rect 20530 25916 20536 25968
rect 20588 25956 20594 25968
rect 20717 25959 20775 25965
rect 20717 25956 20729 25959
rect 20588 25928 20729 25956
rect 20588 25916 20594 25928
rect 20717 25925 20729 25928
rect 20763 25925 20775 25959
rect 20717 25919 20775 25925
rect 20898 25916 20904 25968
rect 20956 25965 20962 25968
rect 20956 25959 20975 25965
rect 20963 25925 20975 25959
rect 21100 25956 21128 25984
rect 21100 25928 21404 25956
rect 20956 25919 20975 25925
rect 20956 25916 20962 25919
rect 7101 25891 7159 25897
rect 7101 25888 7113 25891
rect 6656 25860 7113 25888
rect 7101 25857 7113 25860
rect 7147 25857 7159 25891
rect 7101 25851 7159 25857
rect 4433 25823 4491 25829
rect 3344 25792 3648 25820
rect 3620 25752 3648 25792
rect 4433 25789 4445 25823
rect 4479 25789 4491 25823
rect 4433 25783 4491 25789
rect 4525 25823 4583 25829
rect 4525 25789 4537 25823
rect 4571 25820 4583 25823
rect 4571 25792 4752 25820
rect 4571 25789 4583 25792
rect 4525 25783 4583 25789
rect 3878 25752 3884 25764
rect 3620 25724 3884 25752
rect 3878 25712 3884 25724
rect 3936 25712 3942 25764
rect 3973 25755 4031 25761
rect 3973 25721 3985 25755
rect 4019 25752 4031 25755
rect 4448 25752 4476 25783
rect 4614 25752 4620 25764
rect 4019 25724 4620 25752
rect 4019 25721 4031 25724
rect 3973 25715 4031 25721
rect 4614 25712 4620 25724
rect 4672 25712 4678 25764
rect 4724 25752 4752 25792
rect 4798 25780 4804 25832
rect 4856 25820 4862 25832
rect 5353 25823 5411 25829
rect 5353 25820 5365 25823
rect 4856 25792 5365 25820
rect 4856 25780 4862 25792
rect 5353 25789 5365 25792
rect 5399 25789 5411 25823
rect 5353 25783 5411 25789
rect 5537 25823 5595 25829
rect 5537 25789 5549 25823
rect 5583 25820 5595 25823
rect 5994 25820 6000 25832
rect 5583 25792 6000 25820
rect 5583 25789 5595 25792
rect 5537 25783 5595 25789
rect 5994 25780 6000 25792
rect 6052 25780 6058 25832
rect 7116 25820 7144 25851
rect 7190 25848 7196 25900
rect 7248 25888 7254 25900
rect 8113 25891 8171 25897
rect 8113 25888 8125 25891
rect 7248 25860 8125 25888
rect 7248 25848 7254 25860
rect 8113 25857 8125 25860
rect 8159 25857 8171 25891
rect 8113 25851 8171 25857
rect 8202 25848 8208 25900
rect 8260 25848 8266 25900
rect 8297 25891 8355 25897
rect 8297 25857 8309 25891
rect 8343 25888 8355 25891
rect 8386 25888 8392 25900
rect 8343 25860 8392 25888
rect 8343 25857 8355 25860
rect 8297 25851 8355 25857
rect 8312 25820 8340 25851
rect 8386 25848 8392 25860
rect 8444 25848 8450 25900
rect 8481 25891 8539 25897
rect 8481 25857 8493 25891
rect 8527 25888 8539 25891
rect 8570 25888 8576 25900
rect 8527 25860 8576 25888
rect 8527 25857 8539 25860
rect 8481 25851 8539 25857
rect 8570 25848 8576 25860
rect 8628 25848 8634 25900
rect 8754 25848 8760 25900
rect 8812 25848 8818 25900
rect 9398 25848 9404 25900
rect 9456 25888 9462 25900
rect 9493 25891 9551 25897
rect 9493 25888 9505 25891
rect 9456 25860 9505 25888
rect 9456 25848 9462 25860
rect 9493 25857 9505 25860
rect 9539 25857 9551 25891
rect 9493 25851 9551 25857
rect 9582 25848 9588 25900
rect 9640 25848 9646 25900
rect 10962 25848 10968 25900
rect 11020 25888 11026 25900
rect 11149 25891 11207 25897
rect 11149 25888 11161 25891
rect 11020 25860 11161 25888
rect 11020 25848 11026 25860
rect 11149 25857 11161 25860
rect 11195 25857 11207 25891
rect 11149 25851 11207 25857
rect 11333 25891 11391 25897
rect 11333 25857 11345 25891
rect 11379 25888 11391 25891
rect 12069 25891 12127 25897
rect 12069 25888 12081 25891
rect 11379 25860 12081 25888
rect 11379 25857 11391 25860
rect 11333 25851 11391 25857
rect 12069 25857 12081 25860
rect 12115 25857 12127 25891
rect 12069 25851 12127 25857
rect 7116 25792 8340 25820
rect 9309 25823 9367 25829
rect 9309 25789 9321 25823
rect 9355 25789 9367 25823
rect 11164 25820 11192 25851
rect 12710 25848 12716 25900
rect 12768 25848 12774 25900
rect 13538 25848 13544 25900
rect 13596 25848 13602 25900
rect 13630 25848 13636 25900
rect 13688 25848 13694 25900
rect 14277 25891 14335 25897
rect 14277 25857 14289 25891
rect 14323 25888 14335 25891
rect 14366 25888 14372 25900
rect 14323 25860 14372 25888
rect 14323 25857 14335 25860
rect 14277 25851 14335 25857
rect 14366 25848 14372 25860
rect 14424 25848 14430 25900
rect 14550 25848 14556 25900
rect 14608 25848 14614 25900
rect 15746 25848 15752 25900
rect 15804 25848 15810 25900
rect 15933 25891 15991 25897
rect 15933 25857 15945 25891
rect 15979 25857 15991 25891
rect 15933 25851 15991 25857
rect 16393 25891 16451 25897
rect 16393 25857 16405 25891
rect 16439 25888 16451 25891
rect 16850 25888 16856 25900
rect 16439 25860 16856 25888
rect 16439 25857 16451 25860
rect 16393 25851 16451 25857
rect 11164 25792 12848 25820
rect 9309 25783 9367 25789
rect 5258 25752 5264 25764
rect 4724 25724 5264 25752
rect 5258 25712 5264 25724
rect 5316 25712 5322 25764
rect 6178 25712 6184 25764
rect 6236 25752 6242 25764
rect 6546 25752 6552 25764
rect 6236 25724 6552 25752
rect 6236 25712 6242 25724
rect 6546 25712 6552 25724
rect 6604 25752 6610 25764
rect 7466 25752 7472 25764
rect 6604 25724 7472 25752
rect 6604 25712 6610 25724
rect 7466 25712 7472 25724
rect 7524 25712 7530 25764
rect 8294 25712 8300 25764
rect 8352 25752 8358 25764
rect 9324 25752 9352 25783
rect 12820 25761 12848 25792
rect 13078 25780 13084 25832
rect 13136 25820 13142 25832
rect 13265 25823 13323 25829
rect 13265 25820 13277 25823
rect 13136 25792 13277 25820
rect 13136 25780 13142 25792
rect 13265 25789 13277 25792
rect 13311 25820 13323 25823
rect 13354 25820 13360 25832
rect 13311 25792 13360 25820
rect 13311 25789 13323 25792
rect 13265 25783 13323 25789
rect 13354 25780 13360 25792
rect 13412 25780 13418 25832
rect 15948 25820 15976 25851
rect 16850 25848 16856 25860
rect 16908 25848 16914 25900
rect 17129 25891 17187 25897
rect 17129 25857 17141 25891
rect 17175 25888 17187 25891
rect 17236 25888 17264 25916
rect 17175 25860 17264 25888
rect 17175 25857 17187 25860
rect 17129 25851 17187 25857
rect 17310 25848 17316 25900
rect 17368 25848 17374 25900
rect 21376 25897 21404 25928
rect 20625 25891 20683 25897
rect 20625 25857 20637 25891
rect 20671 25888 20683 25891
rect 21177 25891 21235 25897
rect 21177 25888 21189 25891
rect 20671 25860 21189 25888
rect 20671 25857 20683 25860
rect 20625 25851 20683 25857
rect 21177 25857 21189 25860
rect 21223 25857 21235 25891
rect 21177 25851 21235 25857
rect 21361 25891 21419 25897
rect 21361 25857 21373 25891
rect 21407 25857 21419 25891
rect 21361 25851 21419 25857
rect 16482 25820 16488 25832
rect 15948 25792 16488 25820
rect 16482 25780 16488 25792
rect 16540 25780 16546 25832
rect 17037 25823 17095 25829
rect 17037 25789 17049 25823
rect 17083 25789 17095 25823
rect 17037 25783 17095 25789
rect 8352 25724 9352 25752
rect 12805 25755 12863 25761
rect 8352 25712 8358 25724
rect 12805 25721 12817 25755
rect 12851 25721 12863 25755
rect 17052 25752 17080 25783
rect 17218 25780 17224 25832
rect 17276 25780 17282 25832
rect 18141 25823 18199 25829
rect 18141 25789 18153 25823
rect 18187 25789 18199 25823
rect 18141 25783 18199 25789
rect 17589 25755 17647 25761
rect 17589 25752 17601 25755
rect 12805 25715 12863 25721
rect 15948 25724 16574 25752
rect 17052 25724 17601 25752
rect 1673 25687 1731 25693
rect 1673 25653 1685 25687
rect 1719 25684 1731 25687
rect 1762 25684 1768 25696
rect 1719 25656 1768 25684
rect 1719 25653 1731 25656
rect 1673 25647 1731 25653
rect 1762 25644 1768 25656
rect 1820 25644 1826 25696
rect 2777 25687 2835 25693
rect 2777 25653 2789 25687
rect 2823 25684 2835 25687
rect 3694 25684 3700 25696
rect 2823 25656 3700 25684
rect 2823 25653 2835 25656
rect 2777 25647 2835 25653
rect 3694 25644 3700 25656
rect 3752 25684 3758 25696
rect 4890 25684 4896 25696
rect 3752 25656 4896 25684
rect 3752 25644 3758 25656
rect 4890 25644 4896 25656
rect 4948 25644 4954 25696
rect 7374 25644 7380 25696
rect 7432 25644 7438 25696
rect 7837 25687 7895 25693
rect 7837 25653 7849 25687
rect 7883 25684 7895 25687
rect 8018 25684 8024 25696
rect 7883 25656 8024 25684
rect 7883 25653 7895 25656
rect 7837 25647 7895 25653
rect 8018 25644 8024 25656
rect 8076 25644 8082 25696
rect 12986 25644 12992 25696
rect 13044 25644 13050 25696
rect 13170 25644 13176 25696
rect 13228 25684 13234 25696
rect 13357 25687 13415 25693
rect 13357 25684 13369 25687
rect 13228 25656 13369 25684
rect 13228 25644 13234 25656
rect 13357 25653 13369 25656
rect 13403 25653 13415 25687
rect 13357 25647 13415 25653
rect 13446 25644 13452 25696
rect 13504 25644 13510 25696
rect 15948 25693 15976 25724
rect 15933 25687 15991 25693
rect 15933 25653 15945 25687
rect 15979 25653 15991 25687
rect 16546 25684 16574 25724
rect 17589 25721 17601 25724
rect 17635 25721 17647 25755
rect 17589 25715 17647 25721
rect 16942 25684 16948 25696
rect 16546 25656 16948 25684
rect 15933 25647 15991 25653
rect 16942 25644 16948 25656
rect 17000 25684 17006 25696
rect 18156 25684 18184 25783
rect 19978 25780 19984 25832
rect 20036 25780 20042 25832
rect 17000 25656 18184 25684
rect 17000 25644 17006 25656
rect 19334 25644 19340 25696
rect 19392 25684 19398 25696
rect 20806 25684 20812 25696
rect 19392 25656 20812 25684
rect 19392 25644 19398 25656
rect 20806 25644 20812 25656
rect 20864 25684 20870 25696
rect 20901 25687 20959 25693
rect 20901 25684 20913 25687
rect 20864 25656 20913 25684
rect 20864 25644 20870 25656
rect 20901 25653 20913 25656
rect 20947 25653 20959 25687
rect 20901 25647 20959 25653
rect 20990 25644 20996 25696
rect 21048 25684 21054 25696
rect 21177 25687 21235 25693
rect 21177 25684 21189 25687
rect 21048 25656 21189 25684
rect 21048 25644 21054 25656
rect 21177 25653 21189 25656
rect 21223 25653 21235 25687
rect 21177 25647 21235 25653
rect 1104 25594 27876 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 27876 25594
rect 1104 25520 27876 25542
rect 3970 25440 3976 25492
rect 4028 25480 4034 25492
rect 4249 25483 4307 25489
rect 4249 25480 4261 25483
rect 4028 25452 4261 25480
rect 4028 25440 4034 25452
rect 4249 25449 4261 25452
rect 4295 25449 4307 25483
rect 4249 25443 4307 25449
rect 4617 25483 4675 25489
rect 4617 25449 4629 25483
rect 4663 25480 4675 25483
rect 4706 25480 4712 25492
rect 4663 25452 4712 25480
rect 4663 25449 4675 25452
rect 4617 25443 4675 25449
rect 4706 25440 4712 25452
rect 4764 25440 4770 25492
rect 5350 25440 5356 25492
rect 5408 25440 5414 25492
rect 5721 25483 5779 25489
rect 5721 25449 5733 25483
rect 5767 25480 5779 25483
rect 5902 25480 5908 25492
rect 5767 25452 5908 25480
rect 5767 25449 5779 25452
rect 5721 25443 5779 25449
rect 842 25372 848 25424
rect 900 25412 906 25424
rect 1489 25415 1547 25421
rect 1489 25412 1501 25415
rect 900 25384 1501 25412
rect 900 25372 906 25384
rect 1489 25381 1501 25384
rect 1535 25381 1547 25415
rect 1489 25375 1547 25381
rect 4338 25372 4344 25424
rect 4396 25412 4402 25424
rect 5368 25412 5396 25440
rect 4396 25384 5396 25412
rect 4396 25372 4402 25384
rect 1857 25347 1915 25353
rect 1857 25344 1869 25347
rect 1688 25316 1869 25344
rect 1688 25285 1716 25316
rect 1857 25313 1869 25316
rect 1903 25313 1915 25347
rect 5353 25347 5411 25353
rect 5353 25344 5365 25347
rect 1857 25307 1915 25313
rect 2746 25316 5365 25344
rect 1673 25279 1731 25285
rect 1673 25245 1685 25279
rect 1719 25245 1731 25279
rect 1673 25239 1731 25245
rect 1762 25236 1768 25288
rect 1820 25236 1826 25288
rect 1949 25279 2007 25285
rect 1949 25245 1961 25279
rect 1995 25276 2007 25279
rect 2746 25276 2774 25316
rect 5353 25313 5365 25316
rect 5399 25313 5411 25347
rect 5353 25307 5411 25313
rect 1995 25248 2774 25276
rect 1995 25245 2007 25248
rect 1949 25239 2007 25245
rect 3694 25236 3700 25288
rect 3752 25276 3758 25288
rect 3881 25279 3939 25285
rect 3881 25276 3893 25279
rect 3752 25248 3893 25276
rect 3752 25236 3758 25248
rect 3881 25245 3893 25248
rect 3927 25245 3939 25279
rect 3881 25239 3939 25245
rect 3973 25279 4031 25285
rect 3973 25245 3985 25279
rect 4019 25245 4031 25279
rect 3973 25239 4031 25245
rect 3786 25168 3792 25220
rect 3844 25208 3850 25220
rect 3988 25208 4016 25239
rect 4062 25236 4068 25288
rect 4120 25276 4126 25288
rect 4341 25279 4399 25285
rect 4341 25276 4353 25279
rect 4120 25248 4353 25276
rect 4120 25236 4126 25248
rect 4341 25245 4353 25248
rect 4387 25245 4399 25279
rect 4341 25239 4399 25245
rect 4801 25279 4859 25285
rect 4801 25245 4813 25279
rect 4847 25245 4859 25279
rect 4801 25239 4859 25245
rect 4816 25208 4844 25239
rect 4890 25236 4896 25288
rect 4948 25236 4954 25288
rect 4982 25236 4988 25288
rect 5040 25236 5046 25288
rect 5077 25279 5135 25285
rect 5077 25245 5089 25279
rect 5123 25245 5135 25279
rect 5077 25239 5135 25245
rect 5261 25279 5319 25285
rect 5261 25245 5273 25279
rect 5307 25276 5319 25279
rect 5442 25276 5448 25288
rect 5307 25248 5448 25276
rect 5307 25245 5319 25248
rect 5261 25239 5319 25245
rect 3844 25180 4844 25208
rect 5092 25208 5120 25239
rect 5442 25236 5448 25248
rect 5500 25236 5506 25288
rect 5626 25236 5632 25288
rect 5684 25236 5690 25288
rect 5736 25208 5764 25443
rect 5902 25440 5908 25452
rect 5960 25480 5966 25492
rect 6178 25480 6184 25492
rect 5960 25452 6184 25480
rect 5960 25440 5966 25452
rect 6178 25440 6184 25452
rect 6236 25440 6242 25492
rect 13081 25483 13139 25489
rect 13081 25449 13093 25483
rect 13127 25480 13139 25483
rect 13262 25480 13268 25492
rect 13127 25452 13268 25480
rect 13127 25449 13139 25452
rect 13081 25443 13139 25449
rect 5813 25415 5871 25421
rect 5813 25381 5825 25415
rect 5859 25412 5871 25415
rect 7374 25412 7380 25424
rect 5859 25384 7380 25412
rect 5859 25381 5871 25384
rect 5813 25375 5871 25381
rect 7374 25372 7380 25384
rect 7432 25372 7438 25424
rect 7558 25372 7564 25424
rect 7616 25412 7622 25424
rect 8754 25412 8760 25424
rect 7616 25384 8760 25412
rect 7616 25372 7622 25384
rect 8754 25372 8760 25384
rect 8812 25372 8818 25424
rect 6730 25344 6736 25356
rect 6104 25316 6736 25344
rect 5810 25236 5816 25288
rect 5868 25276 5874 25288
rect 6104 25285 6132 25316
rect 6730 25304 6736 25316
rect 6788 25304 6794 25356
rect 6822 25304 6828 25356
rect 6880 25304 6886 25356
rect 7282 25304 7288 25356
rect 7340 25344 7346 25356
rect 7466 25344 7472 25356
rect 7340 25316 7472 25344
rect 7340 25304 7346 25316
rect 7466 25304 7472 25316
rect 7524 25304 7530 25356
rect 7742 25304 7748 25356
rect 7800 25344 7806 25356
rect 8294 25344 8300 25356
rect 7800 25316 8300 25344
rect 7800 25304 7806 25316
rect 8294 25304 8300 25316
rect 8352 25304 8358 25356
rect 9582 25304 9588 25356
rect 9640 25344 9646 25356
rect 9677 25347 9735 25353
rect 9677 25344 9689 25347
rect 9640 25316 9689 25344
rect 9640 25304 9646 25316
rect 9677 25313 9689 25316
rect 9723 25313 9735 25347
rect 9677 25307 9735 25313
rect 11606 25304 11612 25356
rect 11664 25344 11670 25356
rect 13188 25353 13216 25452
rect 13262 25440 13268 25452
rect 13320 25440 13326 25492
rect 15930 25440 15936 25492
rect 15988 25480 15994 25492
rect 16301 25483 16359 25489
rect 16301 25480 16313 25483
rect 15988 25452 16313 25480
rect 15988 25440 15994 25452
rect 16301 25449 16313 25452
rect 16347 25449 16359 25483
rect 16301 25443 16359 25449
rect 19613 25483 19671 25489
rect 19613 25449 19625 25483
rect 19659 25480 19671 25483
rect 19978 25480 19984 25492
rect 19659 25452 19984 25480
rect 19659 25449 19671 25452
rect 19613 25443 19671 25449
rect 19978 25440 19984 25452
rect 20036 25440 20042 25492
rect 20898 25440 20904 25492
rect 20956 25480 20962 25492
rect 21085 25483 21143 25489
rect 21085 25480 21097 25483
rect 20956 25452 21097 25480
rect 20956 25440 20962 25452
rect 21085 25449 21097 25452
rect 21131 25449 21143 25483
rect 21085 25443 21143 25449
rect 11701 25347 11759 25353
rect 11701 25344 11713 25347
rect 11664 25316 11713 25344
rect 11664 25304 11670 25316
rect 11701 25313 11713 25316
rect 11747 25313 11759 25347
rect 11701 25307 11759 25313
rect 13173 25347 13231 25353
rect 13173 25313 13185 25347
rect 13219 25313 13231 25347
rect 13173 25307 13231 25313
rect 18598 25304 18604 25356
rect 18656 25344 18662 25356
rect 19705 25347 19763 25353
rect 19705 25344 19717 25347
rect 18656 25316 19717 25344
rect 18656 25304 18662 25316
rect 19705 25313 19717 25316
rect 19751 25313 19763 25347
rect 21100 25344 21128 25443
rect 21729 25347 21787 25353
rect 21729 25344 21741 25347
rect 21100 25316 21741 25344
rect 19705 25307 19763 25313
rect 21729 25313 21741 25316
rect 21775 25313 21787 25347
rect 21729 25307 21787 25313
rect 5905 25279 5963 25285
rect 5905 25276 5917 25279
rect 5868 25248 5917 25276
rect 5868 25236 5874 25248
rect 5905 25245 5917 25248
rect 5951 25245 5963 25279
rect 5905 25239 5963 25245
rect 6089 25279 6147 25285
rect 6089 25245 6101 25279
rect 6135 25245 6147 25279
rect 6089 25239 6147 25245
rect 5092 25180 5764 25208
rect 5920 25208 5948 25239
rect 6178 25236 6184 25288
rect 6236 25276 6242 25288
rect 6365 25279 6423 25285
rect 6365 25276 6377 25279
rect 6236 25248 6377 25276
rect 6236 25236 6242 25248
rect 6365 25245 6377 25248
rect 6411 25245 6423 25279
rect 6365 25239 6423 25245
rect 6457 25279 6515 25285
rect 6457 25245 6469 25279
rect 6503 25276 6515 25279
rect 6914 25276 6920 25288
rect 6503 25248 6920 25276
rect 6503 25245 6515 25248
rect 6457 25239 6515 25245
rect 6914 25236 6920 25248
rect 6972 25236 6978 25288
rect 8113 25279 8171 25285
rect 8113 25245 8125 25279
rect 8159 25276 8171 25279
rect 8202 25276 8208 25288
rect 8159 25248 8208 25276
rect 8159 25245 8171 25248
rect 8113 25239 8171 25245
rect 8202 25236 8208 25248
rect 8260 25236 8266 25288
rect 10042 25236 10048 25288
rect 10100 25276 10106 25288
rect 10137 25279 10195 25285
rect 10137 25276 10149 25279
rect 10100 25248 10149 25276
rect 10100 25236 10106 25248
rect 10137 25245 10149 25248
rect 10183 25245 10195 25279
rect 10137 25239 10195 25245
rect 14550 25236 14556 25288
rect 14608 25276 14614 25288
rect 14918 25276 14924 25288
rect 14608 25248 14924 25276
rect 14608 25236 14614 25248
rect 14918 25236 14924 25248
rect 14976 25276 14982 25288
rect 15565 25279 15623 25285
rect 15565 25276 15577 25279
rect 14976 25248 15577 25276
rect 14976 25236 14982 25248
rect 15565 25245 15577 25248
rect 15611 25245 15623 25279
rect 15565 25239 15623 25245
rect 10404 25211 10462 25217
rect 5920 25180 6592 25208
rect 3844 25168 3850 25180
rect 4525 25143 4583 25149
rect 4525 25109 4537 25143
rect 4571 25140 4583 25143
rect 4706 25140 4712 25152
rect 4571 25112 4712 25140
rect 4571 25109 4583 25112
rect 4525 25103 4583 25109
rect 4706 25100 4712 25112
rect 4764 25100 4770 25152
rect 5350 25100 5356 25152
rect 5408 25140 5414 25152
rect 6564 25149 6592 25180
rect 10404 25177 10416 25211
rect 10450 25208 10462 25211
rect 10962 25208 10968 25220
rect 10450 25180 10968 25208
rect 10450 25177 10462 25180
rect 10404 25171 10462 25177
rect 10962 25168 10968 25180
rect 11020 25168 11026 25220
rect 11968 25211 12026 25217
rect 11968 25177 11980 25211
rect 12014 25208 12026 25211
rect 12434 25208 12440 25220
rect 12014 25180 12440 25208
rect 12014 25177 12026 25180
rect 11968 25171 12026 25177
rect 12434 25168 12440 25180
rect 12492 25168 12498 25220
rect 6181 25143 6239 25149
rect 6181 25140 6193 25143
rect 5408 25112 6193 25140
rect 5408 25100 5414 25112
rect 6181 25109 6193 25112
rect 6227 25109 6239 25143
rect 6181 25103 6239 25109
rect 6549 25143 6607 25149
rect 6549 25109 6561 25143
rect 6595 25140 6607 25143
rect 6730 25140 6736 25152
rect 6595 25112 6736 25140
rect 6595 25109 6607 25112
rect 6549 25103 6607 25109
rect 6730 25100 6736 25112
rect 6788 25100 6794 25152
rect 7926 25100 7932 25152
rect 7984 25100 7990 25152
rect 8205 25143 8263 25149
rect 8205 25109 8217 25143
rect 8251 25140 8263 25143
rect 8294 25140 8300 25152
rect 8251 25112 8300 25140
rect 8251 25109 8263 25112
rect 8205 25103 8263 25109
rect 8294 25100 8300 25112
rect 8352 25100 8358 25152
rect 8478 25100 8484 25152
rect 8536 25140 8542 25152
rect 9125 25143 9183 25149
rect 9125 25140 9137 25143
rect 8536 25112 9137 25140
rect 8536 25100 8542 25112
rect 9125 25109 9137 25112
rect 9171 25140 9183 25143
rect 9306 25140 9312 25152
rect 9171 25112 9312 25140
rect 9171 25109 9183 25112
rect 9125 25103 9183 25109
rect 9306 25100 9312 25112
rect 9364 25100 9370 25152
rect 10502 25100 10508 25152
rect 10560 25140 10566 25152
rect 11517 25143 11575 25149
rect 11517 25140 11529 25143
rect 10560 25112 11529 25140
rect 10560 25100 10566 25112
rect 11517 25109 11529 25112
rect 11563 25109 11575 25143
rect 11517 25103 11575 25109
rect 12618 25100 12624 25152
rect 12676 25140 12682 25152
rect 13538 25140 13544 25152
rect 12676 25112 13544 25140
rect 12676 25100 12682 25112
rect 13538 25100 13544 25112
rect 13596 25140 13602 25152
rect 13817 25143 13875 25149
rect 13817 25140 13829 25143
rect 13596 25112 13829 25140
rect 13596 25100 13602 25112
rect 13817 25109 13829 25112
rect 13863 25109 13875 25143
rect 13817 25103 13875 25109
rect 15470 25100 15476 25152
rect 15528 25100 15534 25152
rect 15580 25140 15608 25239
rect 19334 25236 19340 25288
rect 19392 25236 19398 25288
rect 19613 25279 19671 25285
rect 19613 25245 19625 25279
rect 19659 25276 19671 25279
rect 21177 25279 21235 25285
rect 21177 25276 21189 25279
rect 19659 25248 21189 25276
rect 19659 25245 19671 25248
rect 19613 25239 19671 25245
rect 21177 25245 21189 25248
rect 21223 25245 21235 25279
rect 21177 25239 21235 25245
rect 16482 25168 16488 25220
rect 16540 25168 16546 25220
rect 19972 25211 20030 25217
rect 19972 25177 19984 25211
rect 20018 25208 20030 25211
rect 20990 25208 20996 25220
rect 20018 25180 20996 25208
rect 20018 25177 20030 25180
rect 19972 25171 20030 25177
rect 20990 25168 20996 25180
rect 21048 25168 21054 25220
rect 16117 25143 16175 25149
rect 16117 25140 16129 25143
rect 15580 25112 16129 25140
rect 16117 25109 16129 25112
rect 16163 25109 16175 25143
rect 16117 25103 16175 25109
rect 16285 25143 16343 25149
rect 16285 25109 16297 25143
rect 16331 25140 16343 25143
rect 16666 25140 16672 25152
rect 16331 25112 16672 25140
rect 16331 25109 16343 25112
rect 16285 25103 16343 25109
rect 16666 25100 16672 25112
rect 16724 25100 16730 25152
rect 19429 25143 19487 25149
rect 19429 25109 19441 25143
rect 19475 25140 19487 25143
rect 20530 25140 20536 25152
rect 19475 25112 20536 25140
rect 19475 25109 19487 25112
rect 19429 25103 19487 25109
rect 20530 25100 20536 25112
rect 20588 25100 20594 25152
rect 1104 25050 27876 25072
rect 1104 24998 4874 25050
rect 4926 24998 4938 25050
rect 4990 24998 5002 25050
rect 5054 24998 5066 25050
rect 5118 24998 5130 25050
rect 5182 24998 27876 25050
rect 1104 24976 27876 24998
rect 2685 24939 2743 24945
rect 2685 24905 2697 24939
rect 2731 24905 2743 24939
rect 2685 24899 2743 24905
rect 1946 24828 1952 24880
rect 2004 24868 2010 24880
rect 2700 24868 2728 24899
rect 6454 24896 6460 24948
rect 6512 24936 6518 24948
rect 6822 24936 6828 24948
rect 6512 24908 6828 24936
rect 6512 24896 6518 24908
rect 6822 24896 6828 24908
rect 6880 24936 6886 24948
rect 7653 24939 7711 24945
rect 7653 24936 7665 24939
rect 6880 24908 7665 24936
rect 6880 24896 6886 24908
rect 7653 24905 7665 24908
rect 7699 24905 7711 24939
rect 8665 24939 8723 24945
rect 8665 24936 8677 24939
rect 7653 24899 7711 24905
rect 8312 24908 8677 24936
rect 2866 24877 2872 24880
rect 2004 24840 2728 24868
rect 2853 24871 2872 24877
rect 2004 24828 2010 24840
rect 2853 24837 2865 24871
rect 2853 24831 2872 24837
rect 2866 24828 2872 24831
rect 2924 24828 2930 24880
rect 3053 24871 3111 24877
rect 3053 24837 3065 24871
rect 3099 24868 3111 24871
rect 3142 24868 3148 24880
rect 3099 24840 3148 24868
rect 3099 24837 3111 24840
rect 3053 24831 3111 24837
rect 3142 24828 3148 24840
rect 3200 24868 3206 24880
rect 3694 24868 3700 24880
rect 3200 24840 3700 24868
rect 3200 24828 3206 24840
rect 3694 24828 3700 24840
rect 3752 24828 3758 24880
rect 5537 24871 5595 24877
rect 4356 24840 5396 24868
rect 1673 24803 1731 24809
rect 1673 24769 1685 24803
rect 1719 24769 1731 24803
rect 1673 24763 1731 24769
rect 1857 24803 1915 24809
rect 1857 24769 1869 24803
rect 1903 24800 1915 24803
rect 1964 24800 1992 24828
rect 1903 24772 1992 24800
rect 2041 24803 2099 24809
rect 1903 24769 1915 24772
rect 1857 24763 1915 24769
rect 2041 24769 2053 24803
rect 2087 24800 2099 24803
rect 2958 24800 2964 24812
rect 2087 24772 2964 24800
rect 2087 24769 2099 24772
rect 2041 24763 2099 24769
rect 1688 24732 1716 24763
rect 2958 24760 2964 24772
rect 3016 24760 3022 24812
rect 4065 24803 4123 24809
rect 4065 24769 4077 24803
rect 4111 24800 4123 24803
rect 4356 24800 4384 24840
rect 5368 24812 5396 24840
rect 5537 24837 5549 24871
rect 5583 24868 5595 24871
rect 7668 24868 7696 24899
rect 8110 24868 8116 24880
rect 5583 24840 7420 24868
rect 7668 24840 8116 24868
rect 5583 24837 5595 24840
rect 5537 24831 5595 24837
rect 7392 24812 7420 24840
rect 8110 24828 8116 24840
rect 8168 24828 8174 24880
rect 4111 24772 4384 24800
rect 4433 24803 4491 24809
rect 4111 24769 4123 24772
rect 4065 24763 4123 24769
rect 4433 24769 4445 24803
rect 4479 24800 4491 24803
rect 4522 24800 4528 24812
rect 4479 24772 4528 24800
rect 4479 24769 4491 24772
rect 4433 24763 4491 24769
rect 4522 24760 4528 24772
rect 4580 24760 4586 24812
rect 4617 24803 4675 24809
rect 4617 24769 4629 24803
rect 4663 24769 4675 24803
rect 4617 24763 4675 24769
rect 1688 24704 4016 24732
rect 842 24624 848 24676
rect 900 24664 906 24676
rect 1489 24667 1547 24673
rect 1489 24664 1501 24667
rect 900 24636 1501 24664
rect 900 24624 906 24636
rect 1489 24633 1501 24636
rect 1535 24633 1547 24667
rect 3881 24667 3939 24673
rect 3881 24664 3893 24667
rect 1489 24627 1547 24633
rect 2746 24636 3893 24664
rect 2038 24556 2044 24608
rect 2096 24556 2102 24608
rect 2222 24556 2228 24608
rect 2280 24596 2286 24608
rect 2746 24596 2774 24636
rect 3881 24633 3893 24636
rect 3927 24633 3939 24667
rect 3988 24664 4016 24704
rect 4338 24692 4344 24744
rect 4396 24692 4402 24744
rect 4632 24732 4660 24763
rect 5350 24760 5356 24812
rect 5408 24760 5414 24812
rect 5629 24803 5687 24809
rect 5629 24769 5641 24803
rect 5675 24769 5687 24803
rect 5629 24763 5687 24769
rect 4706 24732 4712 24744
rect 4632 24704 4712 24732
rect 4706 24692 4712 24704
rect 4764 24732 4770 24744
rect 5442 24732 5448 24744
rect 4764 24704 5448 24732
rect 4764 24692 4770 24704
rect 5442 24692 5448 24704
rect 5500 24692 5506 24744
rect 5644 24732 5672 24763
rect 5810 24760 5816 24812
rect 5868 24760 5874 24812
rect 5997 24803 6055 24809
rect 5997 24769 6009 24803
rect 6043 24800 6055 24803
rect 6270 24800 6276 24812
rect 6043 24772 6276 24800
rect 6043 24769 6055 24772
rect 5997 24763 6055 24769
rect 6270 24760 6276 24772
rect 6328 24760 6334 24812
rect 6362 24760 6368 24812
rect 6420 24760 6426 24812
rect 6546 24760 6552 24812
rect 6604 24760 6610 24812
rect 6730 24760 6736 24812
rect 6788 24760 6794 24812
rect 6822 24760 6828 24812
rect 6880 24760 6886 24812
rect 6914 24760 6920 24812
rect 6972 24800 6978 24812
rect 7285 24803 7343 24809
rect 7285 24800 7297 24803
rect 6972 24772 7297 24800
rect 6972 24760 6978 24772
rect 7285 24769 7297 24772
rect 7331 24769 7343 24803
rect 7285 24763 7343 24769
rect 7374 24760 7380 24812
rect 7432 24800 7438 24812
rect 7469 24803 7527 24809
rect 7469 24800 7481 24803
rect 7432 24772 7481 24800
rect 7432 24760 7438 24772
rect 7469 24769 7481 24772
rect 7515 24769 7527 24803
rect 7469 24763 7527 24769
rect 7558 24760 7564 24812
rect 7616 24760 7622 24812
rect 7742 24760 7748 24812
rect 7800 24800 7806 24812
rect 7837 24803 7895 24809
rect 7837 24800 7849 24803
rect 7800 24772 7849 24800
rect 7800 24760 7806 24772
rect 7837 24769 7849 24772
rect 7883 24769 7895 24803
rect 7837 24763 7895 24769
rect 8018 24760 8024 24812
rect 8076 24760 8082 24812
rect 8128 24800 8156 24828
rect 8205 24803 8263 24809
rect 8205 24800 8217 24803
rect 8128 24772 8217 24800
rect 8205 24769 8217 24772
rect 8251 24769 8263 24803
rect 8205 24763 8263 24769
rect 5905 24735 5963 24741
rect 5905 24732 5917 24735
rect 5644 24704 5917 24732
rect 5905 24701 5917 24704
rect 5951 24701 5963 24735
rect 6288 24732 6316 24760
rect 8113 24735 8171 24741
rect 8113 24732 8125 24735
rect 6288 24704 7604 24732
rect 5905 24695 5963 24701
rect 4798 24664 4804 24676
rect 3988 24636 4804 24664
rect 3881 24627 3939 24633
rect 4798 24624 4804 24636
rect 4856 24624 4862 24676
rect 5258 24624 5264 24676
rect 5316 24664 5322 24676
rect 5353 24667 5411 24673
rect 5353 24664 5365 24667
rect 5316 24636 5365 24664
rect 5316 24624 5322 24636
rect 5353 24633 5365 24636
rect 5399 24633 5411 24667
rect 5353 24627 5411 24633
rect 5810 24624 5816 24676
rect 5868 24664 5874 24676
rect 6546 24664 6552 24676
rect 5868 24636 6552 24664
rect 5868 24624 5874 24636
rect 6546 24624 6552 24636
rect 6604 24664 6610 24676
rect 6822 24664 6828 24676
rect 6604 24636 6828 24664
rect 6604 24624 6610 24636
rect 6822 24624 6828 24636
rect 6880 24624 6886 24676
rect 7576 24664 7604 24704
rect 7751 24704 8125 24732
rect 7751 24664 7779 24704
rect 8113 24701 8125 24704
rect 8159 24732 8171 24735
rect 8312 24732 8340 24908
rect 8665 24905 8677 24908
rect 8711 24905 8723 24939
rect 8665 24899 8723 24905
rect 15930 24896 15936 24948
rect 15988 24936 15994 24948
rect 16485 24939 16543 24945
rect 16485 24936 16497 24939
rect 15988 24908 16497 24936
rect 15988 24896 15994 24908
rect 16485 24905 16497 24908
rect 16531 24905 16543 24939
rect 16485 24899 16543 24905
rect 19981 24939 20039 24945
rect 19981 24905 19993 24939
rect 20027 24936 20039 24939
rect 20530 24936 20536 24948
rect 20027 24908 20536 24936
rect 20027 24905 20039 24908
rect 19981 24899 20039 24905
rect 20530 24896 20536 24908
rect 20588 24896 20594 24948
rect 8386 24760 8392 24812
rect 8444 24760 8450 24812
rect 8573 24803 8631 24809
rect 8573 24769 8585 24803
rect 8619 24800 8631 24803
rect 9778 24803 9836 24809
rect 9778 24800 9790 24803
rect 8619 24772 9790 24800
rect 8619 24769 8631 24772
rect 8573 24763 8631 24769
rect 9778 24769 9790 24772
rect 9824 24769 9836 24803
rect 9778 24763 9836 24769
rect 9950 24760 9956 24812
rect 10008 24800 10014 24812
rect 10229 24803 10287 24809
rect 10229 24800 10241 24803
rect 10008 24772 10241 24800
rect 10008 24760 10014 24772
rect 10229 24769 10241 24772
rect 10275 24769 10287 24803
rect 10229 24763 10287 24769
rect 10318 24760 10324 24812
rect 10376 24800 10382 24812
rect 10413 24803 10471 24809
rect 10413 24800 10425 24803
rect 10376 24772 10425 24800
rect 10376 24760 10382 24772
rect 10413 24769 10425 24772
rect 10459 24800 10471 24803
rect 10502 24800 10508 24812
rect 10459 24772 10508 24800
rect 10459 24769 10471 24772
rect 10413 24763 10471 24769
rect 10502 24760 10508 24772
rect 10560 24760 10566 24812
rect 12713 24803 12771 24809
rect 12713 24769 12725 24803
rect 12759 24769 12771 24803
rect 12713 24763 12771 24769
rect 14645 24803 14703 24809
rect 14645 24769 14657 24803
rect 14691 24800 14703 24803
rect 15010 24800 15016 24812
rect 14691 24772 15016 24800
rect 14691 24769 14703 24772
rect 14645 24763 14703 24769
rect 8159 24704 8340 24732
rect 8159 24701 8171 24704
rect 8113 24695 8171 24701
rect 10042 24692 10048 24744
rect 10100 24692 10106 24744
rect 10778 24692 10784 24744
rect 10836 24732 10842 24744
rect 11517 24735 11575 24741
rect 11517 24732 11529 24735
rect 10836 24704 11529 24732
rect 10836 24692 10842 24704
rect 11517 24701 11529 24704
rect 11563 24701 11575 24735
rect 11517 24695 11575 24701
rect 11606 24692 11612 24744
rect 11664 24732 11670 24744
rect 12342 24732 12348 24744
rect 11664 24704 12348 24732
rect 11664 24692 11670 24704
rect 12342 24692 12348 24704
rect 12400 24732 12406 24744
rect 12728 24732 12756 24763
rect 15010 24760 15016 24772
rect 15068 24760 15074 24812
rect 15378 24809 15384 24812
rect 15372 24763 15384 24809
rect 15378 24760 15384 24763
rect 15436 24760 15442 24812
rect 16850 24760 16856 24812
rect 16908 24800 16914 24812
rect 18242 24803 18300 24809
rect 18242 24800 18254 24803
rect 16908 24772 18254 24800
rect 16908 24760 16914 24772
rect 18242 24769 18254 24772
rect 18288 24769 18300 24803
rect 18242 24763 18300 24769
rect 18509 24803 18567 24809
rect 18509 24769 18521 24803
rect 18555 24800 18567 24803
rect 18598 24800 18604 24812
rect 18555 24772 18604 24800
rect 18555 24769 18567 24772
rect 18509 24763 18567 24769
rect 18598 24760 18604 24772
rect 18656 24760 18662 24812
rect 18690 24760 18696 24812
rect 18748 24800 18754 24812
rect 18857 24803 18915 24809
rect 18857 24800 18869 24803
rect 18748 24772 18869 24800
rect 18748 24760 18754 24772
rect 18857 24769 18869 24772
rect 18903 24769 18915 24803
rect 18857 24763 18915 24769
rect 20530 24760 20536 24812
rect 20588 24800 20594 24812
rect 20625 24803 20683 24809
rect 20625 24800 20637 24803
rect 20588 24772 20637 24800
rect 20588 24760 20594 24772
rect 20625 24769 20637 24772
rect 20671 24769 20683 24803
rect 20625 24763 20683 24769
rect 15105 24735 15163 24741
rect 15105 24732 15117 24735
rect 12400 24704 15117 24732
rect 12400 24692 12406 24704
rect 13372 24673 13400 24704
rect 15105 24701 15117 24704
rect 15151 24701 15163 24735
rect 15105 24695 15163 24701
rect 7576 24636 7779 24664
rect 13357 24667 13415 24673
rect 13357 24633 13369 24667
rect 13403 24633 13415 24667
rect 13357 24627 13415 24633
rect 16482 24624 16488 24676
rect 16540 24664 16546 24676
rect 17129 24667 17187 24673
rect 17129 24664 17141 24667
rect 16540 24636 17141 24664
rect 16540 24624 16546 24636
rect 17129 24633 17141 24636
rect 17175 24633 17187 24667
rect 17129 24627 17187 24633
rect 2280 24568 2774 24596
rect 2869 24599 2927 24605
rect 2280 24556 2286 24568
rect 2869 24565 2881 24599
rect 2915 24596 2927 24599
rect 3418 24596 3424 24608
rect 2915 24568 3424 24596
rect 2915 24565 2927 24568
rect 2869 24559 2927 24565
rect 3418 24556 3424 24568
rect 3476 24596 3482 24608
rect 3970 24596 3976 24608
rect 3476 24568 3976 24596
rect 3476 24556 3482 24568
rect 3970 24556 3976 24568
rect 4028 24556 4034 24608
rect 4249 24599 4307 24605
rect 4249 24565 4261 24599
rect 4295 24596 4307 24599
rect 4525 24599 4583 24605
rect 4525 24596 4537 24599
rect 4295 24568 4537 24596
rect 4295 24565 4307 24568
rect 4249 24559 4307 24565
rect 4525 24565 4537 24568
rect 4571 24565 4583 24599
rect 4525 24559 4583 24565
rect 7098 24556 7104 24608
rect 7156 24556 7162 24608
rect 7377 24599 7435 24605
rect 7377 24565 7389 24599
rect 7423 24596 7435 24599
rect 8386 24596 8392 24608
rect 7423 24568 8392 24596
rect 7423 24565 7435 24568
rect 7377 24559 7435 24565
rect 8386 24556 8392 24568
rect 8444 24556 8450 24608
rect 10321 24599 10379 24605
rect 10321 24565 10333 24599
rect 10367 24596 10379 24599
rect 10410 24596 10416 24608
rect 10367 24568 10416 24596
rect 10367 24565 10379 24568
rect 10321 24559 10379 24565
rect 10410 24556 10416 24568
rect 10468 24556 10474 24608
rect 12066 24556 12072 24608
rect 12124 24596 12130 24608
rect 12161 24599 12219 24605
rect 12161 24596 12173 24599
rect 12124 24568 12173 24596
rect 12124 24556 12130 24568
rect 12161 24565 12173 24568
rect 12207 24565 12219 24599
rect 12161 24559 12219 24565
rect 20070 24556 20076 24608
rect 20128 24556 20134 24608
rect 1104 24506 27876 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 27876 24506
rect 1104 24432 27876 24454
rect 2958 24352 2964 24404
rect 3016 24352 3022 24404
rect 3418 24352 3424 24404
rect 3476 24352 3482 24404
rect 7834 24352 7840 24404
rect 7892 24392 7898 24404
rect 8021 24395 8079 24401
rect 8021 24392 8033 24395
rect 7892 24364 8033 24392
rect 7892 24352 7898 24364
rect 2777 24327 2835 24333
rect 2777 24293 2789 24327
rect 2823 24324 2835 24327
rect 3142 24324 3148 24336
rect 2823 24296 3148 24324
rect 2823 24293 2835 24296
rect 2777 24287 2835 24293
rect 3142 24284 3148 24296
rect 3200 24284 3206 24336
rect 5442 24284 5448 24336
rect 5500 24324 5506 24336
rect 5500 24296 6592 24324
rect 5500 24284 5506 24296
rect 1394 24216 1400 24268
rect 1452 24216 1458 24268
rect 2869 24259 2927 24265
rect 2869 24256 2881 24259
rect 2700 24228 2881 24256
rect 1664 24191 1722 24197
rect 1664 24157 1676 24191
rect 1710 24188 1722 24191
rect 2038 24188 2044 24200
rect 1710 24160 2044 24188
rect 1710 24157 1722 24160
rect 1664 24151 1722 24157
rect 2038 24148 2044 24160
rect 2096 24148 2102 24200
rect 2700 24120 2728 24228
rect 2869 24225 2881 24228
rect 2915 24225 2927 24259
rect 2869 24219 2927 24225
rect 2774 24148 2780 24200
rect 2832 24188 2838 24200
rect 3160 24197 3188 24284
rect 6362 24216 6368 24268
rect 6420 24216 6426 24268
rect 6454 24216 6460 24268
rect 6512 24216 6518 24268
rect 6564 24265 6592 24296
rect 6549 24259 6607 24265
rect 6549 24225 6561 24259
rect 6595 24225 6607 24259
rect 6549 24219 6607 24225
rect 3053 24191 3111 24197
rect 3053 24188 3065 24191
rect 2832 24160 3065 24188
rect 2832 24148 2838 24160
rect 3053 24157 3065 24160
rect 3099 24157 3111 24191
rect 3053 24151 3111 24157
rect 3145 24191 3203 24197
rect 3145 24157 3157 24191
rect 3191 24157 3203 24191
rect 3145 24151 3203 24157
rect 3234 24148 3240 24200
rect 3292 24188 3298 24200
rect 3329 24191 3387 24197
rect 3329 24188 3341 24191
rect 3292 24160 3341 24188
rect 3292 24148 3298 24160
rect 3329 24157 3341 24160
rect 3375 24157 3387 24191
rect 3329 24151 3387 24157
rect 5997 24191 6055 24197
rect 5997 24157 6009 24191
rect 6043 24157 6055 24191
rect 5997 24151 6055 24157
rect 6641 24191 6699 24197
rect 6641 24157 6653 24191
rect 6687 24188 6699 24191
rect 6730 24188 6736 24200
rect 6687 24160 6736 24188
rect 6687 24157 6699 24160
rect 6641 24151 6699 24157
rect 6012 24120 6040 24151
rect 6730 24148 6736 24160
rect 6788 24148 6794 24200
rect 6822 24148 6828 24200
rect 6880 24148 6886 24200
rect 6914 24148 6920 24200
rect 6972 24188 6978 24200
rect 7944 24197 7972 24364
rect 8021 24361 8033 24364
rect 8067 24361 8079 24395
rect 8021 24355 8079 24361
rect 8294 24352 8300 24404
rect 8352 24352 8358 24404
rect 12434 24352 12440 24404
rect 12492 24352 12498 24404
rect 16850 24352 16856 24404
rect 16908 24352 16914 24404
rect 18690 24352 18696 24404
rect 18748 24352 18754 24404
rect 20806 24352 20812 24404
rect 20864 24392 20870 24404
rect 21085 24395 21143 24401
rect 21085 24392 21097 24395
rect 20864 24364 21097 24392
rect 20864 24352 20870 24364
rect 21085 24361 21097 24364
rect 21131 24361 21143 24395
rect 21085 24355 21143 24361
rect 16482 24284 16488 24336
rect 16540 24324 16546 24336
rect 16540 24296 17540 24324
rect 16540 24284 16546 24296
rect 8110 24216 8116 24268
rect 8168 24256 8174 24268
rect 8168 24228 8432 24256
rect 8168 24216 8174 24228
rect 7745 24191 7803 24197
rect 7745 24188 7757 24191
rect 6972 24160 7757 24188
rect 6972 24148 6978 24160
rect 7745 24157 7757 24160
rect 7791 24157 7803 24191
rect 7745 24151 7803 24157
rect 7929 24191 7987 24197
rect 7929 24157 7941 24191
rect 7975 24157 7987 24191
rect 7929 24151 7987 24157
rect 8294 24148 8300 24200
rect 8352 24148 8358 24200
rect 8404 24197 8432 24228
rect 12342 24216 12348 24268
rect 12400 24216 12406 24268
rect 13446 24256 13452 24268
rect 12728 24228 13452 24256
rect 8389 24191 8447 24197
rect 8389 24157 8401 24191
rect 8435 24157 8447 24191
rect 8389 24151 8447 24157
rect 8665 24191 8723 24197
rect 8665 24157 8677 24191
rect 8711 24188 8723 24191
rect 8846 24188 8852 24200
rect 8711 24160 8852 24188
rect 8711 24157 8723 24160
rect 8665 24151 8723 24157
rect 8846 24148 8852 24160
rect 8904 24188 8910 24200
rect 8904 24160 9444 24188
rect 8904 24148 8910 24160
rect 7098 24120 7104 24132
rect 2700 24092 5948 24120
rect 6012 24092 7104 24120
rect 3068 24064 3096 24092
rect 3050 24012 3056 24064
rect 3108 24012 3114 24064
rect 3970 24012 3976 24064
rect 4028 24052 4034 24064
rect 5813 24055 5871 24061
rect 5813 24052 5825 24055
rect 4028 24024 5825 24052
rect 4028 24012 4034 24024
rect 5813 24021 5825 24024
rect 5859 24021 5871 24055
rect 5920 24052 5948 24092
rect 7098 24080 7104 24092
rect 7156 24080 7162 24132
rect 8938 24080 8944 24132
rect 8996 24080 9002 24132
rect 9416 24064 9444 24160
rect 12066 24148 12072 24200
rect 12124 24197 12130 24200
rect 12124 24188 12136 24197
rect 12124 24160 12169 24188
rect 12124 24151 12136 24160
rect 12124 24148 12130 24151
rect 12618 24148 12624 24200
rect 12676 24148 12682 24200
rect 12728 24197 12756 24228
rect 13446 24216 13452 24228
rect 13504 24216 13510 24268
rect 16393 24259 16451 24265
rect 16393 24225 16405 24259
rect 16439 24256 16451 24259
rect 16666 24256 16672 24268
rect 16439 24228 16672 24256
rect 16439 24225 16451 24228
rect 16393 24219 16451 24225
rect 16666 24216 16672 24228
rect 16724 24216 16730 24268
rect 17512 24265 17540 24296
rect 17497 24259 17555 24265
rect 17497 24225 17509 24259
rect 17543 24225 17555 24259
rect 17497 24219 17555 24225
rect 18598 24216 18604 24268
rect 18656 24256 18662 24268
rect 19242 24256 19248 24268
rect 18656 24228 19248 24256
rect 18656 24216 18662 24228
rect 19242 24216 19248 24228
rect 19300 24256 19306 24268
rect 19705 24259 19763 24265
rect 19705 24256 19717 24259
rect 19300 24228 19717 24256
rect 19300 24216 19306 24228
rect 19705 24225 19717 24228
rect 19751 24225 19763 24259
rect 21100 24256 21128 24355
rect 21729 24259 21787 24265
rect 21729 24256 21741 24259
rect 21100 24228 21741 24256
rect 19705 24219 19763 24225
rect 21729 24225 21741 24228
rect 21775 24225 21787 24259
rect 21729 24219 21787 24225
rect 12713 24191 12771 24197
rect 12713 24157 12725 24191
rect 12759 24157 12771 24191
rect 12713 24151 12771 24157
rect 12802 24148 12808 24200
rect 12860 24148 12866 24200
rect 12986 24148 12992 24200
rect 13044 24148 13050 24200
rect 13078 24148 13084 24200
rect 13136 24148 13142 24200
rect 13541 24191 13599 24197
rect 13541 24157 13553 24191
rect 13587 24188 13599 24191
rect 13814 24188 13820 24200
rect 13587 24160 13820 24188
rect 13587 24157 13599 24160
rect 13541 24151 13599 24157
rect 13814 24148 13820 24160
rect 13872 24148 13878 24200
rect 14093 24191 14151 24197
rect 14093 24157 14105 24191
rect 14139 24188 14151 24191
rect 15194 24188 15200 24200
rect 14139 24160 15200 24188
rect 14139 24157 14151 24160
rect 14093 24151 14151 24157
rect 15194 24148 15200 24160
rect 15252 24148 15258 24200
rect 16117 24191 16175 24197
rect 16117 24188 16129 24191
rect 15488 24160 16129 24188
rect 12437 24123 12495 24129
rect 12437 24089 12449 24123
rect 12483 24120 12495 24123
rect 13170 24120 13176 24132
rect 12483 24092 13176 24120
rect 12483 24089 12495 24092
rect 12437 24083 12495 24089
rect 13170 24080 13176 24092
rect 13228 24080 13234 24132
rect 14360 24123 14418 24129
rect 14360 24089 14372 24123
rect 14406 24120 14418 24123
rect 14642 24120 14648 24132
rect 14406 24092 14648 24120
rect 14406 24089 14418 24092
rect 14360 24083 14418 24089
rect 14642 24080 14648 24092
rect 14700 24080 14706 24132
rect 6178 24052 6184 24064
rect 5920 24024 6184 24052
rect 5813 24015 5871 24021
rect 6178 24012 6184 24024
rect 6236 24012 6242 24064
rect 7190 24012 7196 24064
rect 7248 24052 7254 24064
rect 7745 24055 7803 24061
rect 7745 24052 7757 24055
rect 7248 24024 7757 24052
rect 7248 24012 7254 24024
rect 7745 24021 7757 24024
rect 7791 24021 7803 24055
rect 7745 24015 7803 24021
rect 9398 24012 9404 24064
rect 9456 24052 9462 24064
rect 10042 24052 10048 24064
rect 9456 24024 10048 24052
rect 9456 24012 9462 24024
rect 10042 24012 10048 24024
rect 10100 24052 10106 24064
rect 10229 24055 10287 24061
rect 10229 24052 10241 24055
rect 10100 24024 10241 24052
rect 10100 24012 10106 24024
rect 10229 24021 10241 24024
rect 10275 24021 10287 24055
rect 10229 24015 10287 24021
rect 10965 24055 11023 24061
rect 10965 24021 10977 24055
rect 11011 24052 11023 24055
rect 12066 24052 12072 24064
rect 11011 24024 12072 24052
rect 11011 24021 11023 24024
rect 10965 24015 11023 24021
rect 12066 24012 12072 24024
rect 12124 24012 12130 24064
rect 12894 24012 12900 24064
rect 12952 24012 12958 24064
rect 13354 24012 13360 24064
rect 13412 24012 13418 24064
rect 13449 24055 13507 24061
rect 13449 24021 13461 24055
rect 13495 24052 13507 24055
rect 15102 24052 15108 24064
rect 13495 24024 15108 24052
rect 13495 24021 13507 24024
rect 13449 24015 13507 24021
rect 15102 24012 15108 24024
rect 15160 24052 15166 24064
rect 15488 24061 15516 24160
rect 16117 24157 16129 24160
rect 16163 24157 16175 24191
rect 16117 24151 16175 24157
rect 16485 24191 16543 24197
rect 16485 24157 16497 24191
rect 16531 24188 16543 24191
rect 16945 24191 17003 24197
rect 16945 24188 16957 24191
rect 16531 24160 16957 24188
rect 16531 24157 16543 24160
rect 16485 24151 16543 24157
rect 16945 24157 16957 24160
rect 16991 24157 17003 24191
rect 16945 24151 17003 24157
rect 18785 24191 18843 24197
rect 18785 24157 18797 24191
rect 18831 24188 18843 24191
rect 18831 24160 20116 24188
rect 18831 24157 18843 24160
rect 18785 24151 18843 24157
rect 20088 24132 20116 24160
rect 19794 24080 19800 24132
rect 19852 24120 19858 24132
rect 19950 24123 20008 24129
rect 19950 24120 19962 24123
rect 19852 24092 19962 24120
rect 19852 24080 19858 24092
rect 19950 24089 19962 24092
rect 19996 24089 20008 24123
rect 19950 24083 20008 24089
rect 20070 24080 20076 24132
rect 20128 24080 20134 24132
rect 15473 24055 15531 24061
rect 15473 24052 15485 24055
rect 15160 24024 15485 24052
rect 15160 24012 15166 24024
rect 15473 24021 15485 24024
rect 15519 24021 15531 24055
rect 15473 24015 15531 24021
rect 15562 24012 15568 24064
rect 15620 24012 15626 24064
rect 21174 24012 21180 24064
rect 21232 24012 21238 24064
rect 1104 23962 27876 23984
rect 1104 23910 4874 23962
rect 4926 23910 4938 23962
rect 4990 23910 5002 23962
rect 5054 23910 5066 23962
rect 5118 23910 5130 23962
rect 5182 23910 27876 23962
rect 1104 23888 27876 23910
rect 1210 23808 1216 23860
rect 1268 23848 1274 23860
rect 1489 23851 1547 23857
rect 1489 23848 1501 23851
rect 1268 23820 1501 23848
rect 1268 23808 1274 23820
rect 1489 23817 1501 23820
rect 1535 23817 1547 23851
rect 2774 23848 2780 23860
rect 1489 23811 1547 23817
rect 2516 23820 2780 23848
rect 2222 23780 2228 23792
rect 1688 23752 2228 23780
rect 1688 23721 1716 23752
rect 2222 23740 2228 23752
rect 2280 23740 2286 23792
rect 1673 23715 1731 23721
rect 1673 23681 1685 23715
rect 1719 23681 1731 23715
rect 1673 23675 1731 23681
rect 1946 23672 1952 23724
rect 2004 23672 2010 23724
rect 2516 23721 2544 23820
rect 2774 23808 2780 23820
rect 2832 23808 2838 23860
rect 3234 23808 3240 23860
rect 3292 23848 3298 23860
rect 3329 23851 3387 23857
rect 3329 23848 3341 23851
rect 3292 23820 3341 23848
rect 3292 23808 3298 23820
rect 3329 23817 3341 23820
rect 3375 23817 3387 23851
rect 3329 23811 3387 23817
rect 4801 23851 4859 23857
rect 4801 23817 4813 23851
rect 4847 23848 4859 23851
rect 5810 23848 5816 23860
rect 4847 23820 5816 23848
rect 4847 23817 4859 23820
rect 4801 23811 4859 23817
rect 5810 23808 5816 23820
rect 5868 23808 5874 23860
rect 7009 23851 7067 23857
rect 7009 23817 7021 23851
rect 7055 23817 7067 23851
rect 7009 23811 7067 23817
rect 2593 23783 2651 23789
rect 2593 23749 2605 23783
rect 2639 23780 2651 23783
rect 4442 23783 4500 23789
rect 4442 23780 4454 23783
rect 2639 23752 4454 23780
rect 2639 23749 2651 23752
rect 2593 23743 2651 23749
rect 4442 23749 4454 23752
rect 4488 23749 4500 23783
rect 4442 23743 4500 23749
rect 5936 23783 5994 23789
rect 5936 23749 5948 23783
rect 5982 23780 5994 23783
rect 7024 23780 7052 23811
rect 7190 23808 7196 23860
rect 7248 23808 7254 23860
rect 10410 23808 10416 23860
rect 10468 23848 10474 23860
rect 10468 23820 11284 23848
rect 10468 23808 10474 23820
rect 5982 23752 7052 23780
rect 9861 23783 9919 23789
rect 5982 23749 5994 23752
rect 5936 23743 5994 23749
rect 9861 23749 9873 23783
rect 9907 23780 9919 23783
rect 9950 23780 9956 23792
rect 9907 23752 9956 23780
rect 9907 23749 9919 23752
rect 9861 23743 9919 23749
rect 9950 23740 9956 23752
rect 10008 23740 10014 23792
rect 10229 23783 10287 23789
rect 10229 23749 10241 23783
rect 10275 23780 10287 23783
rect 10275 23752 11192 23780
rect 10275 23749 10287 23752
rect 10229 23743 10287 23749
rect 2501 23715 2559 23721
rect 2501 23681 2513 23715
rect 2547 23681 2559 23715
rect 2501 23675 2559 23681
rect 2685 23715 2743 23721
rect 2685 23681 2697 23715
rect 2731 23712 2743 23715
rect 2866 23712 2872 23724
rect 2731 23684 2872 23712
rect 2731 23681 2743 23684
rect 2685 23675 2743 23681
rect 2866 23672 2872 23684
rect 2924 23672 2930 23724
rect 2958 23672 2964 23724
rect 3016 23712 3022 23724
rect 3970 23712 3976 23724
rect 3016 23684 3976 23712
rect 3016 23672 3022 23684
rect 3970 23672 3976 23684
rect 4028 23672 4034 23724
rect 6914 23672 6920 23724
rect 6972 23712 6978 23724
rect 8205 23715 8263 23721
rect 8205 23712 8217 23715
rect 6972 23684 8217 23712
rect 6972 23672 6978 23684
rect 8205 23681 8217 23684
rect 8251 23681 8263 23715
rect 8205 23675 8263 23681
rect 10045 23715 10103 23721
rect 10045 23681 10057 23715
rect 10091 23712 10103 23715
rect 10318 23712 10324 23724
rect 10091 23684 10324 23712
rect 10091 23681 10103 23684
rect 10045 23675 10103 23681
rect 10318 23672 10324 23684
rect 10376 23672 10382 23724
rect 10505 23715 10563 23721
rect 10505 23681 10517 23715
rect 10551 23681 10563 23715
rect 10505 23675 10563 23681
rect 3145 23647 3203 23653
rect 3145 23613 3157 23647
rect 3191 23644 3203 23647
rect 3418 23644 3424 23656
rect 3191 23616 3424 23644
rect 3191 23613 3203 23616
rect 3145 23607 3203 23613
rect 3418 23604 3424 23616
rect 3476 23604 3482 23656
rect 4709 23647 4767 23653
rect 4709 23613 4721 23647
rect 4755 23644 4767 23647
rect 4798 23644 4804 23656
rect 4755 23616 4804 23644
rect 4755 23613 4767 23616
rect 4709 23607 4767 23613
rect 4798 23604 4804 23616
rect 4856 23604 4862 23656
rect 6181 23647 6239 23653
rect 6181 23613 6193 23647
rect 6227 23644 6239 23647
rect 7374 23644 7380 23656
rect 6227 23616 7380 23644
rect 6227 23613 6239 23616
rect 6181 23607 6239 23613
rect 7374 23604 7380 23616
rect 7432 23604 7438 23656
rect 10410 23604 10416 23656
rect 10468 23604 10474 23656
rect 7098 23536 7104 23588
rect 7156 23576 7162 23588
rect 7561 23579 7619 23585
rect 7561 23576 7573 23579
rect 7156 23548 7573 23576
rect 7156 23536 7162 23548
rect 7561 23545 7573 23548
rect 7607 23545 7619 23579
rect 7561 23539 7619 23545
rect 8386 23536 8392 23588
rect 8444 23536 8450 23588
rect 10520 23576 10548 23675
rect 10962 23672 10968 23724
rect 11020 23672 11026 23724
rect 11164 23721 11192 23752
rect 11256 23721 11284 23820
rect 14642 23808 14648 23860
rect 14700 23808 14706 23860
rect 15286 23808 15292 23860
rect 15344 23808 15350 23860
rect 15470 23857 15476 23860
rect 15457 23851 15476 23857
rect 15457 23817 15469 23851
rect 15457 23811 15476 23817
rect 15470 23808 15476 23811
rect 15528 23808 15534 23860
rect 16117 23851 16175 23857
rect 16117 23817 16129 23851
rect 16163 23848 16175 23851
rect 16482 23848 16488 23860
rect 16163 23820 16488 23848
rect 16163 23817 16175 23820
rect 16117 23811 16175 23817
rect 16482 23808 16488 23820
rect 16540 23808 16546 23860
rect 12704 23783 12762 23789
rect 12704 23749 12716 23783
rect 12750 23780 12762 23783
rect 12894 23780 12900 23792
rect 12750 23752 12900 23780
rect 12750 23749 12762 23752
rect 12704 23743 12762 23749
rect 12894 23740 12900 23752
rect 12952 23740 12958 23792
rect 13354 23740 13360 23792
rect 13412 23780 13418 23792
rect 15657 23783 15715 23789
rect 13412 23752 14872 23780
rect 13412 23740 13418 23752
rect 11149 23715 11207 23721
rect 11149 23681 11161 23715
rect 11195 23681 11207 23715
rect 11149 23675 11207 23681
rect 11241 23715 11299 23721
rect 11241 23681 11253 23715
rect 11287 23681 11299 23715
rect 11241 23675 11299 23681
rect 12066 23672 12072 23724
rect 12124 23672 12130 23724
rect 13078 23672 13084 23724
rect 13136 23712 13142 23724
rect 14844 23721 14872 23752
rect 15657 23749 15669 23783
rect 15703 23749 15715 23783
rect 20070 23780 20076 23792
rect 15657 23743 15715 23749
rect 19444 23752 20076 23780
rect 14829 23715 14887 23721
rect 13136 23684 14596 23712
rect 13136 23672 13142 23684
rect 12434 23604 12440 23656
rect 12492 23604 12498 23656
rect 14461 23647 14519 23653
rect 14461 23644 14473 23647
rect 13832 23616 14473 23644
rect 13832 23588 13860 23616
rect 14461 23613 14473 23616
rect 14507 23613 14519 23647
rect 14568 23644 14596 23684
rect 14829 23681 14841 23715
rect 14875 23681 14887 23715
rect 14829 23675 14887 23681
rect 14918 23672 14924 23724
rect 14976 23712 14982 23724
rect 15013 23715 15071 23721
rect 15013 23712 15025 23715
rect 14976 23684 15025 23712
rect 14976 23672 14982 23684
rect 15013 23681 15025 23684
rect 15059 23681 15071 23715
rect 15013 23675 15071 23681
rect 15105 23715 15163 23721
rect 15105 23681 15117 23715
rect 15151 23712 15163 23715
rect 15562 23712 15568 23724
rect 15151 23684 15568 23712
rect 15151 23681 15163 23684
rect 15105 23675 15163 23681
rect 15562 23672 15568 23684
rect 15620 23672 15626 23724
rect 15672 23644 15700 23743
rect 15930 23672 15936 23724
rect 15988 23672 15994 23724
rect 16209 23715 16267 23721
rect 16209 23681 16221 23715
rect 16255 23712 16267 23715
rect 16666 23712 16672 23724
rect 16255 23684 16672 23712
rect 16255 23681 16267 23684
rect 16209 23675 16267 23681
rect 16666 23672 16672 23684
rect 16724 23672 16730 23724
rect 19444 23721 19472 23752
rect 20070 23740 20076 23752
rect 20128 23740 20134 23792
rect 19429 23715 19487 23721
rect 19429 23681 19441 23715
rect 19475 23681 19487 23715
rect 21174 23712 21180 23724
rect 19429 23675 19487 23681
rect 19536 23684 21180 23712
rect 19536 23653 19564 23684
rect 21174 23672 21180 23684
rect 21232 23672 21238 23724
rect 14568 23616 15700 23644
rect 19521 23647 19579 23653
rect 14461 23607 14519 23613
rect 19521 23613 19533 23647
rect 19567 23613 19579 23647
rect 19521 23607 19579 23613
rect 19794 23604 19800 23656
rect 19852 23604 19858 23656
rect 11517 23579 11575 23585
rect 11517 23576 11529 23579
rect 10520 23548 11529 23576
rect 11517 23545 11529 23548
rect 11563 23545 11575 23579
rect 11517 23539 11575 23545
rect 13814 23536 13820 23588
rect 13872 23536 13878 23588
rect 1670 23468 1676 23520
rect 1728 23508 1734 23520
rect 1765 23511 1823 23517
rect 1765 23508 1777 23511
rect 1728 23480 1777 23508
rect 1728 23468 1734 23480
rect 1765 23477 1777 23480
rect 1811 23477 1823 23511
rect 1765 23471 1823 23477
rect 6178 23468 6184 23520
rect 6236 23508 6242 23520
rect 7193 23511 7251 23517
rect 7193 23508 7205 23511
rect 6236 23480 7205 23508
rect 6236 23468 6242 23480
rect 7193 23477 7205 23480
rect 7239 23508 7251 23511
rect 7742 23508 7748 23520
rect 7239 23480 7748 23508
rect 7239 23477 7251 23480
rect 7193 23471 7251 23477
rect 7742 23468 7748 23480
rect 7800 23468 7806 23520
rect 10778 23468 10784 23520
rect 10836 23468 10842 23520
rect 13909 23511 13967 23517
rect 13909 23477 13921 23511
rect 13955 23508 13967 23511
rect 13998 23508 14004 23520
rect 13955 23480 14004 23508
rect 13955 23477 13967 23480
rect 13909 23471 13967 23477
rect 13998 23468 14004 23480
rect 14056 23468 14062 23520
rect 15473 23511 15531 23517
rect 15473 23477 15485 23511
rect 15519 23508 15531 23511
rect 15749 23511 15807 23517
rect 15749 23508 15761 23511
rect 15519 23480 15761 23508
rect 15519 23477 15531 23480
rect 15473 23471 15531 23477
rect 15749 23477 15761 23480
rect 15795 23477 15807 23511
rect 15749 23471 15807 23477
rect 1104 23418 27876 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 27876 23418
rect 1104 23344 27876 23366
rect 2866 23264 2872 23316
rect 2924 23304 2930 23316
rect 3881 23307 3939 23313
rect 3881 23304 3893 23307
rect 2924 23276 3893 23304
rect 2924 23264 2930 23276
rect 3881 23273 3893 23276
rect 3927 23273 3939 23307
rect 3881 23267 3939 23273
rect 3970 23264 3976 23316
rect 4028 23264 4034 23316
rect 12802 23264 12808 23316
rect 12860 23264 12866 23316
rect 12897 23307 12955 23313
rect 12897 23273 12909 23307
rect 12943 23304 12955 23307
rect 12986 23304 12992 23316
rect 12943 23276 12992 23304
rect 12943 23273 12955 23276
rect 12897 23267 12955 23273
rect 12986 23264 12992 23276
rect 13044 23264 13050 23316
rect 13081 23307 13139 23313
rect 13081 23273 13093 23307
rect 13127 23273 13139 23307
rect 13081 23267 13139 23273
rect 13096 23236 13124 23267
rect 20898 23264 20904 23316
rect 20956 23304 20962 23316
rect 21545 23307 21603 23313
rect 21545 23304 21557 23307
rect 20956 23276 21557 23304
rect 20956 23264 20962 23276
rect 21545 23273 21557 23276
rect 21591 23273 21603 23307
rect 21545 23267 21603 23273
rect 10152 23208 13124 23236
rect 10152 23180 10180 23208
rect 20254 23196 20260 23248
rect 20312 23236 20318 23248
rect 20625 23239 20683 23245
rect 20625 23236 20637 23239
rect 20312 23208 20637 23236
rect 20312 23196 20318 23208
rect 20625 23205 20637 23208
rect 20671 23236 20683 23239
rect 20671 23208 21404 23236
rect 20671 23205 20683 23208
rect 20625 23199 20683 23205
rect 3050 23128 3056 23180
rect 3108 23168 3114 23180
rect 3789 23171 3847 23177
rect 3789 23168 3801 23171
rect 3108 23140 3801 23168
rect 3108 23128 3114 23140
rect 3789 23137 3801 23140
rect 3835 23137 3847 23171
rect 3789 23131 3847 23137
rect 7837 23171 7895 23177
rect 7837 23137 7849 23171
rect 7883 23168 7895 23171
rect 9677 23171 9735 23177
rect 9677 23168 9689 23171
rect 7883 23140 9689 23168
rect 7883 23137 7895 23140
rect 7837 23131 7895 23137
rect 9677 23137 9689 23140
rect 9723 23168 9735 23171
rect 10134 23168 10140 23180
rect 9723 23140 10140 23168
rect 9723 23137 9735 23140
rect 9677 23131 9735 23137
rect 10134 23128 10140 23140
rect 10192 23128 10198 23180
rect 12636 23140 12940 23168
rect 12636 23112 12664 23140
rect 3234 23060 3240 23112
rect 3292 23060 3298 23112
rect 3418 23060 3424 23112
rect 3476 23100 3482 23112
rect 4065 23103 4123 23109
rect 4065 23100 4077 23103
rect 3476 23072 4077 23100
rect 3476 23060 3482 23072
rect 4065 23069 4077 23072
rect 4111 23069 4123 23103
rect 4065 23063 4123 23069
rect 4798 23060 4804 23112
rect 4856 23100 4862 23112
rect 5261 23103 5319 23109
rect 5261 23100 5273 23103
rect 4856 23072 5273 23100
rect 4856 23060 4862 23072
rect 5261 23069 5273 23072
rect 5307 23069 5319 23103
rect 5261 23063 5319 23069
rect 6822 23060 6828 23112
rect 6880 23100 6886 23112
rect 7469 23103 7527 23109
rect 7469 23100 7481 23103
rect 6880 23072 7481 23100
rect 6880 23060 6886 23072
rect 7469 23069 7481 23072
rect 7515 23069 7527 23103
rect 7469 23063 7527 23069
rect 7653 23103 7711 23109
rect 7653 23069 7665 23103
rect 7699 23069 7711 23103
rect 7653 23063 7711 23069
rect 7282 22992 7288 23044
rect 7340 23032 7346 23044
rect 7668 23032 7696 23063
rect 8386 23060 8392 23112
rect 8444 23100 8450 23112
rect 8662 23100 8668 23112
rect 8444 23072 8668 23100
rect 8444 23060 8450 23072
rect 8662 23060 8668 23072
rect 8720 23100 8726 23112
rect 9217 23103 9275 23109
rect 9217 23100 9229 23103
rect 8720 23072 9229 23100
rect 8720 23060 8726 23072
rect 9217 23069 9229 23072
rect 9263 23069 9275 23103
rect 9217 23063 9275 23069
rect 9306 23060 9312 23112
rect 9364 23100 9370 23112
rect 9585 23103 9643 23109
rect 9585 23100 9597 23103
rect 9364 23072 9597 23100
rect 9364 23060 9370 23072
rect 9585 23069 9597 23072
rect 9631 23069 9643 23103
rect 9585 23063 9643 23069
rect 9766 23060 9772 23112
rect 9824 23060 9830 23112
rect 9861 23103 9919 23109
rect 9861 23069 9873 23103
rect 9907 23100 9919 23103
rect 10778 23100 10784 23112
rect 9907 23072 10784 23100
rect 9907 23069 9919 23072
rect 9861 23063 9919 23069
rect 10778 23060 10784 23072
rect 10836 23060 10842 23112
rect 12529 23103 12587 23109
rect 12529 23069 12541 23103
rect 12575 23100 12587 23103
rect 12618 23100 12624 23112
rect 12575 23072 12624 23100
rect 12575 23069 12587 23072
rect 12529 23063 12587 23069
rect 12618 23060 12624 23072
rect 12676 23060 12682 23112
rect 12805 23103 12863 23109
rect 12805 23069 12817 23103
rect 12851 23069 12863 23103
rect 12805 23063 12863 23069
rect 7340 23004 7696 23032
rect 7340 22992 7346 23004
rect 2682 22924 2688 22976
rect 2740 22924 2746 22976
rect 9030 22924 9036 22976
rect 9088 22924 9094 22976
rect 9214 22924 9220 22976
rect 9272 22964 9278 22976
rect 9401 22967 9459 22973
rect 9401 22964 9413 22967
rect 9272 22936 9413 22964
rect 9272 22924 9278 22936
rect 9401 22933 9413 22936
rect 9447 22933 9459 22967
rect 9401 22927 9459 22933
rect 12621 22967 12679 22973
rect 12621 22933 12633 22967
rect 12667 22964 12679 22967
rect 12710 22964 12716 22976
rect 12667 22936 12716 22964
rect 12667 22933 12679 22936
rect 12621 22927 12679 22933
rect 12710 22924 12716 22936
rect 12768 22924 12774 22976
rect 12820 22964 12848 23063
rect 12912 23032 12940 23140
rect 13170 23128 13176 23180
rect 13228 23168 13234 23180
rect 13449 23171 13507 23177
rect 13449 23168 13461 23171
rect 13228 23140 13461 23168
rect 13228 23128 13234 23140
rect 13449 23137 13461 23140
rect 13495 23137 13507 23171
rect 13449 23131 13507 23137
rect 13906 23128 13912 23180
rect 13964 23128 13970 23180
rect 19242 23128 19248 23180
rect 19300 23128 19306 23180
rect 20806 23128 20812 23180
rect 20864 23128 20870 23180
rect 13541 23103 13599 23109
rect 13541 23069 13553 23103
rect 13587 23100 13599 23103
rect 14093 23103 14151 23109
rect 14093 23100 14105 23103
rect 13587 23072 14105 23100
rect 13587 23069 13599 23072
rect 13541 23063 13599 23069
rect 14093 23069 14105 23072
rect 14139 23069 14151 23103
rect 14093 23063 14151 23069
rect 14642 23060 14648 23112
rect 14700 23060 14706 23112
rect 15010 23060 15016 23112
rect 15068 23100 15074 23112
rect 15381 23103 15439 23109
rect 15381 23100 15393 23103
rect 15068 23072 15393 23100
rect 15068 23060 15074 23072
rect 15381 23069 15393 23072
rect 15427 23069 15439 23103
rect 15381 23063 15439 23069
rect 16666 23060 16672 23112
rect 16724 23100 16730 23112
rect 17129 23103 17187 23109
rect 17129 23100 17141 23103
rect 16724 23072 17141 23100
rect 16724 23060 16730 23072
rect 17129 23069 17141 23072
rect 17175 23100 17187 23103
rect 17405 23103 17463 23109
rect 17405 23100 17417 23103
rect 17175 23072 17417 23100
rect 17175 23069 17187 23072
rect 17129 23063 17187 23069
rect 17405 23069 17417 23072
rect 17451 23100 17463 23103
rect 19260 23100 19288 23128
rect 17451 23072 19288 23100
rect 17451 23069 17463 23072
rect 17405 23063 17463 23069
rect 20714 23060 20720 23112
rect 20772 23100 20778 23112
rect 21376 23109 21404 23208
rect 20901 23103 20959 23109
rect 20901 23100 20913 23103
rect 20772 23072 20913 23100
rect 20772 23060 20778 23072
rect 20901 23069 20913 23072
rect 20947 23069 20959 23103
rect 20901 23063 20959 23069
rect 21361 23103 21419 23109
rect 21361 23069 21373 23103
rect 21407 23069 21419 23103
rect 21361 23063 21419 23069
rect 13049 23035 13107 23041
rect 13049 23032 13061 23035
rect 12912 23004 13061 23032
rect 13049 23001 13061 23004
rect 13095 23001 13107 23035
rect 13049 22995 13107 23001
rect 13265 23035 13323 23041
rect 13265 23001 13277 23035
rect 13311 23032 13323 23035
rect 13814 23032 13820 23044
rect 13311 23004 13820 23032
rect 13311 23001 13323 23004
rect 13265 22995 13323 23001
rect 13814 22992 13820 23004
rect 13872 22992 13878 23044
rect 17310 22992 17316 23044
rect 17368 23032 17374 23044
rect 17650 23035 17708 23041
rect 17650 23032 17662 23035
rect 17368 23004 17662 23032
rect 17368 22992 17374 23004
rect 17650 23001 17662 23004
rect 17696 23001 17708 23035
rect 17650 22995 17708 23001
rect 18966 22992 18972 23044
rect 19024 23032 19030 23044
rect 19490 23035 19548 23041
rect 19490 23032 19502 23035
rect 19024 23004 19502 23032
rect 19024 22992 19030 23004
rect 19490 23001 19502 23004
rect 19536 23001 19548 23035
rect 19490 22995 19548 23001
rect 13998 22964 14004 22976
rect 12820 22936 14004 22964
rect 13998 22924 14004 22936
rect 14056 22924 14062 22976
rect 18782 22924 18788 22976
rect 18840 22924 18846 22976
rect 21266 22924 21272 22976
rect 21324 22924 21330 22976
rect 1104 22874 27876 22896
rect 1104 22822 4874 22874
rect 4926 22822 4938 22874
rect 4990 22822 5002 22874
rect 5054 22822 5066 22874
rect 5118 22822 5130 22874
rect 5182 22822 27876 22874
rect 1104 22800 27876 22822
rect 6825 22763 6883 22769
rect 6825 22729 6837 22763
rect 6871 22760 6883 22763
rect 6914 22760 6920 22772
rect 6871 22732 6920 22760
rect 6871 22729 6883 22732
rect 6825 22723 6883 22729
rect 6914 22720 6920 22732
rect 6972 22720 6978 22772
rect 8570 22720 8576 22772
rect 8628 22760 8634 22772
rect 8757 22763 8815 22769
rect 8757 22760 8769 22763
rect 8628 22732 8769 22760
rect 8628 22720 8634 22732
rect 8757 22729 8769 22732
rect 8803 22729 8815 22763
rect 8757 22723 8815 22729
rect 9309 22763 9367 22769
rect 9309 22729 9321 22763
rect 9355 22760 9367 22763
rect 9355 22732 9536 22760
rect 9355 22729 9367 22732
rect 9309 22723 9367 22729
rect 2492 22695 2550 22701
rect 2492 22661 2504 22695
rect 2538 22692 2550 22695
rect 2682 22692 2688 22704
rect 2538 22664 2688 22692
rect 2538 22661 2550 22664
rect 2492 22655 2550 22661
rect 2682 22652 2688 22664
rect 2740 22652 2746 22704
rect 9508 22692 9536 22732
rect 10778 22720 10784 22772
rect 10836 22760 10842 22772
rect 11701 22763 11759 22769
rect 11701 22760 11713 22763
rect 10836 22732 11713 22760
rect 10836 22720 10842 22732
rect 11701 22729 11713 22732
rect 11747 22729 11759 22763
rect 11701 22723 11759 22729
rect 11793 22763 11851 22769
rect 11793 22729 11805 22763
rect 11839 22760 11851 22763
rect 12066 22760 12072 22772
rect 11839 22732 12072 22760
rect 11839 22729 11851 22732
rect 11793 22723 11851 22729
rect 9646 22695 9704 22701
rect 9646 22692 9658 22695
rect 9508 22664 9658 22692
rect 9646 22661 9658 22664
rect 9692 22661 9704 22695
rect 9646 22655 9704 22661
rect 10318 22652 10324 22704
rect 10376 22692 10382 22704
rect 10873 22695 10931 22701
rect 10873 22692 10885 22695
rect 10376 22664 10885 22692
rect 10376 22652 10382 22664
rect 10873 22661 10885 22664
rect 10919 22692 10931 22695
rect 10962 22692 10968 22704
rect 10919 22664 10968 22692
rect 10919 22661 10931 22664
rect 10873 22655 10931 22661
rect 10962 22652 10968 22664
rect 11020 22652 11026 22704
rect 11808 22692 11836 22723
rect 12066 22720 12072 22732
rect 12124 22720 12130 22772
rect 14369 22763 14427 22769
rect 14369 22729 14381 22763
rect 14415 22760 14427 22763
rect 14642 22760 14648 22772
rect 14415 22732 14648 22760
rect 14415 22729 14427 22732
rect 14369 22723 14427 22729
rect 14642 22720 14648 22732
rect 14700 22720 14706 22772
rect 16206 22760 16212 22772
rect 16040 22732 16212 22760
rect 11072 22664 11836 22692
rect 11992 22664 12572 22692
rect 1394 22584 1400 22636
rect 1452 22624 1458 22636
rect 2225 22627 2283 22633
rect 2225 22624 2237 22627
rect 1452 22596 2237 22624
rect 1452 22584 1458 22596
rect 2225 22593 2237 22596
rect 2271 22624 2283 22627
rect 2314 22624 2320 22636
rect 2271 22596 2320 22624
rect 2271 22593 2283 22596
rect 2225 22587 2283 22593
rect 2314 22584 2320 22596
rect 2372 22584 2378 22636
rect 5068 22627 5126 22633
rect 5068 22593 5080 22627
rect 5114 22624 5126 22627
rect 5442 22624 5448 22636
rect 5114 22596 5448 22624
rect 5114 22593 5126 22596
rect 5068 22587 5126 22593
rect 5442 22584 5448 22596
rect 5500 22584 5506 22636
rect 6641 22627 6699 22633
rect 6641 22593 6653 22627
rect 6687 22624 6699 22627
rect 6822 22624 6828 22636
rect 6687 22596 6828 22624
rect 6687 22593 6699 22596
rect 6641 22587 6699 22593
rect 6822 22584 6828 22596
rect 6880 22584 6886 22636
rect 7650 22633 7656 22636
rect 7644 22587 7656 22633
rect 7650 22584 7656 22587
rect 7708 22584 7714 22636
rect 9398 22584 9404 22636
rect 9456 22584 9462 22636
rect 9950 22624 9956 22636
rect 9508 22596 9956 22624
rect 4433 22559 4491 22565
rect 4433 22525 4445 22559
rect 4479 22525 4491 22559
rect 4433 22519 4491 22525
rect 3605 22491 3663 22497
rect 3605 22457 3617 22491
rect 3651 22488 3663 22491
rect 4448 22488 4476 22519
rect 4798 22516 4804 22568
rect 4856 22516 4862 22568
rect 6457 22559 6515 22565
rect 6457 22556 6469 22559
rect 6196 22528 6469 22556
rect 4706 22488 4712 22500
rect 3651 22460 4712 22488
rect 3651 22457 3663 22460
rect 3605 22451 3663 22457
rect 4706 22448 4712 22460
rect 4764 22448 4770 22500
rect 6196 22497 6224 22528
rect 6457 22525 6469 22528
rect 6503 22556 6515 22559
rect 6730 22556 6736 22568
rect 6503 22528 6736 22556
rect 6503 22525 6515 22528
rect 6457 22519 6515 22525
rect 6730 22516 6736 22528
rect 6788 22556 6794 22568
rect 7282 22556 7288 22568
rect 6788 22528 7288 22556
rect 6788 22516 6794 22528
rect 7282 22516 7288 22528
rect 7340 22516 7346 22568
rect 7374 22516 7380 22568
rect 7432 22516 7438 22568
rect 8849 22559 8907 22565
rect 8849 22525 8861 22559
rect 8895 22556 8907 22559
rect 9508 22556 9536 22596
rect 9950 22584 9956 22596
rect 10008 22584 10014 22636
rect 11072 22633 11100 22664
rect 11057 22627 11115 22633
rect 11057 22593 11069 22627
rect 11103 22593 11115 22627
rect 11057 22587 11115 22593
rect 11149 22627 11207 22633
rect 11149 22593 11161 22627
rect 11195 22593 11207 22627
rect 11149 22587 11207 22593
rect 8895 22528 9536 22556
rect 8895 22525 8907 22528
rect 8849 22519 8907 22525
rect 10962 22516 10968 22568
rect 11020 22556 11026 22568
rect 11164 22556 11192 22587
rect 11238 22584 11244 22636
rect 11296 22624 11302 22636
rect 11885 22627 11943 22633
rect 11885 22624 11897 22627
rect 11296 22596 11897 22624
rect 11296 22584 11302 22596
rect 11885 22593 11897 22596
rect 11931 22593 11943 22627
rect 11885 22587 11943 22593
rect 11517 22559 11575 22565
rect 11517 22556 11529 22559
rect 11020 22528 11529 22556
rect 11020 22516 11026 22528
rect 11517 22525 11529 22528
rect 11563 22525 11575 22559
rect 11992 22556 12020 22664
rect 12544 22633 12572 22664
rect 13906 22652 13912 22704
rect 13964 22692 13970 22704
rect 16040 22701 16068 22732
rect 16206 22720 16212 22732
rect 16264 22720 16270 22772
rect 16393 22763 16451 22769
rect 16393 22729 16405 22763
rect 16439 22760 16451 22763
rect 16439 22732 16574 22760
rect 16439 22729 16451 22732
rect 16393 22723 16451 22729
rect 15482 22695 15540 22701
rect 15482 22692 15494 22695
rect 13964 22664 15494 22692
rect 13964 22652 13970 22664
rect 15482 22661 15494 22664
rect 15528 22661 15540 22695
rect 15482 22655 15540 22661
rect 16025 22695 16083 22701
rect 16025 22661 16037 22695
rect 16071 22661 16083 22695
rect 16546 22692 16574 22732
rect 18966 22720 18972 22772
rect 19024 22720 19030 22772
rect 21266 22720 21272 22772
rect 21324 22720 21330 22772
rect 16914 22695 16972 22701
rect 16914 22692 16926 22695
rect 16546 22664 16926 22692
rect 16025 22655 16083 22661
rect 16914 22661 16926 22664
rect 16960 22661 16972 22695
rect 16914 22655 16972 22661
rect 17034 22652 17040 22704
rect 17092 22692 17098 22704
rect 18233 22695 18291 22701
rect 18233 22692 18245 22695
rect 17092 22664 18245 22692
rect 17092 22652 17098 22664
rect 18233 22661 18245 22664
rect 18279 22661 18291 22695
rect 18233 22655 18291 22661
rect 19245 22695 19303 22701
rect 19245 22661 19257 22695
rect 19291 22692 19303 22695
rect 19613 22695 19671 22701
rect 19613 22692 19625 22695
rect 19291 22664 19625 22692
rect 19291 22661 19303 22664
rect 19245 22655 19303 22661
rect 19613 22661 19625 22664
rect 19659 22661 19671 22695
rect 19613 22655 19671 22661
rect 12437 22627 12495 22633
rect 12437 22593 12449 22627
rect 12483 22593 12495 22627
rect 12437 22587 12495 22593
rect 12529 22627 12587 22633
rect 12529 22593 12541 22627
rect 12575 22593 12587 22627
rect 12529 22587 12587 22593
rect 11517 22519 11575 22525
rect 11624 22528 12020 22556
rect 6181 22491 6239 22497
rect 6181 22457 6193 22491
rect 6227 22457 6239 22491
rect 6181 22451 6239 22457
rect 9214 22448 9220 22500
rect 9272 22448 9278 22500
rect 10410 22448 10416 22500
rect 10468 22488 10474 22500
rect 11624 22488 11652 22528
rect 12452 22488 12480 22587
rect 15838 22584 15844 22636
rect 15896 22584 15902 22636
rect 16114 22584 16120 22636
rect 16172 22584 16178 22636
rect 16209 22627 16267 22633
rect 16209 22593 16221 22627
rect 16255 22624 16267 22627
rect 16298 22624 16304 22636
rect 16255 22596 16304 22624
rect 16255 22593 16267 22596
rect 16209 22587 16267 22593
rect 16298 22584 16304 22596
rect 16356 22584 16362 22636
rect 16666 22624 16672 22636
rect 16546 22596 16672 22624
rect 13630 22516 13636 22568
rect 13688 22516 13694 22568
rect 15749 22559 15807 22565
rect 15749 22525 15761 22559
rect 15795 22556 15807 22559
rect 16546 22556 16574 22596
rect 16666 22584 16672 22596
rect 16724 22584 16730 22636
rect 18690 22584 18696 22636
rect 18748 22624 18754 22636
rect 19153 22627 19211 22633
rect 19153 22624 19165 22627
rect 18748 22596 19165 22624
rect 18748 22584 18754 22596
rect 19153 22593 19165 22596
rect 19199 22593 19211 22627
rect 19153 22587 19211 22593
rect 19334 22584 19340 22636
rect 19392 22584 19398 22636
rect 19521 22627 19579 22633
rect 19521 22593 19533 22627
rect 19567 22624 19579 22627
rect 21177 22627 21235 22633
rect 19567 22596 20852 22624
rect 19567 22593 19579 22596
rect 19521 22587 19579 22593
rect 15795 22528 16574 22556
rect 15795 22525 15807 22528
rect 15749 22519 15807 22525
rect 18138 22516 18144 22568
rect 18196 22556 18202 22568
rect 18782 22556 18788 22568
rect 18196 22528 18788 22556
rect 18196 22516 18202 22528
rect 18782 22516 18788 22528
rect 18840 22516 18846 22568
rect 20254 22516 20260 22568
rect 20312 22516 20318 22568
rect 12713 22491 12771 22497
rect 12713 22488 12725 22491
rect 10468 22460 11652 22488
rect 11900 22460 12388 22488
rect 12452 22460 12725 22488
rect 10468 22448 10474 22460
rect 3878 22380 3884 22432
rect 3936 22380 3942 22432
rect 8294 22380 8300 22432
rect 8352 22420 8358 22432
rect 9030 22420 9036 22432
rect 8352 22392 9036 22420
rect 8352 22380 8358 22392
rect 9030 22380 9036 22392
rect 9088 22380 9094 22432
rect 10778 22380 10784 22432
rect 10836 22420 10842 22432
rect 10873 22423 10931 22429
rect 10873 22420 10885 22423
rect 10836 22392 10885 22420
rect 10836 22380 10842 22392
rect 10873 22389 10885 22392
rect 10919 22389 10931 22423
rect 10873 22383 10931 22389
rect 11333 22423 11391 22429
rect 11333 22389 11345 22423
rect 11379 22420 11391 22423
rect 11900 22420 11928 22460
rect 11379 22392 11928 22420
rect 11379 22389 11391 22392
rect 11333 22383 11391 22389
rect 12066 22380 12072 22432
rect 12124 22380 12130 22432
rect 12158 22380 12164 22432
rect 12216 22420 12222 22432
rect 12253 22423 12311 22429
rect 12253 22420 12265 22423
rect 12216 22392 12265 22420
rect 12216 22380 12222 22392
rect 12253 22389 12265 22392
rect 12299 22389 12311 22423
rect 12360 22420 12388 22460
rect 12713 22457 12725 22460
rect 12759 22488 12771 22491
rect 14366 22488 14372 22500
rect 12759 22460 14372 22488
rect 12759 22457 12771 22460
rect 12713 22451 12771 22457
rect 14366 22448 14372 22460
rect 14424 22448 14430 22500
rect 20824 22497 20852 22596
rect 21177 22593 21189 22627
rect 21223 22624 21235 22627
rect 21223 22596 21864 22624
rect 21223 22593 21235 22596
rect 21177 22587 21235 22593
rect 21358 22516 21364 22568
rect 21416 22516 21422 22568
rect 21836 22565 21864 22596
rect 22186 22584 22192 22636
rect 22244 22584 22250 22636
rect 21821 22559 21879 22565
rect 21821 22525 21833 22559
rect 21867 22525 21879 22559
rect 21821 22519 21879 22525
rect 22094 22516 22100 22568
rect 22152 22516 22158 22568
rect 20809 22491 20867 22497
rect 20809 22457 20821 22491
rect 20855 22457 20867 22491
rect 20809 22451 20867 22457
rect 12894 22420 12900 22432
rect 12360 22392 12900 22420
rect 12253 22383 12311 22389
rect 12894 22380 12900 22392
rect 12952 22380 12958 22432
rect 13078 22380 13084 22432
rect 13136 22380 13142 22432
rect 16022 22380 16028 22432
rect 16080 22420 16086 22432
rect 18049 22423 18107 22429
rect 18049 22420 18061 22423
rect 16080 22392 18061 22420
rect 16080 22380 16086 22392
rect 18049 22389 18061 22392
rect 18095 22389 18107 22423
rect 18049 22383 18107 22389
rect 1104 22330 27876 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 27876 22330
rect 1104 22256 27876 22278
rect 2777 22219 2835 22225
rect 2777 22185 2789 22219
rect 2823 22216 2835 22219
rect 3234 22216 3240 22228
rect 2823 22188 3240 22216
rect 2823 22185 2835 22188
rect 2777 22179 2835 22185
rect 3234 22176 3240 22188
rect 3292 22176 3298 22228
rect 4798 22216 4804 22228
rect 3804 22188 4804 22216
rect 1394 22040 1400 22092
rect 1452 22040 1458 22092
rect 2406 22040 2412 22092
rect 2464 22080 2470 22092
rect 3804 22089 3832 22188
rect 4798 22176 4804 22188
rect 4856 22216 4862 22228
rect 5537 22219 5595 22225
rect 5537 22216 5549 22219
rect 4856 22188 5549 22216
rect 4856 22176 4862 22188
rect 5537 22185 5549 22188
rect 5583 22185 5595 22219
rect 5537 22179 5595 22185
rect 6914 22176 6920 22228
rect 6972 22216 6978 22228
rect 7561 22219 7619 22225
rect 7561 22216 7573 22219
rect 6972 22188 7573 22216
rect 6972 22176 6978 22188
rect 7561 22185 7573 22188
rect 7607 22185 7619 22219
rect 7561 22179 7619 22185
rect 7650 22176 7656 22228
rect 7708 22216 7714 22228
rect 7745 22219 7803 22225
rect 7745 22216 7757 22219
rect 7708 22188 7757 22216
rect 7708 22176 7714 22188
rect 7745 22185 7757 22188
rect 7791 22185 7803 22219
rect 7745 22179 7803 22185
rect 12437 22219 12495 22225
rect 12437 22185 12449 22219
rect 12483 22185 12495 22219
rect 12437 22179 12495 22185
rect 7024 22120 7328 22148
rect 7024 22092 7052 22120
rect 3789 22083 3847 22089
rect 3789 22080 3801 22083
rect 2464 22052 3801 22080
rect 2464 22040 2470 22052
rect 3789 22049 3801 22052
rect 3835 22049 3847 22083
rect 3789 22043 3847 22049
rect 7006 22040 7012 22092
rect 7064 22040 7070 22092
rect 1670 22021 1676 22024
rect 1664 21975 1676 22021
rect 1670 21972 1676 21975
rect 1728 21972 1734 22024
rect 3878 21972 3884 22024
rect 3936 22012 3942 22024
rect 4045 22015 4103 22021
rect 4045 22012 4057 22015
rect 3936 21984 4057 22012
rect 3936 21972 3942 21984
rect 4045 21981 4057 21984
rect 4091 21981 4103 22015
rect 4045 21975 4103 21981
rect 7101 22015 7159 22021
rect 7101 21981 7113 22015
rect 7147 22012 7159 22015
rect 7190 22012 7196 22024
rect 7147 21984 7196 22012
rect 7147 21981 7159 21984
rect 7101 21975 7159 21981
rect 7190 21972 7196 21984
rect 7248 21972 7254 22024
rect 7300 22012 7328 22120
rect 9766 22108 9772 22160
rect 9824 22148 9830 22160
rect 10413 22151 10471 22157
rect 10413 22148 10425 22151
rect 9824 22120 10425 22148
rect 9824 22108 9830 22120
rect 10413 22117 10425 22120
rect 10459 22148 10471 22151
rect 10962 22148 10968 22160
rect 10459 22120 10968 22148
rect 10459 22117 10471 22120
rect 10413 22111 10471 22117
rect 10962 22108 10968 22120
rect 11020 22108 11026 22160
rect 12066 22148 12072 22160
rect 11900 22120 12072 22148
rect 7377 22015 7435 22021
rect 7377 22012 7389 22015
rect 7300 21984 7389 22012
rect 7377 21981 7389 21984
rect 7423 22012 7435 22015
rect 8021 22015 8079 22021
rect 8021 22012 8033 22015
rect 7423 21984 8033 22012
rect 7423 21981 7435 21984
rect 7377 21975 7435 21981
rect 8021 21981 8033 21984
rect 8067 22012 8079 22015
rect 8202 22012 8208 22024
rect 8067 21984 8208 22012
rect 8067 21981 8079 21984
rect 8021 21975 8079 21981
rect 8202 21972 8208 21984
rect 8260 21972 8266 22024
rect 8386 21972 8392 22024
rect 8444 21972 8450 22024
rect 8478 21972 8484 22024
rect 8536 21972 8542 22024
rect 9861 22015 9919 22021
rect 9861 21981 9873 22015
rect 9907 22012 9919 22015
rect 9950 22012 9956 22024
rect 9907 21984 9956 22012
rect 9907 21981 9919 21984
rect 9861 21975 9919 21981
rect 9950 21972 9956 21984
rect 10008 21972 10014 22024
rect 10229 22015 10287 22021
rect 10229 21981 10241 22015
rect 10275 22012 10287 22015
rect 10778 22012 10784 22024
rect 10275 21984 10784 22012
rect 10275 21981 10287 21984
rect 10229 21975 10287 21981
rect 10778 21972 10784 21984
rect 10836 21972 10842 22024
rect 11900 22021 11928 22120
rect 12066 22108 12072 22120
rect 12124 22148 12130 22160
rect 12452 22148 12480 22179
rect 12526 22176 12532 22228
rect 12584 22216 12590 22228
rect 13630 22216 13636 22228
rect 12584 22188 13636 22216
rect 12584 22176 12590 22188
rect 13630 22176 13636 22188
rect 13688 22176 13694 22228
rect 13722 22176 13728 22228
rect 13780 22216 13786 22228
rect 16298 22216 16304 22228
rect 13780 22188 16304 22216
rect 13780 22176 13786 22188
rect 16298 22176 16304 22188
rect 16356 22176 16362 22228
rect 17310 22176 17316 22228
rect 17368 22176 17374 22228
rect 12124 22120 12664 22148
rect 12124 22108 12130 22120
rect 12526 22080 12532 22092
rect 12268 22052 12532 22080
rect 11425 22015 11483 22021
rect 11425 21981 11437 22015
rect 11471 21981 11483 22015
rect 11425 21975 11483 21981
rect 11609 22015 11667 22021
rect 11609 21981 11621 22015
rect 11655 22012 11667 22015
rect 11885 22015 11943 22021
rect 11655 21984 11836 22012
rect 11655 21981 11667 21984
rect 11609 21975 11667 21981
rect 7006 21904 7012 21956
rect 7064 21944 7070 21956
rect 7064 21916 7696 21944
rect 7064 21904 7070 21916
rect 5169 21879 5227 21885
rect 5169 21845 5181 21879
rect 5215 21876 5227 21879
rect 5258 21876 5264 21888
rect 5215 21848 5264 21876
rect 5215 21845 5227 21848
rect 5169 21839 5227 21845
rect 5258 21836 5264 21848
rect 5316 21836 5322 21888
rect 6730 21836 6736 21888
rect 6788 21876 6794 21888
rect 7193 21879 7251 21885
rect 7193 21876 7205 21879
rect 6788 21848 7205 21876
rect 6788 21836 6794 21848
rect 7193 21845 7205 21848
rect 7239 21845 7251 21879
rect 7668 21876 7696 21916
rect 7742 21904 7748 21956
rect 7800 21904 7806 21956
rect 7929 21947 7987 21953
rect 7929 21913 7941 21947
rect 7975 21944 7987 21947
rect 8404 21944 8432 21972
rect 7975 21916 8432 21944
rect 7975 21913 7987 21916
rect 7929 21907 7987 21913
rect 9766 21904 9772 21956
rect 9824 21944 9830 21956
rect 10045 21947 10103 21953
rect 10045 21944 10057 21947
rect 9824 21916 10057 21944
rect 9824 21904 9830 21916
rect 10045 21913 10057 21916
rect 10091 21944 10103 21947
rect 10410 21944 10416 21956
rect 10091 21916 10416 21944
rect 10091 21913 10103 21916
rect 10045 21907 10103 21913
rect 10410 21904 10416 21916
rect 10468 21904 10474 21956
rect 11440 21944 11468 21975
rect 11440 21916 11652 21944
rect 8938 21876 8944 21888
rect 7668 21848 8944 21876
rect 7193 21839 7251 21845
rect 8938 21836 8944 21848
rect 8996 21836 9002 21888
rect 10134 21836 10140 21888
rect 10192 21836 10198 21888
rect 11514 21836 11520 21888
rect 11572 21836 11578 21888
rect 11624 21876 11652 21916
rect 11698 21904 11704 21956
rect 11756 21904 11762 21956
rect 11808 21944 11836 21984
rect 11885 21981 11897 22015
rect 11931 21981 11943 22015
rect 11885 21975 11943 21981
rect 11977 22015 12035 22021
rect 11977 21981 11989 22015
rect 12023 22012 12035 22015
rect 12158 22012 12164 22024
rect 12023 21984 12164 22012
rect 12023 21981 12035 21984
rect 11977 21975 12035 21981
rect 12158 21972 12164 21984
rect 12216 21972 12222 22024
rect 11808 21916 12020 21944
rect 11799 21879 11857 21885
rect 11799 21876 11811 21879
rect 11624 21848 11811 21876
rect 11799 21845 11811 21848
rect 11845 21845 11857 21879
rect 11992 21876 12020 21916
rect 12066 21904 12072 21956
rect 12124 21944 12130 21956
rect 12268 21953 12296 22052
rect 12526 22040 12532 22052
rect 12584 22040 12590 22092
rect 12253 21947 12311 21953
rect 12253 21944 12265 21947
rect 12124 21916 12265 21944
rect 12124 21904 12130 21916
rect 12253 21913 12265 21916
rect 12299 21913 12311 21947
rect 12253 21907 12311 21913
rect 12342 21904 12348 21956
rect 12400 21944 12406 21956
rect 12453 21947 12511 21953
rect 12453 21944 12465 21947
rect 12400 21916 12465 21944
rect 12400 21904 12406 21916
rect 12453 21913 12465 21916
rect 12499 21913 12511 21947
rect 12636 21944 12664 22120
rect 12894 22108 12900 22160
rect 12952 22148 12958 22160
rect 13449 22151 13507 22157
rect 13449 22148 13461 22151
rect 12952 22120 13461 22148
rect 12952 22108 12958 22120
rect 13449 22117 13461 22120
rect 13495 22117 13507 22151
rect 13449 22111 13507 22117
rect 13541 22151 13599 22157
rect 13541 22117 13553 22151
rect 13587 22148 13599 22151
rect 13587 22120 14412 22148
rect 13587 22117 13599 22120
rect 13541 22111 13599 22117
rect 12986 22040 12992 22092
rect 13044 22080 13050 22092
rect 13722 22080 13728 22092
rect 13044 22052 13728 22080
rect 13044 22040 13050 22052
rect 13722 22040 13728 22052
rect 13780 22040 13786 22092
rect 13354 21972 13360 22024
rect 13412 21972 13418 22024
rect 13814 21972 13820 22024
rect 13872 22012 13878 22024
rect 14384 22021 14412 22120
rect 16942 22108 16948 22160
rect 17000 22148 17006 22160
rect 17000 22120 18552 22148
rect 17000 22108 17006 22120
rect 15470 22040 15476 22092
rect 15528 22080 15534 22092
rect 18138 22080 18144 22092
rect 15528 22052 18144 22080
rect 15528 22040 15534 22052
rect 18138 22040 18144 22052
rect 18196 22080 18202 22092
rect 18524 22080 18552 22120
rect 18196 22052 18276 22080
rect 18196 22040 18202 22052
rect 14093 22015 14151 22021
rect 14093 22012 14105 22015
rect 13872 21984 14105 22012
rect 13872 21972 13878 21984
rect 14093 21981 14105 21984
rect 14139 21981 14151 22015
rect 14369 22015 14427 22021
rect 14369 22012 14381 22015
rect 14327 21984 14381 22012
rect 14093 21975 14151 21981
rect 14369 21981 14381 21984
rect 14415 22012 14427 22015
rect 14642 22012 14648 22024
rect 14415 21984 14648 22012
rect 14415 21981 14427 21984
rect 14369 21975 14427 21981
rect 14642 21972 14648 21984
rect 14700 21972 14706 22024
rect 15562 21972 15568 22024
rect 15620 21972 15626 22024
rect 15749 22015 15807 22021
rect 15749 21981 15761 22015
rect 15795 22012 15807 22015
rect 16114 22012 16120 22024
rect 15795 21984 16120 22012
rect 15795 21981 15807 21984
rect 15749 21975 15807 21981
rect 16114 21972 16120 21984
rect 16172 21972 16178 22024
rect 16666 21972 16672 22024
rect 16724 22012 16730 22024
rect 16761 22015 16819 22021
rect 16761 22012 16773 22015
rect 16724 21984 16773 22012
rect 16724 21972 16730 21984
rect 16761 21981 16773 21984
rect 16807 21981 16819 22015
rect 16761 21975 16819 21981
rect 17034 21972 17040 22024
rect 17092 21972 17098 22024
rect 17175 22015 17233 22021
rect 17175 21981 17187 22015
rect 17221 21981 17233 22015
rect 17175 21975 17233 21981
rect 12636 21916 12756 21944
rect 12453 21907 12511 21913
rect 12618 21876 12624 21888
rect 11992 21848 12624 21876
rect 11799 21839 11857 21845
rect 12618 21836 12624 21848
rect 12676 21836 12682 21888
rect 12728 21876 12756 21916
rect 12802 21904 12808 21956
rect 12860 21904 12866 21956
rect 14461 21947 14519 21953
rect 14461 21944 14473 21947
rect 13004 21916 14473 21944
rect 13004 21876 13032 21916
rect 14461 21913 14473 21916
rect 14507 21913 14519 21947
rect 14461 21907 14519 21913
rect 16206 21904 16212 21956
rect 16264 21944 16270 21956
rect 16942 21944 16948 21956
rect 16264 21916 16948 21944
rect 16264 21904 16270 21916
rect 16942 21904 16948 21916
rect 17000 21904 17006 21956
rect 17190 21944 17218 21975
rect 17586 21972 17592 22024
rect 17644 21972 17650 22024
rect 17862 21972 17868 22024
rect 17920 21972 17926 22024
rect 18248 22021 18276 22052
rect 18524 22052 19196 22080
rect 18233 22015 18291 22021
rect 18233 21981 18245 22015
rect 18279 21981 18291 22015
rect 18233 21975 18291 21981
rect 18325 22015 18383 22021
rect 18325 21981 18337 22015
rect 18371 22012 18383 22015
rect 18414 22012 18420 22024
rect 18371 21984 18420 22012
rect 18371 21981 18383 21984
rect 18325 21975 18383 21981
rect 18414 21972 18420 21984
rect 18472 21972 18478 22024
rect 18524 22021 18552 22052
rect 18509 22015 18567 22021
rect 18509 21981 18521 22015
rect 18555 21981 18567 22015
rect 18509 21975 18567 21981
rect 18690 21972 18696 22024
rect 18748 21972 18754 22024
rect 19168 22012 19196 22052
rect 19242 22040 19248 22092
rect 19300 22040 19306 22092
rect 20990 22080 20996 22092
rect 20824 22052 20996 22080
rect 19334 22012 19340 22024
rect 19168 21984 19340 22012
rect 19334 21972 19340 21984
rect 19392 21972 19398 22024
rect 20824 22021 20852 22052
rect 20990 22040 20996 22052
rect 21048 22080 21054 22092
rect 22278 22080 22284 22092
rect 21048 22052 22284 22080
rect 21048 22040 21054 22052
rect 22278 22040 22284 22052
rect 22336 22040 22342 22092
rect 20809 22015 20867 22021
rect 20809 21981 20821 22015
rect 20855 21981 20867 22015
rect 20809 21975 20867 21981
rect 17190 21916 18184 21944
rect 12728 21848 13032 21876
rect 13081 21879 13139 21885
rect 13081 21845 13093 21879
rect 13127 21876 13139 21879
rect 13170 21876 13176 21888
rect 13127 21848 13176 21876
rect 13127 21845 13139 21848
rect 13081 21839 13139 21845
rect 13170 21836 13176 21848
rect 13228 21836 13234 21888
rect 13630 21836 13636 21888
rect 13688 21876 13694 21888
rect 14277 21879 14335 21885
rect 14277 21876 14289 21879
rect 13688 21848 14289 21876
rect 13688 21836 13694 21848
rect 14277 21845 14289 21848
rect 14323 21845 14335 21879
rect 14277 21839 14335 21845
rect 14645 21879 14703 21885
rect 14645 21845 14657 21879
rect 14691 21876 14703 21879
rect 14918 21876 14924 21888
rect 14691 21848 14924 21876
rect 14691 21845 14703 21848
rect 14645 21839 14703 21845
rect 14918 21836 14924 21848
rect 14976 21836 14982 21888
rect 15654 21836 15660 21888
rect 15712 21836 15718 21888
rect 16298 21836 16304 21888
rect 16356 21876 16362 21888
rect 16758 21876 16764 21888
rect 16356 21848 16764 21876
rect 16356 21836 16362 21848
rect 16758 21836 16764 21848
rect 16816 21876 16822 21888
rect 17190 21876 17218 21916
rect 16816 21848 17218 21876
rect 16816 21836 16822 21848
rect 17310 21836 17316 21888
rect 17368 21876 17374 21888
rect 17405 21879 17463 21885
rect 17405 21876 17417 21879
rect 17368 21848 17417 21876
rect 17368 21836 17374 21848
rect 17405 21845 17417 21848
rect 17451 21845 17463 21879
rect 17405 21839 17463 21845
rect 17770 21836 17776 21888
rect 17828 21836 17834 21888
rect 18046 21836 18052 21888
rect 18104 21836 18110 21888
rect 18156 21876 18184 21916
rect 18598 21904 18604 21956
rect 18656 21904 18662 21956
rect 18708 21876 18736 21972
rect 19490 21947 19548 21953
rect 19490 21944 19502 21947
rect 18892 21916 19502 21944
rect 18892 21885 18920 21916
rect 19490 21913 19502 21916
rect 19536 21913 19548 21947
rect 19490 21907 19548 21913
rect 18156 21848 18736 21876
rect 18877 21879 18935 21885
rect 18877 21845 18889 21879
rect 18923 21845 18935 21879
rect 18877 21839 18935 21845
rect 20162 21836 20168 21888
rect 20220 21876 20226 21888
rect 20625 21879 20683 21885
rect 20625 21876 20637 21879
rect 20220 21848 20637 21876
rect 20220 21836 20226 21848
rect 20625 21845 20637 21848
rect 20671 21845 20683 21879
rect 20625 21839 20683 21845
rect 20714 21836 20720 21888
rect 20772 21876 20778 21888
rect 20901 21879 20959 21885
rect 20901 21876 20913 21879
rect 20772 21848 20913 21876
rect 20772 21836 20778 21848
rect 20901 21845 20913 21848
rect 20947 21845 20959 21879
rect 20901 21839 20959 21845
rect 1104 21786 27876 21808
rect 1104 21734 4874 21786
rect 4926 21734 4938 21786
rect 4990 21734 5002 21786
rect 5054 21734 5066 21786
rect 5118 21734 5130 21786
rect 5182 21734 27876 21786
rect 1104 21712 27876 21734
rect 5442 21632 5448 21684
rect 5500 21632 5506 21684
rect 7098 21672 7104 21684
rect 5828 21644 7104 21672
rect 5258 21604 5264 21616
rect 5000 21576 5264 21604
rect 842 21496 848 21548
rect 900 21536 906 21548
rect 1397 21539 1455 21545
rect 1397 21536 1409 21539
rect 900 21508 1409 21536
rect 900 21496 906 21508
rect 1397 21505 1409 21508
rect 1443 21505 1455 21539
rect 1397 21499 1455 21505
rect 2314 21496 2320 21548
rect 2372 21496 2378 21548
rect 2584 21539 2642 21545
rect 2584 21505 2596 21539
rect 2630 21536 2642 21539
rect 2866 21536 2872 21548
rect 2630 21508 2872 21536
rect 2630 21505 2642 21508
rect 2584 21499 2642 21505
rect 2866 21496 2872 21508
rect 2924 21496 2930 21548
rect 5000 21545 5028 21576
rect 5258 21564 5264 21576
rect 5316 21564 5322 21616
rect 5828 21545 5856 21644
rect 7098 21632 7104 21644
rect 7156 21632 7162 21684
rect 7190 21632 7196 21684
rect 7248 21632 7254 21684
rect 7466 21672 7472 21684
rect 7392 21644 7472 21672
rect 6914 21604 6920 21616
rect 6656 21576 6920 21604
rect 6656 21545 6684 21576
rect 6914 21564 6920 21576
rect 6972 21564 6978 21616
rect 4985 21539 5043 21545
rect 4985 21505 4997 21539
rect 5031 21505 5043 21539
rect 4985 21499 5043 21505
rect 5078 21539 5136 21545
rect 5078 21505 5090 21539
rect 5124 21505 5136 21539
rect 5078 21499 5136 21505
rect 5813 21539 5871 21545
rect 5813 21505 5825 21539
rect 5859 21505 5871 21539
rect 5813 21499 5871 21505
rect 6641 21539 6699 21545
rect 6641 21505 6653 21539
rect 6687 21505 6699 21539
rect 6641 21499 6699 21505
rect 3973 21471 4031 21477
rect 3973 21437 3985 21471
rect 4019 21437 4031 21471
rect 3973 21431 4031 21437
rect 3697 21403 3755 21409
rect 3697 21369 3709 21403
rect 3743 21400 3755 21403
rect 3988 21400 4016 21431
rect 4798 21428 4804 21480
rect 4856 21468 4862 21480
rect 5092 21468 5120 21499
rect 7098 21496 7104 21548
rect 7156 21496 7162 21548
rect 7190 21496 7196 21548
rect 7248 21536 7254 21548
rect 7285 21539 7343 21545
rect 7285 21536 7297 21539
rect 7248 21508 7297 21536
rect 7248 21496 7254 21508
rect 7285 21505 7297 21508
rect 7331 21505 7343 21539
rect 7285 21499 7343 21505
rect 4856 21440 5120 21468
rect 4856 21428 4862 21440
rect 5258 21428 5264 21480
rect 5316 21468 5322 21480
rect 5353 21471 5411 21477
rect 5353 21468 5365 21471
rect 5316 21440 5365 21468
rect 5316 21428 5322 21440
rect 5353 21437 5365 21440
rect 5399 21468 5411 21471
rect 5629 21471 5687 21477
rect 5629 21468 5641 21471
rect 5399 21440 5641 21468
rect 5399 21437 5411 21440
rect 5353 21431 5411 21437
rect 5629 21437 5641 21440
rect 5675 21437 5687 21471
rect 5629 21431 5687 21437
rect 5442 21400 5448 21412
rect 3743 21372 5448 21400
rect 3743 21369 3755 21372
rect 3697 21363 3755 21369
rect 5442 21360 5448 21372
rect 5500 21360 5506 21412
rect 5644 21400 5672 21431
rect 5718 21428 5724 21480
rect 5776 21428 5782 21480
rect 5905 21471 5963 21477
rect 5905 21437 5917 21471
rect 5951 21468 5963 21471
rect 6457 21471 6515 21477
rect 6457 21468 6469 21471
rect 5951 21440 6469 21468
rect 5951 21437 5963 21440
rect 5905 21431 5963 21437
rect 6457 21437 6469 21440
rect 6503 21437 6515 21471
rect 6457 21431 6515 21437
rect 6733 21471 6791 21477
rect 6733 21437 6745 21471
rect 6779 21437 6791 21471
rect 6733 21431 6791 21437
rect 6825 21471 6883 21477
rect 6825 21437 6837 21471
rect 6871 21437 6883 21471
rect 6825 21431 6883 21437
rect 6638 21400 6644 21412
rect 5644 21372 6644 21400
rect 6638 21360 6644 21372
rect 6696 21360 6702 21412
rect 1578 21292 1584 21344
rect 1636 21292 1642 21344
rect 4525 21335 4583 21341
rect 4525 21301 4537 21335
rect 4571 21332 4583 21335
rect 4614 21332 4620 21344
rect 4571 21304 4620 21332
rect 4571 21301 4583 21304
rect 4525 21295 4583 21301
rect 4614 21292 4620 21304
rect 4672 21292 4678 21344
rect 6748 21332 6776 21431
rect 6840 21400 6868 21431
rect 6914 21428 6920 21480
rect 6972 21428 6978 21480
rect 7098 21400 7104 21412
rect 6840 21372 7104 21400
rect 7098 21360 7104 21372
rect 7156 21400 7162 21412
rect 7392 21400 7420 21644
rect 7466 21632 7472 21644
rect 7524 21632 7530 21684
rect 7834 21632 7840 21684
rect 7892 21672 7898 21684
rect 8849 21675 8907 21681
rect 7892 21644 8800 21672
rect 7892 21632 7898 21644
rect 7736 21607 7794 21613
rect 7736 21573 7748 21607
rect 7782 21604 7794 21607
rect 7926 21604 7932 21616
rect 7782 21576 7932 21604
rect 7782 21573 7794 21576
rect 7736 21567 7794 21573
rect 7926 21564 7932 21576
rect 7984 21564 7990 21616
rect 7466 21496 7472 21548
rect 7524 21536 7530 21548
rect 8018 21536 8024 21548
rect 7524 21508 8024 21536
rect 7524 21496 7530 21508
rect 8018 21496 8024 21508
rect 8076 21496 8082 21548
rect 8772 21468 8800 21644
rect 8849 21641 8861 21675
rect 8895 21641 8907 21675
rect 8849 21635 8907 21641
rect 8864 21536 8892 21635
rect 13630 21632 13636 21684
rect 13688 21672 13694 21684
rect 13909 21675 13967 21681
rect 13909 21672 13921 21675
rect 13688 21644 13921 21672
rect 13688 21632 13694 21644
rect 13909 21641 13921 21644
rect 13955 21641 13967 21675
rect 13909 21635 13967 21641
rect 14642 21632 14648 21684
rect 14700 21672 14706 21684
rect 14700 21644 15332 21672
rect 14700 21632 14706 21644
rect 15304 21616 15332 21644
rect 15562 21632 15568 21684
rect 15620 21672 15626 21684
rect 15620 21644 15700 21672
rect 15620 21632 15626 21644
rect 12158 21564 12164 21616
rect 12216 21564 12222 21616
rect 12774 21607 12832 21613
rect 12774 21604 12786 21607
rect 12468 21576 12786 21604
rect 8941 21539 8999 21545
rect 8941 21536 8953 21539
rect 8864 21508 8953 21536
rect 8941 21505 8953 21508
rect 8987 21505 8999 21539
rect 8941 21499 8999 21505
rect 11514 21496 11520 21548
rect 11572 21536 11578 21548
rect 11885 21539 11943 21545
rect 11885 21536 11897 21539
rect 11572 21508 11897 21536
rect 11572 21496 11578 21508
rect 11885 21505 11897 21508
rect 11931 21505 11943 21539
rect 11885 21499 11943 21505
rect 12069 21539 12127 21545
rect 12069 21505 12081 21539
rect 12115 21505 12127 21539
rect 12069 21499 12127 21505
rect 12084 21468 12112 21499
rect 12250 21496 12256 21548
rect 12308 21496 12314 21548
rect 8772 21440 12112 21468
rect 7156 21372 7420 21400
rect 7156 21360 7162 21372
rect 8938 21360 8944 21412
rect 8996 21400 9002 21412
rect 11882 21400 11888 21412
rect 8996 21372 11888 21400
rect 8996 21360 9002 21372
rect 11882 21360 11888 21372
rect 11940 21360 11946 21412
rect 7834 21332 7840 21344
rect 6748 21304 7840 21332
rect 7834 21292 7840 21304
rect 7892 21332 7898 21344
rect 9033 21335 9091 21341
rect 9033 21332 9045 21335
rect 7892 21304 9045 21332
rect 7892 21292 7898 21304
rect 9033 21301 9045 21304
rect 9079 21301 9091 21335
rect 12084 21332 12112 21440
rect 12468 21409 12496 21576
rect 12774 21573 12786 21576
rect 12820 21573 12832 21607
rect 12774 21567 12832 21573
rect 13354 21564 13360 21616
rect 13412 21604 13418 21616
rect 14553 21607 14611 21613
rect 14553 21604 14565 21607
rect 13412 21576 14565 21604
rect 13412 21564 13418 21576
rect 14553 21573 14565 21576
rect 14599 21573 14611 21607
rect 14553 21567 14611 21573
rect 14769 21607 14827 21613
rect 14769 21573 14781 21607
rect 14815 21604 14827 21607
rect 14815 21576 14964 21604
rect 14815 21573 14827 21576
rect 14769 21567 14827 21573
rect 12526 21496 12532 21548
rect 12584 21496 12590 21548
rect 14568 21468 14596 21567
rect 14936 21548 14964 21576
rect 15286 21564 15292 21616
rect 15344 21564 15350 21616
rect 15672 21604 15700 21644
rect 15838 21632 15844 21684
rect 15896 21632 15902 21684
rect 16666 21632 16672 21684
rect 16724 21632 16730 21684
rect 16776 21644 17448 21672
rect 16022 21604 16028 21616
rect 15672 21576 16028 21604
rect 16022 21564 16028 21576
rect 16080 21604 16086 21616
rect 16390 21604 16396 21616
rect 16080 21576 16396 21604
rect 16080 21564 16086 21576
rect 16390 21564 16396 21576
rect 16448 21564 16454 21616
rect 14918 21496 14924 21548
rect 14976 21536 14982 21548
rect 15013 21539 15071 21545
rect 15013 21536 15025 21539
rect 14976 21508 15025 21536
rect 14976 21496 14982 21508
rect 15013 21505 15025 21508
rect 15059 21505 15071 21539
rect 15013 21499 15071 21505
rect 15105 21539 15163 21545
rect 15105 21505 15117 21539
rect 15151 21505 15163 21539
rect 15105 21499 15163 21505
rect 15120 21468 15148 21499
rect 15378 21496 15384 21548
rect 15436 21496 15442 21548
rect 15519 21539 15577 21545
rect 15519 21505 15531 21539
rect 15565 21536 15577 21539
rect 15654 21536 15660 21548
rect 15565 21508 15660 21536
rect 15565 21505 15577 21508
rect 15519 21499 15577 21505
rect 15654 21496 15660 21508
rect 15712 21496 15718 21548
rect 15838 21496 15844 21548
rect 15896 21496 15902 21548
rect 16114 21496 16120 21548
rect 16172 21536 16178 21548
rect 16776 21536 16804 21644
rect 16945 21607 17003 21613
rect 16945 21573 16957 21607
rect 16991 21604 17003 21607
rect 17310 21604 17316 21616
rect 16991 21576 17316 21604
rect 16991 21573 17003 21576
rect 16945 21567 17003 21573
rect 17310 21564 17316 21576
rect 17368 21564 17374 21616
rect 16172 21508 16804 21536
rect 16853 21539 16911 21545
rect 16172 21496 16178 21508
rect 16853 21505 16865 21539
rect 16899 21505 16911 21539
rect 16853 21499 16911 21505
rect 16022 21468 16028 21480
rect 14568 21440 16028 21468
rect 16022 21428 16028 21440
rect 16080 21428 16086 21480
rect 16301 21471 16359 21477
rect 16301 21437 16313 21471
rect 16347 21468 16359 21471
rect 16390 21468 16396 21480
rect 16347 21440 16396 21468
rect 16347 21437 16359 21440
rect 16301 21431 16359 21437
rect 16390 21428 16396 21440
rect 16448 21428 16454 21480
rect 12437 21403 12496 21409
rect 12437 21369 12449 21403
rect 12483 21372 12496 21403
rect 14550 21400 14556 21412
rect 13832 21372 14556 21400
rect 12483 21369 12495 21372
rect 12437 21363 12495 21369
rect 12710 21332 12716 21344
rect 12084 21304 12716 21332
rect 9033 21295 9091 21301
rect 12710 21292 12716 21304
rect 12768 21332 12774 21344
rect 13832 21332 13860 21372
rect 14550 21360 14556 21372
rect 14608 21360 14614 21412
rect 15289 21403 15347 21409
rect 15289 21369 15301 21403
rect 15335 21400 15347 21403
rect 16868 21400 16896 21499
rect 17034 21496 17040 21548
rect 17092 21496 17098 21548
rect 17218 21545 17224 21548
rect 17175 21539 17224 21545
rect 17175 21505 17187 21539
rect 17221 21505 17224 21539
rect 17175 21499 17224 21505
rect 17218 21496 17224 21499
rect 17276 21496 17282 21548
rect 17420 21545 17448 21644
rect 18414 21632 18420 21684
rect 18472 21632 18478 21684
rect 18598 21632 18604 21684
rect 18656 21672 18662 21684
rect 19613 21675 19671 21681
rect 19613 21672 19625 21675
rect 18656 21644 19625 21672
rect 18656 21632 18662 21644
rect 19613 21641 19625 21644
rect 19659 21641 19671 21675
rect 19613 21635 19671 21641
rect 21821 21675 21879 21681
rect 21821 21641 21833 21675
rect 21867 21641 21879 21675
rect 22554 21672 22560 21684
rect 21821 21635 21879 21641
rect 22066 21644 22560 21672
rect 17494 21564 17500 21616
rect 17552 21604 17558 21616
rect 21836 21604 21864 21635
rect 22066 21604 22094 21644
rect 22554 21632 22560 21644
rect 22612 21632 22618 21684
rect 22649 21675 22707 21681
rect 22649 21641 22661 21675
rect 22695 21641 22707 21675
rect 22649 21635 22707 21641
rect 17552 21576 21864 21604
rect 21928 21576 22094 21604
rect 17552 21564 17558 21576
rect 17405 21539 17463 21545
rect 17405 21505 17417 21539
rect 17451 21505 17463 21539
rect 17957 21539 18015 21545
rect 17957 21536 17969 21539
rect 17405 21499 17463 21505
rect 17696 21508 17969 21536
rect 17313 21471 17371 21477
rect 17313 21437 17325 21471
rect 17359 21468 17371 21471
rect 17586 21468 17592 21480
rect 17359 21440 17592 21468
rect 17359 21437 17371 21440
rect 17313 21431 17371 21437
rect 17586 21428 17592 21440
rect 17644 21428 17650 21480
rect 17497 21403 17555 21409
rect 17497 21400 17509 21403
rect 15335 21372 16804 21400
rect 16868 21372 17509 21400
rect 15335 21369 15347 21372
rect 15289 21363 15347 21369
rect 12768 21304 13860 21332
rect 12768 21292 12774 21304
rect 13906 21292 13912 21344
rect 13964 21332 13970 21344
rect 14642 21332 14648 21344
rect 13964 21304 14648 21332
rect 13964 21292 13970 21304
rect 14642 21292 14648 21304
rect 14700 21332 14706 21344
rect 14737 21335 14795 21341
rect 14737 21332 14749 21335
rect 14700 21304 14749 21332
rect 14700 21292 14706 21304
rect 14737 21301 14749 21304
rect 14783 21301 14795 21335
rect 14737 21295 14795 21301
rect 14921 21335 14979 21341
rect 14921 21301 14933 21335
rect 14967 21332 14979 21335
rect 15102 21332 15108 21344
rect 14967 21304 15108 21332
rect 14967 21301 14979 21304
rect 14921 21295 14979 21301
rect 15102 21292 15108 21304
rect 15160 21292 15166 21344
rect 15654 21292 15660 21344
rect 15712 21332 15718 21344
rect 15933 21335 15991 21341
rect 15933 21332 15945 21335
rect 15712 21304 15945 21332
rect 15712 21292 15718 21304
rect 15933 21301 15945 21304
rect 15979 21301 15991 21335
rect 16776 21332 16804 21372
rect 17497 21369 17509 21372
rect 17543 21369 17555 21403
rect 17497 21363 17555 21369
rect 17696 21332 17724 21508
rect 17957 21505 17969 21508
rect 18003 21505 18015 21539
rect 17957 21499 18015 21505
rect 18248 21508 18552 21536
rect 18046 21428 18052 21480
rect 18104 21428 18110 21480
rect 16776 21304 17724 21332
rect 15933 21295 15991 21301
rect 17862 21292 17868 21344
rect 17920 21332 17926 21344
rect 18141 21335 18199 21341
rect 18141 21332 18153 21335
rect 17920 21304 18153 21332
rect 17920 21292 17926 21304
rect 18141 21301 18153 21304
rect 18187 21332 18199 21335
rect 18248 21332 18276 21508
rect 18417 21471 18475 21477
rect 18417 21468 18429 21471
rect 18340 21440 18429 21468
rect 18340 21409 18368 21440
rect 18417 21437 18429 21440
rect 18463 21437 18475 21471
rect 18524 21468 18552 21508
rect 18690 21496 18696 21548
rect 18748 21496 18754 21548
rect 20162 21496 20168 21548
rect 20220 21536 20226 21548
rect 21928 21536 21956 21576
rect 22186 21564 22192 21616
rect 22244 21604 22250 21616
rect 22664 21604 22692 21635
rect 22738 21632 22744 21684
rect 22796 21672 22802 21684
rect 22796 21644 23060 21672
rect 22796 21632 22802 21644
rect 23032 21616 23060 21644
rect 22244 21576 22692 21604
rect 22244 21564 22250 21576
rect 20220 21508 21956 21536
rect 20220 21496 20226 21508
rect 22094 21496 22100 21548
rect 22152 21496 22158 21548
rect 20806 21468 20812 21480
rect 18524 21440 20812 21468
rect 18417 21431 18475 21437
rect 20806 21428 20812 21440
rect 20864 21428 20870 21480
rect 22005 21471 22063 21477
rect 22005 21437 22017 21471
rect 22051 21468 22063 21471
rect 22296 21468 22324 21576
rect 23014 21564 23020 21616
rect 23072 21604 23078 21616
rect 23072 21576 23704 21604
rect 23072 21564 23078 21576
rect 22557 21539 22615 21545
rect 22557 21505 22569 21539
rect 22603 21536 22615 21539
rect 22646 21536 22652 21548
rect 22603 21508 22652 21536
rect 22603 21505 22615 21508
rect 22557 21499 22615 21505
rect 22646 21496 22652 21508
rect 22704 21496 22710 21548
rect 22738 21496 22744 21548
rect 22796 21496 22802 21548
rect 23382 21496 23388 21548
rect 23440 21537 23446 21548
rect 23676 21545 23704 21576
rect 23661 21539 23719 21545
rect 23440 21509 23520 21537
rect 23440 21496 23446 21509
rect 22051 21440 22324 21468
rect 22051 21437 22063 21440
rect 22005 21431 22063 21437
rect 22370 21428 22376 21480
rect 22428 21428 22434 21480
rect 22462 21428 22468 21480
rect 22520 21428 22526 21480
rect 23198 21428 23204 21480
rect 23256 21468 23262 21480
rect 23293 21471 23351 21477
rect 23293 21468 23305 21471
rect 23256 21440 23305 21468
rect 23256 21428 23262 21440
rect 23293 21437 23305 21440
rect 23339 21437 23351 21471
rect 23492 21468 23520 21509
rect 23661 21505 23673 21539
rect 23707 21505 23719 21539
rect 23661 21499 23719 21505
rect 23753 21471 23811 21477
rect 23753 21468 23765 21471
rect 23492 21440 23765 21468
rect 23293 21431 23351 21437
rect 23753 21437 23765 21440
rect 23799 21437 23811 21471
rect 23753 21431 23811 21437
rect 18325 21403 18383 21409
rect 18325 21369 18337 21403
rect 18371 21369 18383 21403
rect 18325 21363 18383 21369
rect 18506 21360 18512 21412
rect 18564 21400 18570 21412
rect 20898 21400 20904 21412
rect 18564 21372 20904 21400
rect 18564 21360 18570 21372
rect 20898 21360 20904 21372
rect 20956 21360 20962 21412
rect 23017 21403 23075 21409
rect 23017 21400 23029 21403
rect 22066 21372 23029 21400
rect 18187 21304 18276 21332
rect 18187 21301 18199 21304
rect 18141 21295 18199 21301
rect 18598 21292 18604 21344
rect 18656 21292 18662 21344
rect 20806 21292 20812 21344
rect 20864 21332 20870 21344
rect 22066 21332 22094 21372
rect 23017 21369 23029 21372
rect 23063 21369 23075 21403
rect 23017 21363 23075 21369
rect 20864 21304 22094 21332
rect 20864 21292 20870 21304
rect 1104 21242 27876 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 27876 21242
rect 1104 21168 27876 21190
rect 2866 21088 2872 21140
rect 2924 21088 2930 21140
rect 5718 21088 5724 21140
rect 5776 21128 5782 21140
rect 5813 21131 5871 21137
rect 5813 21128 5825 21131
rect 5776 21100 5825 21128
rect 5776 21088 5782 21100
rect 5813 21097 5825 21100
rect 5859 21097 5871 21131
rect 6822 21128 6828 21140
rect 5813 21091 5871 21097
rect 6656 21100 6828 21128
rect 6656 21069 6684 21100
rect 6822 21088 6828 21100
rect 6880 21088 6886 21140
rect 8662 21088 8668 21140
rect 8720 21128 8726 21140
rect 8720 21100 10364 21128
rect 8720 21088 8726 21100
rect 2777 21063 2835 21069
rect 2777 21029 2789 21063
rect 2823 21060 2835 21063
rect 6641 21063 6699 21069
rect 2823 21032 3464 21060
rect 2823 21029 2835 21032
rect 2777 21023 2835 21029
rect 3436 20933 3464 21032
rect 5368 21032 5948 21060
rect 5368 20936 5396 21032
rect 5442 20952 5448 21004
rect 5500 20952 5506 21004
rect 5644 20964 5856 20992
rect 1397 20927 1455 20933
rect 1397 20893 1409 20927
rect 1443 20893 1455 20927
rect 1397 20887 1455 20893
rect 1664 20927 1722 20933
rect 1664 20893 1676 20927
rect 1710 20893 1722 20927
rect 1664 20887 1722 20893
rect 3421 20927 3479 20933
rect 3421 20893 3433 20927
rect 3467 20893 3479 20927
rect 3421 20887 3479 20893
rect 3789 20927 3847 20933
rect 3789 20893 3801 20927
rect 3835 20893 3847 20927
rect 3789 20887 3847 20893
rect 1412 20788 1440 20887
rect 1578 20816 1584 20868
rect 1636 20856 1642 20868
rect 1688 20856 1716 20887
rect 3804 20856 3832 20887
rect 5258 20884 5264 20936
rect 5316 20884 5322 20936
rect 5350 20884 5356 20936
rect 5408 20884 5414 20936
rect 5644 20933 5672 20964
rect 5629 20927 5687 20933
rect 5629 20893 5641 20927
rect 5675 20893 5687 20927
rect 5629 20887 5687 20893
rect 5721 20927 5779 20933
rect 5721 20893 5733 20927
rect 5767 20893 5779 20927
rect 5721 20887 5779 20893
rect 1636 20828 1716 20856
rect 2792 20828 3832 20856
rect 4056 20859 4114 20865
rect 1636 20816 1642 20828
rect 2792 20800 2820 20828
rect 4056 20825 4068 20859
rect 4102 20856 4114 20859
rect 4614 20856 4620 20868
rect 4102 20828 4620 20856
rect 4102 20825 4114 20828
rect 4056 20819 4114 20825
rect 4614 20816 4620 20828
rect 4672 20856 4678 20868
rect 5736 20856 5764 20887
rect 4672 20828 5764 20856
rect 5828 20856 5856 20964
rect 5920 20933 5948 21032
rect 6641 21029 6653 21063
rect 6687 21029 6699 21063
rect 6641 21023 6699 21029
rect 6730 21020 6736 21072
rect 6788 21020 6794 21072
rect 10336 21060 10364 21100
rect 10594 21088 10600 21140
rect 10652 21128 10658 21140
rect 10781 21131 10839 21137
rect 10781 21128 10793 21131
rect 10652 21100 10793 21128
rect 10652 21088 10658 21100
rect 10781 21097 10793 21100
rect 10827 21128 10839 21131
rect 10962 21128 10968 21140
rect 10827 21100 10968 21128
rect 10827 21097 10839 21100
rect 10781 21091 10839 21097
rect 10962 21088 10968 21100
rect 11020 21088 11026 21140
rect 15013 21131 15071 21137
rect 15013 21097 15025 21131
rect 15059 21128 15071 21131
rect 15470 21128 15476 21140
rect 15059 21100 15476 21128
rect 15059 21097 15071 21100
rect 15013 21091 15071 21097
rect 15470 21088 15476 21100
rect 15528 21088 15534 21140
rect 15562 21088 15568 21140
rect 15620 21128 15626 21140
rect 15930 21128 15936 21140
rect 15620 21100 15936 21128
rect 15620 21088 15626 21100
rect 15930 21088 15936 21100
rect 15988 21088 15994 21140
rect 16022 21088 16028 21140
rect 16080 21128 16086 21140
rect 17494 21128 17500 21140
rect 16080 21100 17500 21128
rect 16080 21088 16086 21100
rect 17494 21088 17500 21100
rect 17552 21088 17558 21140
rect 17586 21088 17592 21140
rect 17644 21088 17650 21140
rect 18509 21131 18567 21137
rect 18509 21097 18521 21131
rect 18555 21128 18567 21131
rect 18598 21128 18604 21140
rect 18555 21100 18604 21128
rect 18555 21097 18567 21100
rect 18509 21091 18567 21097
rect 18598 21088 18604 21100
rect 18656 21088 18662 21140
rect 18690 21088 18696 21140
rect 18748 21128 18754 21140
rect 19245 21131 19303 21137
rect 19245 21128 19257 21131
rect 18748 21100 19257 21128
rect 18748 21088 18754 21100
rect 19245 21097 19257 21100
rect 19291 21097 19303 21131
rect 19245 21091 19303 21097
rect 19794 21088 19800 21140
rect 19852 21128 19858 21140
rect 20622 21128 20628 21140
rect 19852 21100 20628 21128
rect 19852 21088 19858 21100
rect 20622 21088 20628 21100
rect 20680 21128 20686 21140
rect 21358 21128 21364 21140
rect 20680 21100 21364 21128
rect 20680 21088 20686 21100
rect 21358 21088 21364 21100
rect 21416 21088 21422 21140
rect 21545 21131 21603 21137
rect 21545 21097 21557 21131
rect 21591 21128 21603 21131
rect 22094 21128 22100 21140
rect 21591 21100 22100 21128
rect 21591 21097 21603 21100
rect 21545 21091 21603 21097
rect 22094 21088 22100 21100
rect 22152 21088 22158 21140
rect 22646 21088 22652 21140
rect 22704 21088 22710 21140
rect 22830 21088 22836 21140
rect 22888 21128 22894 21140
rect 23290 21128 23296 21140
rect 22888 21100 23296 21128
rect 22888 21088 22894 21100
rect 23290 21088 23296 21100
rect 23348 21088 23354 21140
rect 12802 21060 12808 21072
rect 10336 21032 12808 21060
rect 12802 21020 12808 21032
rect 12860 21060 12866 21072
rect 14090 21060 14096 21072
rect 12860 21032 14096 21060
rect 12860 21020 12866 21032
rect 14090 21020 14096 21032
rect 14148 21020 14154 21072
rect 15749 21063 15807 21069
rect 15749 21029 15761 21063
rect 15795 21060 15807 21063
rect 16114 21060 16120 21072
rect 15795 21032 16120 21060
rect 15795 21029 15807 21032
rect 15749 21023 15807 21029
rect 16114 21020 16120 21032
rect 16172 21020 16178 21072
rect 21269 21063 21327 21069
rect 21269 21060 21281 21063
rect 17420 21032 21281 21060
rect 7190 20992 7196 21004
rect 6564 20964 7196 20992
rect 6564 20933 6592 20964
rect 7190 20952 7196 20964
rect 7248 20952 7254 21004
rect 8018 20952 8024 21004
rect 8076 20992 8082 21004
rect 9398 20992 9404 21004
rect 8076 20964 9404 20992
rect 8076 20952 8082 20964
rect 9398 20952 9404 20964
rect 9456 20952 9462 21004
rect 13814 20952 13820 21004
rect 13872 20992 13878 21004
rect 14918 20992 14924 21004
rect 13872 20964 14924 20992
rect 13872 20952 13878 20964
rect 14918 20952 14924 20964
rect 14976 20952 14982 21004
rect 15286 20952 15292 21004
rect 15344 20992 15350 21004
rect 17420 21001 17448 21032
rect 17313 20995 17371 21001
rect 17313 20992 17325 20995
rect 15344 20964 17325 20992
rect 15344 20952 15350 20964
rect 17313 20961 17325 20964
rect 17359 20961 17371 20995
rect 17313 20955 17371 20961
rect 17405 20995 17463 21001
rect 17405 20961 17417 20995
rect 17451 20961 17463 20995
rect 17405 20955 17463 20961
rect 5905 20927 5963 20933
rect 5905 20893 5917 20927
rect 5951 20893 5963 20927
rect 5905 20887 5963 20893
rect 6549 20927 6607 20933
rect 6549 20893 6561 20927
rect 6595 20893 6607 20927
rect 6549 20887 6607 20893
rect 6825 20927 6883 20933
rect 6825 20893 6837 20927
rect 6871 20924 6883 20927
rect 7377 20927 7435 20933
rect 7377 20924 7389 20927
rect 6871 20896 7389 20924
rect 6871 20893 6883 20896
rect 6825 20887 6883 20893
rect 7377 20893 7389 20896
rect 7423 20893 7435 20927
rect 7377 20887 7435 20893
rect 7558 20884 7564 20936
rect 7616 20884 7622 20936
rect 7834 20884 7840 20936
rect 7892 20884 7898 20936
rect 8941 20927 8999 20933
rect 8941 20893 8953 20927
rect 8987 20893 8999 20927
rect 8941 20887 8999 20893
rect 9125 20927 9183 20933
rect 9125 20893 9137 20927
rect 9171 20924 9183 20927
rect 9306 20924 9312 20936
rect 9171 20896 9312 20924
rect 9171 20893 9183 20896
rect 9125 20887 9183 20893
rect 6365 20859 6423 20865
rect 6365 20856 6377 20859
rect 5828 20828 6377 20856
rect 4672 20816 4678 20828
rect 6365 20825 6377 20828
rect 6411 20825 6423 20859
rect 6365 20819 6423 20825
rect 7098 20816 7104 20868
rect 7156 20856 7162 20868
rect 7745 20859 7803 20865
rect 7745 20856 7757 20859
rect 7156 20828 7757 20856
rect 7156 20816 7162 20828
rect 7745 20825 7757 20828
rect 7791 20825 7803 20859
rect 7745 20819 7803 20825
rect 8956 20856 8984 20887
rect 9306 20884 9312 20896
rect 9364 20884 9370 20936
rect 15746 20924 15752 20936
rect 14844 20896 15752 20924
rect 9674 20865 9680 20868
rect 8956 20828 9168 20856
rect 2774 20788 2780 20800
rect 1412 20760 2780 20788
rect 2774 20748 2780 20760
rect 2832 20748 2838 20800
rect 5169 20791 5227 20797
rect 5169 20757 5181 20791
rect 5215 20788 5227 20791
rect 5258 20788 5264 20800
rect 5215 20760 5264 20788
rect 5215 20757 5227 20760
rect 5169 20751 5227 20757
rect 5258 20748 5264 20760
rect 5316 20748 5322 20800
rect 5537 20791 5595 20797
rect 5537 20757 5549 20791
rect 5583 20788 5595 20791
rect 6270 20788 6276 20800
rect 5583 20760 6276 20788
rect 5583 20757 5595 20760
rect 5537 20751 5595 20757
rect 6270 20748 6276 20760
rect 6328 20748 6334 20800
rect 7558 20748 7564 20800
rect 7616 20788 7622 20800
rect 8956 20788 8984 20828
rect 7616 20760 8984 20788
rect 7616 20748 7622 20760
rect 9030 20748 9036 20800
rect 9088 20748 9094 20800
rect 9140 20788 9168 20828
rect 9668 20819 9680 20865
rect 9674 20816 9680 20819
rect 9732 20816 9738 20868
rect 13998 20816 14004 20868
rect 14056 20856 14062 20868
rect 14844 20865 14872 20896
rect 15746 20884 15752 20896
rect 15804 20884 15810 20936
rect 15838 20884 15844 20936
rect 15896 20924 15902 20936
rect 17328 20924 17356 20955
rect 17494 20952 17500 21004
rect 17552 20992 17558 21004
rect 18325 20995 18383 21001
rect 17552 20964 18276 20992
rect 17552 20952 17558 20964
rect 18046 20924 18052 20936
rect 15896 20896 17264 20924
rect 17328 20896 18052 20924
rect 15896 20884 15902 20896
rect 15102 20865 15108 20868
rect 14829 20859 14887 20865
rect 14829 20856 14841 20859
rect 14056 20828 14841 20856
rect 14056 20816 14062 20828
rect 14829 20825 14841 20828
rect 14875 20825 14887 20859
rect 14829 20819 14887 20825
rect 15045 20859 15108 20865
rect 15045 20825 15057 20859
rect 15091 20825 15108 20859
rect 15045 20819 15108 20825
rect 15102 20816 15108 20819
rect 15160 20856 15166 20868
rect 15160 20828 15960 20856
rect 15160 20816 15166 20828
rect 10134 20788 10140 20800
rect 9140 20760 10140 20788
rect 10134 20748 10140 20760
rect 10192 20788 10198 20800
rect 10778 20788 10784 20800
rect 10192 20760 10784 20788
rect 10192 20748 10198 20760
rect 10778 20748 10784 20760
rect 10836 20748 10842 20800
rect 12342 20748 12348 20800
rect 12400 20788 12406 20800
rect 14734 20788 14740 20800
rect 12400 20760 14740 20788
rect 12400 20748 12406 20760
rect 14734 20748 14740 20760
rect 14792 20748 14798 20800
rect 15197 20791 15255 20797
rect 15197 20757 15209 20791
rect 15243 20788 15255 20791
rect 15562 20788 15568 20800
rect 15243 20760 15568 20788
rect 15243 20757 15255 20760
rect 15197 20751 15255 20757
rect 15562 20748 15568 20760
rect 15620 20748 15626 20800
rect 15932 20797 15960 20828
rect 16022 20816 16028 20868
rect 16080 20856 16086 20868
rect 16117 20859 16175 20865
rect 16117 20856 16129 20859
rect 16080 20828 16129 20856
rect 16080 20816 16086 20828
rect 16117 20825 16129 20828
rect 16163 20825 16175 20859
rect 16117 20819 16175 20825
rect 15917 20791 15975 20797
rect 15917 20757 15929 20791
rect 15963 20788 15975 20791
rect 16298 20788 16304 20800
rect 15963 20760 16304 20788
rect 15963 20757 15975 20760
rect 15917 20751 15975 20757
rect 16298 20748 16304 20760
rect 16356 20748 16362 20800
rect 16942 20748 16948 20800
rect 17000 20748 17006 20800
rect 17236 20788 17264 20896
rect 18046 20884 18052 20896
rect 18104 20884 18110 20936
rect 18248 20933 18276 20964
rect 18325 20961 18337 20995
rect 18371 20992 18383 20995
rect 18877 20995 18935 21001
rect 18877 20992 18889 20995
rect 18371 20964 18889 20992
rect 18371 20961 18383 20964
rect 18325 20955 18383 20961
rect 18877 20961 18889 20964
rect 18923 20992 18935 20995
rect 18923 20964 19472 20992
rect 18923 20961 18935 20964
rect 18877 20955 18935 20961
rect 18233 20927 18291 20933
rect 18233 20893 18245 20927
rect 18279 20924 18291 20927
rect 18506 20924 18512 20936
rect 18279 20896 18512 20924
rect 18279 20893 18291 20896
rect 18233 20887 18291 20893
rect 18506 20884 18512 20896
rect 18564 20884 18570 20936
rect 18598 20884 18604 20936
rect 18656 20924 18662 20936
rect 18693 20927 18751 20933
rect 18693 20924 18705 20927
rect 18656 20896 18705 20924
rect 18656 20884 18662 20896
rect 18693 20893 18705 20896
rect 18739 20893 18751 20927
rect 18693 20887 18751 20893
rect 18785 20927 18843 20933
rect 18785 20893 18797 20927
rect 18831 20893 18843 20927
rect 18785 20887 18843 20893
rect 18800 20856 18828 20887
rect 18966 20884 18972 20936
rect 19024 20884 19030 20936
rect 19444 20933 19472 20964
rect 20272 20936 20300 21032
rect 21269 21029 21281 21032
rect 21315 21029 21327 21063
rect 21269 21023 21327 21029
rect 22462 21020 22468 21072
rect 22520 21060 22526 21072
rect 22557 21063 22615 21069
rect 22557 21060 22569 21063
rect 22520 21032 22569 21060
rect 22520 21020 22526 21032
rect 22557 21029 22569 21032
rect 22603 21029 22615 21063
rect 22557 21023 22615 21029
rect 22005 20995 22063 21001
rect 22005 20992 22017 20995
rect 21192 20964 22017 20992
rect 19429 20927 19487 20933
rect 19429 20893 19441 20927
rect 19475 20893 19487 20927
rect 19429 20887 19487 20893
rect 19521 20927 19579 20933
rect 19521 20893 19533 20927
rect 19567 20924 19579 20927
rect 19886 20924 19892 20936
rect 19567 20896 19892 20924
rect 19567 20893 19579 20896
rect 19521 20887 19579 20893
rect 19886 20884 19892 20896
rect 19944 20924 19950 20936
rect 20165 20927 20223 20933
rect 20165 20924 20177 20927
rect 19944 20896 20177 20924
rect 19944 20884 19950 20896
rect 20165 20893 20177 20896
rect 20211 20893 20223 20927
rect 20165 20887 20223 20893
rect 20254 20884 20260 20936
rect 20312 20884 20318 20936
rect 20530 20884 20536 20936
rect 20588 20884 20594 20936
rect 20622 20884 20628 20936
rect 20680 20884 20686 20936
rect 20717 20927 20775 20933
rect 20717 20893 20729 20927
rect 20763 20924 20775 20927
rect 20806 20924 20812 20936
rect 20763 20896 20812 20924
rect 20763 20893 20775 20896
rect 20717 20887 20775 20893
rect 19245 20859 19303 20865
rect 19245 20856 19257 20859
rect 18800 20828 19257 20856
rect 19245 20825 19257 20828
rect 19291 20856 19303 20859
rect 20349 20859 20407 20865
rect 19291 20828 20208 20856
rect 19291 20825 19303 20828
rect 19245 20819 19303 20825
rect 19981 20791 20039 20797
rect 19981 20788 19993 20791
rect 17236 20760 19993 20788
rect 19981 20757 19993 20760
rect 20027 20757 20039 20791
rect 20180 20788 20208 20828
rect 20349 20825 20361 20859
rect 20395 20856 20407 20859
rect 20438 20856 20444 20868
rect 20395 20828 20444 20856
rect 20395 20825 20407 20828
rect 20349 20819 20407 20825
rect 20438 20816 20444 20828
rect 20496 20816 20502 20868
rect 20732 20788 20760 20887
rect 20806 20884 20812 20896
rect 20864 20884 20870 20936
rect 20898 20884 20904 20936
rect 20956 20884 20962 20936
rect 21082 20884 21088 20936
rect 21140 20924 21146 20936
rect 21192 20933 21220 20964
rect 22005 20961 22017 20964
rect 22051 20961 22063 20995
rect 22005 20955 22063 20961
rect 21177 20927 21235 20933
rect 21177 20924 21189 20927
rect 21140 20896 21189 20924
rect 21140 20884 21146 20896
rect 21177 20893 21189 20896
rect 21223 20893 21235 20927
rect 21177 20887 21235 20893
rect 21361 20927 21419 20933
rect 21361 20893 21373 20927
rect 21407 20924 21419 20927
rect 21453 20927 21511 20933
rect 21453 20924 21465 20927
rect 21407 20896 21465 20924
rect 21407 20893 21419 20896
rect 21361 20887 21419 20893
rect 21453 20893 21465 20896
rect 21499 20893 21511 20927
rect 21453 20887 21511 20893
rect 21637 20927 21695 20933
rect 21637 20893 21649 20927
rect 21683 20893 21695 20927
rect 21637 20887 21695 20893
rect 22189 20927 22247 20933
rect 22189 20893 22201 20927
rect 22235 20924 22247 20927
rect 22664 20924 22692 21088
rect 23032 21032 23520 21060
rect 22235 20896 22692 20924
rect 22235 20893 22247 20896
rect 22189 20887 22247 20893
rect 21376 20856 21404 20887
rect 21100 20828 21404 20856
rect 21652 20856 21680 20887
rect 22830 20884 22836 20936
rect 22888 20884 22894 20936
rect 23032 20924 23060 21032
rect 23109 20927 23167 20933
rect 23109 20924 23121 20927
rect 23032 20896 23121 20924
rect 23109 20893 23121 20896
rect 23155 20893 23167 20927
rect 23109 20887 23167 20893
rect 23201 20927 23259 20933
rect 23201 20893 23213 20927
rect 23247 20924 23259 20927
rect 23382 20924 23388 20936
rect 23247 20896 23388 20924
rect 23247 20893 23259 20896
rect 23201 20887 23259 20893
rect 22002 20856 22008 20868
rect 21652 20828 22008 20856
rect 20180 20760 20760 20788
rect 19981 20751 20039 20757
rect 20990 20748 20996 20800
rect 21048 20788 21054 20800
rect 21100 20797 21128 20828
rect 22002 20816 22008 20828
rect 22060 20816 22066 20868
rect 22281 20859 22339 20865
rect 22281 20825 22293 20859
rect 22327 20856 22339 20859
rect 23017 20859 23075 20865
rect 22327 20828 22508 20856
rect 22327 20825 22339 20828
rect 22281 20819 22339 20825
rect 21085 20791 21143 20797
rect 21085 20788 21097 20791
rect 21048 20760 21097 20788
rect 21048 20748 21054 20760
rect 21085 20757 21097 20760
rect 21131 20757 21143 20791
rect 21085 20751 21143 20757
rect 22370 20748 22376 20800
rect 22428 20748 22434 20800
rect 22480 20788 22508 20828
rect 23017 20825 23029 20859
rect 23063 20856 23075 20859
rect 23216 20856 23244 20887
rect 23382 20884 23388 20896
rect 23440 20884 23446 20936
rect 23492 20933 23520 21032
rect 23477 20927 23535 20933
rect 23477 20893 23489 20927
rect 23523 20924 23535 20927
rect 25314 20924 25320 20936
rect 23523 20896 25320 20924
rect 23523 20893 23535 20896
rect 23477 20887 23535 20893
rect 25314 20884 25320 20896
rect 25372 20884 25378 20936
rect 23063 20828 23244 20856
rect 23063 20825 23075 20828
rect 23017 20819 23075 20825
rect 23290 20816 23296 20868
rect 23348 20816 23354 20868
rect 22738 20788 22744 20800
rect 22480 20760 22744 20788
rect 22738 20748 22744 20760
rect 22796 20788 22802 20800
rect 23201 20791 23259 20797
rect 23201 20788 23213 20791
rect 22796 20760 23213 20788
rect 22796 20748 22802 20760
rect 23201 20757 23213 20760
rect 23247 20757 23259 20791
rect 23201 20751 23259 20757
rect 1104 20698 27876 20720
rect 1104 20646 4874 20698
rect 4926 20646 4938 20698
rect 4990 20646 5002 20698
rect 5054 20646 5066 20698
rect 5118 20646 5130 20698
rect 5182 20646 27876 20698
rect 1104 20624 27876 20646
rect 5261 20587 5319 20593
rect 5261 20553 5273 20587
rect 5307 20584 5319 20587
rect 5350 20584 5356 20596
rect 5307 20556 5356 20584
rect 5307 20553 5319 20556
rect 5261 20547 5319 20553
rect 5350 20544 5356 20556
rect 5408 20544 5414 20596
rect 5994 20544 6000 20596
rect 6052 20584 6058 20596
rect 7006 20584 7012 20596
rect 6052 20556 7012 20584
rect 6052 20544 6058 20556
rect 7006 20544 7012 20556
rect 7064 20544 7070 20596
rect 9309 20587 9367 20593
rect 9309 20553 9321 20587
rect 9355 20584 9367 20587
rect 9674 20584 9680 20596
rect 9355 20556 9680 20584
rect 9355 20553 9367 20556
rect 9309 20547 9367 20553
rect 9674 20544 9680 20556
rect 9732 20544 9738 20596
rect 12802 20544 12808 20596
rect 12860 20584 12866 20596
rect 12897 20587 12955 20593
rect 12897 20584 12909 20587
rect 12860 20556 12909 20584
rect 12860 20544 12866 20556
rect 12897 20553 12909 20556
rect 12943 20584 12955 20587
rect 13354 20584 13360 20596
rect 12943 20556 13360 20584
rect 12943 20553 12955 20556
rect 12897 20547 12955 20553
rect 13354 20544 13360 20556
rect 13412 20544 13418 20596
rect 20254 20544 20260 20596
rect 20312 20584 20318 20596
rect 20349 20587 20407 20593
rect 20349 20584 20361 20587
rect 20312 20556 20361 20584
rect 20312 20544 20318 20556
rect 20349 20553 20361 20556
rect 20395 20553 20407 20587
rect 20349 20547 20407 20553
rect 5629 20519 5687 20525
rect 5629 20485 5641 20519
rect 5675 20516 5687 20519
rect 5718 20516 5724 20528
rect 5675 20488 5724 20516
rect 5675 20485 5687 20488
rect 5629 20479 5687 20485
rect 5718 20476 5724 20488
rect 5776 20476 5782 20528
rect 6822 20476 6828 20528
rect 6880 20516 6886 20528
rect 6917 20519 6975 20525
rect 6917 20516 6929 20519
rect 6880 20488 6929 20516
rect 6880 20476 6886 20488
rect 6917 20485 6929 20488
rect 6963 20516 6975 20519
rect 8018 20516 8024 20528
rect 6963 20488 8024 20516
rect 6963 20485 6975 20488
rect 6917 20479 6975 20485
rect 8018 20476 8024 20488
rect 8076 20476 8082 20528
rect 10778 20476 10784 20528
rect 10836 20476 10842 20528
rect 16942 20516 16948 20528
rect 11532 20488 12020 20516
rect 3878 20408 3884 20460
rect 3936 20448 3942 20460
rect 4617 20451 4675 20457
rect 4617 20448 4629 20451
rect 3936 20420 4629 20448
rect 3936 20408 3942 20420
rect 4617 20417 4629 20420
rect 4663 20417 4675 20451
rect 4617 20411 4675 20417
rect 5169 20451 5227 20457
rect 5169 20417 5181 20451
rect 5215 20448 5227 20451
rect 5258 20448 5264 20460
rect 5215 20420 5264 20448
rect 5215 20417 5227 20420
rect 5169 20411 5227 20417
rect 5258 20408 5264 20420
rect 5316 20408 5322 20460
rect 5813 20451 5871 20457
rect 5813 20417 5825 20451
rect 5859 20448 5871 20451
rect 6546 20448 6552 20460
rect 5859 20420 6552 20448
rect 5859 20417 5871 20420
rect 5813 20411 5871 20417
rect 6546 20408 6552 20420
rect 6604 20408 6610 20460
rect 8941 20451 8999 20457
rect 8941 20417 8953 20451
rect 8987 20448 8999 20451
rect 9953 20451 10011 20457
rect 9953 20448 9965 20451
rect 8987 20420 9965 20448
rect 8987 20417 8999 20420
rect 8941 20411 8999 20417
rect 9953 20417 9965 20420
rect 9999 20417 10011 20451
rect 9953 20411 10011 20417
rect 10594 20408 10600 20460
rect 10652 20408 10658 20460
rect 10689 20451 10747 20457
rect 10689 20417 10701 20451
rect 10735 20417 10747 20451
rect 10689 20411 10747 20417
rect 10965 20451 11023 20457
rect 10965 20417 10977 20451
rect 11011 20448 11023 20451
rect 11422 20448 11428 20460
rect 11011 20420 11428 20448
rect 11011 20417 11023 20420
rect 10965 20411 11023 20417
rect 3234 20340 3240 20392
rect 3292 20340 3298 20392
rect 4525 20383 4583 20389
rect 4525 20349 4537 20383
rect 4571 20380 4583 20383
rect 6362 20380 6368 20392
rect 4571 20352 6368 20380
rect 4571 20349 4583 20352
rect 4525 20343 4583 20349
rect 6362 20340 6368 20352
rect 6420 20340 6426 20392
rect 9030 20340 9036 20392
rect 9088 20340 9094 20392
rect 10318 20340 10324 20392
rect 10376 20380 10382 20392
rect 10704 20380 10732 20411
rect 11422 20408 11428 20420
rect 11480 20408 11486 20460
rect 11532 20457 11560 20488
rect 11517 20451 11575 20457
rect 11517 20417 11529 20451
rect 11563 20417 11575 20451
rect 11773 20451 11831 20457
rect 11773 20448 11785 20451
rect 11517 20411 11575 20417
rect 11624 20420 11785 20448
rect 11624 20380 11652 20420
rect 11773 20417 11785 20420
rect 11819 20417 11831 20451
rect 11992 20448 12020 20488
rect 13924 20488 16948 20516
rect 12618 20448 12624 20460
rect 11992 20420 12624 20448
rect 11773 20411 11831 20417
rect 12618 20408 12624 20420
rect 12676 20408 12682 20460
rect 13722 20448 13728 20460
rect 13372 20420 13728 20448
rect 10376 20352 10732 20380
rect 10980 20352 11652 20380
rect 10376 20340 10382 20352
rect 6641 20315 6699 20321
rect 6641 20281 6653 20315
rect 6687 20312 6699 20315
rect 7190 20312 7196 20324
rect 6687 20284 7196 20312
rect 6687 20281 6699 20284
rect 6641 20275 6699 20281
rect 7190 20272 7196 20284
rect 7248 20312 7254 20324
rect 8110 20312 8116 20324
rect 7248 20284 8116 20312
rect 7248 20272 7254 20284
rect 8110 20272 8116 20284
rect 8168 20272 8174 20324
rect 10980 20321 11008 20352
rect 10965 20315 11023 20321
rect 10965 20281 10977 20315
rect 11011 20281 11023 20315
rect 10965 20275 11023 20281
rect 2682 20204 2688 20256
rect 2740 20204 2746 20256
rect 3881 20247 3939 20253
rect 3881 20213 3893 20247
rect 3927 20244 3939 20247
rect 4062 20244 4068 20256
rect 3927 20216 4068 20244
rect 3927 20213 3939 20216
rect 3881 20207 3939 20213
rect 4062 20204 4068 20216
rect 4120 20204 4126 20256
rect 5445 20247 5503 20253
rect 5445 20213 5457 20247
rect 5491 20244 5503 20247
rect 5626 20244 5632 20256
rect 5491 20216 5632 20244
rect 5491 20213 5503 20216
rect 5445 20207 5503 20213
rect 5626 20204 5632 20216
rect 5684 20204 5690 20256
rect 6457 20247 6515 20253
rect 6457 20213 6469 20247
rect 6503 20244 6515 20247
rect 6822 20244 6828 20256
rect 6503 20216 6828 20244
rect 6503 20213 6515 20216
rect 6457 20207 6515 20213
rect 6822 20204 6828 20216
rect 6880 20204 6886 20256
rect 10778 20204 10784 20256
rect 10836 20244 10842 20256
rect 13372 20244 13400 20420
rect 13722 20408 13728 20420
rect 13780 20408 13786 20460
rect 13924 20457 13952 20488
rect 16942 20476 16948 20488
rect 17000 20516 17006 20528
rect 18782 20516 18788 20528
rect 17000 20488 18788 20516
rect 17000 20476 17006 20488
rect 18782 20476 18788 20488
rect 18840 20476 18846 20528
rect 20438 20476 20444 20528
rect 20496 20516 20502 20528
rect 20533 20519 20591 20525
rect 20533 20516 20545 20519
rect 20496 20488 20545 20516
rect 20496 20476 20502 20488
rect 20533 20485 20545 20488
rect 20579 20485 20591 20519
rect 20533 20479 20591 20485
rect 13814 20451 13872 20457
rect 13814 20417 13826 20451
rect 13860 20417 13872 20451
rect 13814 20411 13872 20417
rect 13909 20451 13967 20457
rect 13909 20417 13921 20451
rect 13955 20417 13967 20451
rect 13909 20411 13967 20417
rect 14093 20451 14151 20457
rect 14093 20417 14105 20451
rect 14139 20448 14151 20451
rect 14182 20448 14188 20460
rect 14139 20420 14188 20448
rect 14139 20417 14151 20420
rect 14093 20411 14151 20417
rect 13816 20312 13844 20411
rect 14182 20408 14188 20420
rect 14240 20408 14246 20460
rect 14550 20408 14556 20460
rect 14608 20408 14614 20460
rect 15378 20408 15384 20460
rect 15436 20448 15442 20460
rect 16025 20451 16083 20457
rect 16025 20448 16037 20451
rect 15436 20420 16037 20448
rect 15436 20408 15442 20420
rect 16025 20417 16037 20420
rect 16071 20448 16083 20451
rect 17678 20448 17684 20460
rect 16071 20420 17684 20448
rect 16071 20417 16083 20420
rect 16025 20411 16083 20417
rect 17678 20408 17684 20420
rect 17736 20408 17742 20460
rect 19886 20408 19892 20460
rect 19944 20448 19950 20460
rect 20257 20451 20315 20457
rect 20257 20448 20269 20451
rect 19944 20420 20269 20448
rect 19944 20408 19950 20420
rect 20257 20417 20269 20420
rect 20303 20417 20315 20451
rect 20257 20411 20315 20417
rect 14568 20380 14596 20408
rect 15838 20380 15844 20392
rect 14568 20352 15844 20380
rect 15838 20340 15844 20352
rect 15896 20340 15902 20392
rect 24210 20340 24216 20392
rect 24268 20380 24274 20392
rect 24305 20383 24363 20389
rect 24305 20380 24317 20383
rect 24268 20352 24317 20380
rect 24268 20340 24274 20352
rect 24305 20349 24317 20352
rect 24351 20349 24363 20383
rect 24305 20343 24363 20349
rect 15286 20312 15292 20324
rect 13816 20284 15292 20312
rect 15286 20272 15292 20284
rect 15344 20272 15350 20324
rect 20530 20272 20536 20324
rect 20588 20272 20594 20324
rect 24029 20315 24087 20321
rect 24029 20281 24041 20315
rect 24075 20312 24087 20315
rect 24394 20312 24400 20324
rect 24075 20284 24400 20312
rect 24075 20281 24087 20284
rect 24029 20275 24087 20281
rect 24394 20272 24400 20284
rect 24452 20272 24458 20324
rect 10836 20216 13400 20244
rect 10836 20204 10842 20216
rect 13446 20204 13452 20256
rect 13504 20204 13510 20256
rect 14182 20204 14188 20256
rect 14240 20244 14246 20256
rect 14369 20247 14427 20253
rect 14369 20244 14381 20247
rect 14240 20216 14381 20244
rect 14240 20204 14246 20216
rect 14369 20213 14381 20216
rect 14415 20213 14427 20247
rect 14369 20207 14427 20213
rect 15746 20204 15752 20256
rect 15804 20204 15810 20256
rect 21634 20204 21640 20256
rect 21692 20244 21698 20256
rect 23845 20247 23903 20253
rect 23845 20244 23857 20247
rect 21692 20216 23857 20244
rect 21692 20204 21698 20216
rect 23845 20213 23857 20216
rect 23891 20213 23903 20247
rect 23845 20207 23903 20213
rect 1104 20154 27876 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 27876 20154
rect 1104 20080 27876 20102
rect 1302 20000 1308 20052
rect 1360 20040 1366 20052
rect 1360 20012 10640 20040
rect 1360 20000 1366 20012
rect 3605 19975 3663 19981
rect 3605 19941 3617 19975
rect 3651 19972 3663 19975
rect 6362 19972 6368 19984
rect 3651 19944 6368 19972
rect 3651 19941 3663 19944
rect 3605 19935 3663 19941
rect 6362 19932 6368 19944
rect 6420 19932 6426 19984
rect 6546 19932 6552 19984
rect 6604 19932 6610 19984
rect 8018 19932 8024 19984
rect 8076 19972 8082 19984
rect 8389 19975 8447 19981
rect 8389 19972 8401 19975
rect 8076 19944 8401 19972
rect 8076 19932 8082 19944
rect 8389 19941 8401 19944
rect 8435 19941 8447 19975
rect 8389 19935 8447 19941
rect 9033 19975 9091 19981
rect 9033 19941 9045 19975
rect 9079 19972 9091 19975
rect 9306 19972 9312 19984
rect 9079 19944 9312 19972
rect 9079 19941 9091 19944
rect 9033 19935 9091 19941
rect 9306 19932 9312 19944
rect 9364 19932 9370 19984
rect 6178 19864 6184 19916
rect 6236 19904 6242 19916
rect 6564 19904 6592 19932
rect 6236 19876 6592 19904
rect 6236 19864 6242 19876
rect 8110 19864 8116 19916
rect 8168 19864 8174 19916
rect 9140 19876 9996 19904
rect 842 19796 848 19848
rect 900 19836 906 19848
rect 1397 19839 1455 19845
rect 1397 19836 1409 19839
rect 900 19808 1409 19836
rect 900 19796 906 19808
rect 1397 19805 1409 19808
rect 1443 19805 1455 19839
rect 1397 19799 1455 19805
rect 2225 19839 2283 19845
rect 2225 19805 2237 19839
rect 2271 19836 2283 19839
rect 2774 19836 2780 19848
rect 2271 19808 2780 19836
rect 2271 19805 2283 19808
rect 2225 19799 2283 19805
rect 2774 19796 2780 19808
rect 2832 19796 2838 19848
rect 6641 19839 6699 19845
rect 6641 19836 6653 19839
rect 4264 19808 6653 19836
rect 2492 19771 2550 19777
rect 2492 19737 2504 19771
rect 2538 19768 2550 19771
rect 2682 19768 2688 19780
rect 2538 19740 2688 19768
rect 2538 19737 2550 19740
rect 2492 19731 2550 19737
rect 2682 19728 2688 19740
rect 2740 19728 2746 19780
rect 3878 19728 3884 19780
rect 3936 19768 3942 19780
rect 4264 19777 4292 19808
rect 6641 19805 6653 19808
rect 6687 19805 6699 19839
rect 8202 19836 8208 19848
rect 6641 19799 6699 19805
rect 7576 19808 8208 19836
rect 7576 19780 7604 19808
rect 8202 19796 8208 19808
rect 8260 19836 8266 19848
rect 9140 19836 9168 19876
rect 8260 19808 9168 19836
rect 9217 19839 9275 19845
rect 8260 19796 8266 19808
rect 9217 19805 9229 19839
rect 9263 19836 9275 19839
rect 9766 19836 9772 19848
rect 9263 19808 9772 19836
rect 9263 19805 9275 19808
rect 9217 19799 9275 19805
rect 9766 19796 9772 19808
rect 9824 19796 9830 19848
rect 9968 19845 9996 19876
rect 9953 19839 10011 19845
rect 9953 19805 9965 19839
rect 9999 19805 10011 19839
rect 9953 19799 10011 19805
rect 10137 19839 10195 19845
rect 10137 19805 10149 19839
rect 10183 19836 10195 19839
rect 10318 19836 10324 19848
rect 10183 19808 10324 19836
rect 10183 19805 10195 19808
rect 10137 19799 10195 19805
rect 10318 19796 10324 19808
rect 10376 19796 10382 19848
rect 10612 19845 10640 20012
rect 11882 20000 11888 20052
rect 11940 20040 11946 20052
rect 15010 20040 15016 20052
rect 11940 20012 15016 20040
rect 11940 20000 11946 20012
rect 15010 20000 15016 20012
rect 15068 20000 15074 20052
rect 15197 20043 15255 20049
rect 15197 20009 15209 20043
rect 15243 20009 15255 20043
rect 15197 20003 15255 20009
rect 14642 19932 14648 19984
rect 14700 19972 14706 19984
rect 15212 19972 15240 20003
rect 15286 20000 15292 20052
rect 15344 20040 15350 20052
rect 15657 20043 15715 20049
rect 15657 20040 15669 20043
rect 15344 20012 15669 20040
rect 15344 20000 15350 20012
rect 15657 20009 15669 20012
rect 15703 20040 15715 20043
rect 15746 20040 15752 20052
rect 15703 20012 15752 20040
rect 15703 20009 15715 20012
rect 15657 20003 15715 20009
rect 15746 20000 15752 20012
rect 15804 20000 15810 20052
rect 16114 20000 16120 20052
rect 16172 20040 16178 20052
rect 16172 20012 16252 20040
rect 16172 20000 16178 20012
rect 14700 19944 15240 19972
rect 14700 19932 14706 19944
rect 15470 19904 15476 19916
rect 13556 19876 15476 19904
rect 10597 19839 10655 19845
rect 10597 19805 10609 19839
rect 10643 19805 10655 19839
rect 10597 19799 10655 19805
rect 12529 19839 12587 19845
rect 12529 19805 12541 19839
rect 12575 19836 12587 19839
rect 12618 19836 12624 19848
rect 12575 19808 12624 19836
rect 12575 19805 12587 19808
rect 12529 19799 12587 19805
rect 12618 19796 12624 19808
rect 12676 19796 12682 19848
rect 13078 19796 13084 19848
rect 13136 19836 13142 19848
rect 13556 19836 13584 19876
rect 15470 19864 15476 19876
rect 15528 19864 15534 19916
rect 15654 19864 15660 19916
rect 15712 19864 15718 19916
rect 16224 19913 16252 20012
rect 17678 20000 17684 20052
rect 17736 20000 17742 20052
rect 18782 20000 18788 20052
rect 18840 20000 18846 20052
rect 20438 20000 20444 20052
rect 20496 20040 20502 20052
rect 20622 20040 20628 20052
rect 20496 20012 20628 20040
rect 20496 20000 20502 20012
rect 20622 20000 20628 20012
rect 20680 20040 20686 20052
rect 20717 20043 20775 20049
rect 20717 20040 20729 20043
rect 20680 20012 20729 20040
rect 20680 20000 20686 20012
rect 20717 20009 20729 20012
rect 20763 20009 20775 20043
rect 20717 20003 20775 20009
rect 16209 19907 16267 19913
rect 15856 19876 16160 19904
rect 13136 19808 13584 19836
rect 13136 19796 13142 19808
rect 14090 19796 14096 19848
rect 14148 19796 14154 19848
rect 15672 19836 15700 19864
rect 15304 19808 15700 19836
rect 4249 19771 4307 19777
rect 4249 19768 4261 19771
rect 3936 19740 4261 19768
rect 3936 19728 3942 19740
rect 4249 19737 4261 19740
rect 4295 19737 4307 19771
rect 4249 19731 4307 19737
rect 5994 19728 6000 19780
rect 6052 19728 6058 19780
rect 6086 19728 6092 19780
rect 6144 19728 6150 19780
rect 6908 19771 6966 19777
rect 6908 19737 6920 19771
rect 6954 19768 6966 19771
rect 7006 19768 7012 19780
rect 6954 19740 7012 19768
rect 6954 19737 6966 19740
rect 6908 19731 6966 19737
rect 7006 19728 7012 19740
rect 7064 19728 7070 19780
rect 7558 19728 7564 19780
rect 7616 19728 7622 19780
rect 12796 19771 12854 19777
rect 8588 19740 10180 19768
rect 1581 19703 1639 19709
rect 1581 19669 1593 19703
rect 1627 19700 1639 19703
rect 1670 19700 1676 19712
rect 1627 19672 1676 19700
rect 1627 19669 1639 19672
rect 1581 19663 1639 19669
rect 1670 19660 1676 19672
rect 1728 19660 1734 19712
rect 5902 19660 5908 19712
rect 5960 19700 5966 19712
rect 6454 19700 6460 19712
rect 5960 19672 6460 19700
rect 5960 19660 5966 19672
rect 6454 19660 6460 19672
rect 6512 19700 6518 19712
rect 8588 19709 8616 19740
rect 10152 19712 10180 19740
rect 12796 19737 12808 19771
rect 12842 19768 12854 19771
rect 13814 19768 13820 19780
rect 12842 19740 13820 19768
rect 12842 19737 12854 19740
rect 12796 19731 12854 19737
rect 13814 19728 13820 19740
rect 13872 19728 13878 19780
rect 14550 19768 14556 19780
rect 13924 19740 14556 19768
rect 8573 19703 8631 19709
rect 8573 19700 8585 19703
rect 6512 19672 8585 19700
rect 6512 19660 6518 19672
rect 8573 19669 8585 19672
rect 8619 19669 8631 19703
rect 8573 19663 8631 19669
rect 9674 19660 9680 19712
rect 9732 19700 9738 19712
rect 10045 19703 10103 19709
rect 10045 19700 10057 19703
rect 9732 19672 10057 19700
rect 9732 19660 9738 19672
rect 10045 19669 10057 19672
rect 10091 19669 10103 19703
rect 10045 19663 10103 19669
rect 10134 19660 10140 19712
rect 10192 19660 10198 19712
rect 13924 19709 13952 19740
rect 14550 19728 14556 19740
rect 14608 19728 14614 19780
rect 15181 19771 15239 19777
rect 15181 19737 15193 19771
rect 15227 19768 15239 19771
rect 15304 19768 15332 19808
rect 15227 19740 15332 19768
rect 15227 19737 15239 19740
rect 15181 19731 15239 19737
rect 15378 19728 15384 19780
rect 15436 19728 15442 19780
rect 15562 19728 15568 19780
rect 15620 19777 15626 19780
rect 15856 19777 15884 19876
rect 15930 19796 15936 19848
rect 15988 19796 15994 19848
rect 16025 19839 16083 19845
rect 16025 19805 16037 19839
rect 16071 19805 16083 19839
rect 16025 19799 16083 19805
rect 15620 19771 15683 19777
rect 15620 19737 15637 19771
rect 15671 19737 15683 19771
rect 15620 19731 15683 19737
rect 15841 19771 15899 19777
rect 15841 19737 15853 19771
rect 15887 19737 15899 19771
rect 16040 19768 16068 19799
rect 15841 19731 15899 19737
rect 15948 19740 16068 19768
rect 16132 19768 16160 19876
rect 16209 19873 16221 19907
rect 16255 19904 16267 19907
rect 17696 19904 17724 20000
rect 18325 19907 18383 19913
rect 18325 19904 18337 19907
rect 16255 19876 16436 19904
rect 17696 19876 18337 19904
rect 16255 19873 16267 19876
rect 16209 19867 16267 19873
rect 16298 19796 16304 19848
rect 16356 19796 16362 19848
rect 16408 19836 16436 19876
rect 18325 19873 18337 19876
rect 18371 19873 18383 19907
rect 18325 19867 18383 19873
rect 18690 19864 18696 19916
rect 18748 19904 18754 19916
rect 19245 19907 19303 19913
rect 19245 19904 19257 19907
rect 18748 19876 19257 19904
rect 18748 19864 18754 19876
rect 19245 19873 19257 19876
rect 19291 19873 19303 19907
rect 19245 19867 19303 19873
rect 19705 19907 19763 19913
rect 19705 19873 19717 19907
rect 19751 19904 19763 19907
rect 19981 19907 20039 19913
rect 19981 19904 19993 19907
rect 19751 19876 19993 19904
rect 19751 19873 19763 19876
rect 19705 19867 19763 19873
rect 19981 19873 19993 19876
rect 20027 19873 20039 19907
rect 20732 19904 20760 20003
rect 22462 20000 22468 20052
rect 22520 20040 22526 20052
rect 22649 20043 22707 20049
rect 22649 20040 22661 20043
rect 22520 20012 22661 20040
rect 22520 20000 22526 20012
rect 22649 20009 22661 20012
rect 22695 20009 22707 20043
rect 22649 20003 22707 20009
rect 24026 20000 24032 20052
rect 24084 20000 24090 20052
rect 24210 20000 24216 20052
rect 24268 20040 24274 20052
rect 24489 20043 24547 20049
rect 24489 20040 24501 20043
rect 24268 20012 24501 20040
rect 24268 20000 24274 20012
rect 24489 20009 24501 20012
rect 24535 20009 24547 20043
rect 24489 20003 24547 20009
rect 20901 19975 20959 19981
rect 20901 19941 20913 19975
rect 20947 19972 20959 19975
rect 24949 19975 25007 19981
rect 24949 19972 24961 19975
rect 20947 19944 24961 19972
rect 20947 19941 20959 19944
rect 20901 19935 20959 19941
rect 24949 19941 24961 19944
rect 24995 19941 25007 19975
rect 24949 19935 25007 19941
rect 21269 19907 21327 19913
rect 21269 19904 21281 19907
rect 19981 19867 20039 19873
rect 20180 19876 20576 19904
rect 20732 19876 21281 19904
rect 17034 19836 17040 19848
rect 16408 19808 17040 19836
rect 17034 19796 17040 19808
rect 17092 19796 17098 19848
rect 18509 19839 18567 19845
rect 18509 19805 18521 19839
rect 18555 19836 18567 19839
rect 18598 19836 18604 19848
rect 18555 19808 18604 19836
rect 18555 19805 18567 19808
rect 18509 19799 18567 19805
rect 18598 19796 18604 19808
rect 18656 19836 18662 19848
rect 18656 19808 19564 19836
rect 18656 19796 18662 19808
rect 16390 19768 16396 19780
rect 16132 19740 16396 19768
rect 15620 19728 15626 19731
rect 13909 19703 13967 19709
rect 13909 19669 13921 19703
rect 13955 19669 13967 19703
rect 13909 19663 13967 19669
rect 14274 19660 14280 19712
rect 14332 19660 14338 19712
rect 14642 19660 14648 19712
rect 14700 19660 14706 19712
rect 14918 19660 14924 19712
rect 14976 19700 14982 19712
rect 15013 19703 15071 19709
rect 15013 19700 15025 19703
rect 14976 19672 15025 19700
rect 14976 19660 14982 19672
rect 15013 19669 15025 19672
rect 15059 19669 15071 19703
rect 15013 19663 15071 19669
rect 15470 19660 15476 19712
rect 15528 19700 15534 19712
rect 15948 19700 15976 19740
rect 16390 19728 16396 19740
rect 16448 19728 16454 19780
rect 16568 19771 16626 19777
rect 16568 19737 16580 19771
rect 16614 19768 16626 19771
rect 16666 19768 16672 19780
rect 16614 19740 16672 19768
rect 16614 19737 16626 19740
rect 16568 19731 16626 19737
rect 16666 19728 16672 19740
rect 16724 19728 16730 19780
rect 18322 19728 18328 19780
rect 18380 19768 18386 19780
rect 18693 19771 18751 19777
rect 18693 19768 18705 19771
rect 18380 19740 18705 19768
rect 18380 19728 18386 19740
rect 18693 19737 18705 19740
rect 18739 19768 18751 19771
rect 18966 19768 18972 19780
rect 18739 19740 18972 19768
rect 18739 19737 18751 19740
rect 18693 19731 18751 19737
rect 18966 19728 18972 19740
rect 19024 19728 19030 19780
rect 19536 19768 19564 19808
rect 19610 19796 19616 19848
rect 19668 19796 19674 19848
rect 19886 19796 19892 19848
rect 19944 19796 19950 19848
rect 20070 19796 20076 19848
rect 20128 19796 20134 19848
rect 19904 19768 19932 19796
rect 19536 19740 19932 19768
rect 19978 19728 19984 19780
rect 20036 19768 20042 19780
rect 20180 19768 20208 19876
rect 20441 19839 20499 19845
rect 20441 19805 20453 19839
rect 20487 19805 20499 19839
rect 20548 19836 20576 19876
rect 21269 19873 21281 19876
rect 21315 19873 21327 19907
rect 21269 19867 21327 19873
rect 22189 19907 22247 19913
rect 22189 19873 22201 19907
rect 22235 19904 22247 19907
rect 22462 19904 22468 19916
rect 22235 19876 22468 19904
rect 22235 19873 22247 19876
rect 22189 19867 22247 19873
rect 22462 19864 22468 19876
rect 22520 19864 22526 19916
rect 22940 19876 23520 19904
rect 20809 19839 20867 19845
rect 20809 19836 20821 19839
rect 20548 19808 20821 19836
rect 20441 19799 20499 19805
rect 20809 19805 20821 19808
rect 20855 19836 20867 19839
rect 21726 19836 21732 19848
rect 20855 19808 21732 19836
rect 20855 19805 20867 19808
rect 20809 19799 20867 19805
rect 20036 19740 20208 19768
rect 20456 19768 20484 19799
rect 21726 19796 21732 19808
rect 21784 19796 21790 19848
rect 21910 19796 21916 19848
rect 21968 19796 21974 19848
rect 22940 19845 22968 19876
rect 23492 19848 23520 19876
rect 22557 19839 22615 19845
rect 22557 19836 22569 19839
rect 22296 19808 22569 19836
rect 20898 19768 20904 19780
rect 20456 19740 20904 19768
rect 20036 19728 20042 19740
rect 20898 19728 20904 19740
rect 20956 19728 20962 19780
rect 15528 19672 15976 19700
rect 16209 19703 16267 19709
rect 15528 19660 15534 19672
rect 16209 19669 16221 19703
rect 16255 19700 16267 19703
rect 16850 19700 16856 19712
rect 16255 19672 16856 19700
rect 16255 19669 16267 19672
rect 16209 19663 16267 19669
rect 16850 19660 16856 19672
rect 16908 19660 16914 19712
rect 17770 19660 17776 19712
rect 17828 19660 17834 19712
rect 20533 19703 20591 19709
rect 20533 19669 20545 19703
rect 20579 19700 20591 19703
rect 21082 19700 21088 19712
rect 20579 19672 21088 19700
rect 20579 19669 20591 19672
rect 20533 19663 20591 19669
rect 21082 19660 21088 19672
rect 21140 19660 21146 19712
rect 21177 19703 21235 19709
rect 21177 19669 21189 19703
rect 21223 19700 21235 19703
rect 21542 19700 21548 19712
rect 21223 19672 21548 19700
rect 21223 19669 21235 19672
rect 21177 19663 21235 19669
rect 21542 19660 21548 19672
rect 21600 19660 21606 19712
rect 22296 19700 22324 19808
rect 22557 19805 22569 19808
rect 22603 19805 22615 19839
rect 22557 19799 22615 19805
rect 22925 19839 22983 19845
rect 22925 19805 22937 19839
rect 22971 19805 22983 19839
rect 22925 19799 22983 19805
rect 23198 19796 23204 19848
rect 23256 19836 23262 19848
rect 23256 19808 23428 19836
rect 23256 19796 23262 19808
rect 22370 19728 22376 19780
rect 22428 19768 22434 19780
rect 23293 19771 23351 19777
rect 23293 19768 23305 19771
rect 22428 19740 23305 19768
rect 22428 19728 22434 19740
rect 23293 19737 23305 19740
rect 23339 19737 23351 19771
rect 23400 19768 23428 19808
rect 23474 19796 23480 19848
rect 23532 19796 23538 19848
rect 23753 19839 23811 19845
rect 23753 19805 23765 19839
rect 23799 19805 23811 19839
rect 23753 19799 23811 19805
rect 23768 19768 23796 19799
rect 24394 19796 24400 19848
rect 24452 19796 24458 19848
rect 24765 19839 24823 19845
rect 24765 19805 24777 19839
rect 24811 19836 24823 19839
rect 25222 19836 25228 19848
rect 24811 19808 25228 19836
rect 24811 19805 24823 19808
rect 24765 19799 24823 19805
rect 25222 19796 25228 19808
rect 25280 19796 25286 19848
rect 23400 19740 23796 19768
rect 23293 19731 23351 19737
rect 23768 19712 23796 19740
rect 23842 19728 23848 19780
rect 23900 19728 23906 19780
rect 23658 19700 23664 19712
rect 22296 19672 23664 19700
rect 23658 19660 23664 19672
rect 23716 19660 23722 19712
rect 23750 19660 23756 19712
rect 23808 19700 23814 19712
rect 24045 19703 24103 19709
rect 24045 19700 24057 19703
rect 23808 19672 24057 19700
rect 23808 19660 23814 19672
rect 24045 19669 24057 19672
rect 24091 19669 24103 19703
rect 24045 19663 24103 19669
rect 1104 19610 27876 19632
rect 1104 19558 4874 19610
rect 4926 19558 4938 19610
rect 4990 19558 5002 19610
rect 5054 19558 5066 19610
rect 5118 19558 5130 19610
rect 5182 19558 27876 19610
rect 1104 19536 27876 19558
rect 5169 19499 5227 19505
rect 5169 19465 5181 19499
rect 5215 19496 5227 19499
rect 6086 19496 6092 19508
rect 5215 19468 6092 19496
rect 5215 19465 5227 19468
rect 5169 19459 5227 19465
rect 6086 19456 6092 19468
rect 6144 19456 6150 19508
rect 6178 19456 6184 19508
rect 6236 19496 6242 19508
rect 6730 19496 6736 19508
rect 6236 19468 6736 19496
rect 6236 19456 6242 19468
rect 6730 19456 6736 19468
rect 6788 19456 6794 19508
rect 7006 19456 7012 19508
rect 7064 19456 7070 19508
rect 7650 19456 7656 19508
rect 7708 19496 7714 19508
rect 9306 19496 9312 19508
rect 7708 19468 9312 19496
rect 7708 19456 7714 19468
rect 2774 19428 2780 19440
rect 1412 19400 2780 19428
rect 1412 19369 1440 19400
rect 2774 19388 2780 19400
rect 2832 19428 2838 19440
rect 5813 19431 5871 19437
rect 2832 19400 3832 19428
rect 2832 19388 2838 19400
rect 1670 19369 1676 19372
rect 1397 19363 1455 19369
rect 1397 19329 1409 19363
rect 1443 19329 1455 19363
rect 1664 19360 1676 19369
rect 1631 19332 1676 19360
rect 1397 19323 1455 19329
rect 1664 19323 1676 19332
rect 1670 19320 1676 19323
rect 1728 19320 1734 19372
rect 3234 19360 3240 19372
rect 2792 19332 3240 19360
rect 2792 19233 2820 19332
rect 3234 19320 3240 19332
rect 3292 19320 3298 19372
rect 3804 19369 3832 19400
rect 5813 19397 5825 19431
rect 5859 19428 5871 19431
rect 5859 19400 6868 19428
rect 5859 19397 5871 19400
rect 5813 19391 5871 19397
rect 6840 19372 6868 19400
rect 6914 19388 6920 19440
rect 6972 19428 6978 19440
rect 7852 19437 7880 19468
rect 9306 19456 9312 19468
rect 9364 19456 9370 19508
rect 10778 19456 10784 19508
rect 10836 19456 10842 19508
rect 11422 19456 11428 19508
rect 11480 19496 11486 19508
rect 12253 19499 12311 19505
rect 12253 19496 12265 19499
rect 11480 19468 12265 19496
rect 11480 19456 11486 19468
rect 12253 19465 12265 19468
rect 12299 19465 12311 19499
rect 12253 19459 12311 19465
rect 13814 19456 13820 19508
rect 13872 19456 13878 19508
rect 13998 19496 14004 19508
rect 13924 19468 14004 19496
rect 7837 19431 7895 19437
rect 6972 19400 7052 19428
rect 6972 19388 6978 19400
rect 3789 19363 3847 19369
rect 3789 19329 3801 19363
rect 3835 19360 3847 19363
rect 3878 19360 3884 19372
rect 3835 19332 3884 19360
rect 3835 19329 3847 19332
rect 3789 19323 3847 19329
rect 3878 19320 3884 19332
rect 3936 19320 3942 19372
rect 4062 19369 4068 19372
rect 4056 19360 4068 19369
rect 4023 19332 4068 19360
rect 4056 19323 4068 19332
rect 4062 19320 4068 19323
rect 4120 19320 4126 19372
rect 5626 19320 5632 19372
rect 5684 19360 5690 19372
rect 5684 19332 5856 19360
rect 5684 19320 5690 19332
rect 5828 19292 5856 19332
rect 5902 19320 5908 19372
rect 5960 19320 5966 19372
rect 5997 19363 6055 19369
rect 5997 19329 6009 19363
rect 6043 19360 6055 19363
rect 6178 19360 6184 19372
rect 6043 19332 6184 19360
rect 6043 19329 6055 19332
rect 5997 19323 6055 19329
rect 6178 19320 6184 19332
rect 6236 19320 6242 19372
rect 6270 19320 6276 19372
rect 6328 19360 6334 19372
rect 6365 19363 6423 19369
rect 6365 19360 6377 19363
rect 6328 19332 6377 19360
rect 6328 19320 6334 19332
rect 6365 19329 6377 19332
rect 6411 19329 6423 19363
rect 6365 19323 6423 19329
rect 6454 19320 6460 19372
rect 6512 19360 6518 19372
rect 6641 19363 6699 19369
rect 6512 19332 6557 19360
rect 6512 19320 6518 19332
rect 6641 19329 6653 19363
rect 6687 19329 6699 19363
rect 6641 19323 6699 19329
rect 6656 19292 6684 19323
rect 6730 19320 6736 19372
rect 6788 19320 6794 19372
rect 6822 19320 6828 19372
rect 6880 19369 6886 19372
rect 6880 19360 6888 19369
rect 6880 19332 6925 19360
rect 6880 19323 6888 19332
rect 6880 19320 6886 19323
rect 7024 19292 7052 19400
rect 7837 19397 7849 19431
rect 7883 19397 7895 19431
rect 7837 19391 7895 19397
rect 8113 19431 8171 19437
rect 8113 19397 8125 19431
rect 8159 19428 8171 19431
rect 8450 19431 8508 19437
rect 8450 19428 8462 19431
rect 8159 19400 8462 19428
rect 8159 19397 8171 19400
rect 8113 19391 8171 19397
rect 8450 19397 8462 19400
rect 8496 19397 8508 19431
rect 8450 19391 8508 19397
rect 10226 19388 10232 19440
rect 10284 19388 10290 19440
rect 10318 19388 10324 19440
rect 10376 19428 10382 19440
rect 10965 19431 11023 19437
rect 10965 19428 10977 19431
rect 10376 19400 10977 19428
rect 10376 19388 10382 19400
rect 10965 19397 10977 19400
rect 11011 19397 11023 19431
rect 13924 19428 13952 19468
rect 13998 19456 14004 19468
rect 14056 19456 14062 19508
rect 15565 19499 15623 19505
rect 14108 19468 15516 19496
rect 14108 19437 14136 19468
rect 10965 19391 11023 19397
rect 11716 19400 12434 19428
rect 7558 19320 7564 19372
rect 7616 19369 7622 19372
rect 7616 19363 7665 19369
rect 7616 19329 7619 19363
rect 7653 19329 7665 19363
rect 7616 19323 7665 19329
rect 7616 19320 7622 19323
rect 7742 19320 7748 19372
rect 7800 19320 7806 19372
rect 7929 19363 7987 19369
rect 7929 19329 7941 19363
rect 7975 19360 7987 19363
rect 9766 19360 9772 19372
rect 7975 19332 9772 19360
rect 7975 19329 7987 19332
rect 7929 19323 7987 19329
rect 9766 19320 9772 19332
rect 9824 19320 9830 19372
rect 11716 19304 11744 19400
rect 11790 19320 11796 19372
rect 11848 19320 11854 19372
rect 12406 19360 12434 19400
rect 12912 19400 13952 19428
rect 14093 19431 14151 19437
rect 12912 19372 12940 19400
rect 14093 19397 14105 19431
rect 14139 19397 14151 19431
rect 14093 19391 14151 19397
rect 14274 19388 14280 19440
rect 14332 19437 14338 19440
rect 14332 19431 14361 19437
rect 14349 19397 14361 19431
rect 14332 19391 14361 19397
rect 14829 19431 14887 19437
rect 14829 19397 14841 19431
rect 14875 19397 14887 19431
rect 15289 19431 15347 19437
rect 15289 19428 15301 19431
rect 14829 19391 14887 19397
rect 15120 19400 15301 19428
rect 14332 19388 14338 19391
rect 12621 19363 12679 19369
rect 12621 19360 12633 19363
rect 12406 19332 12633 19360
rect 12621 19329 12633 19332
rect 12667 19360 12679 19363
rect 12802 19360 12808 19372
rect 12667 19332 12808 19360
rect 12667 19329 12679 19332
rect 12621 19323 12679 19329
rect 12802 19320 12808 19332
rect 12860 19320 12866 19372
rect 12894 19320 12900 19372
rect 12952 19320 12958 19372
rect 13078 19320 13084 19372
rect 13136 19320 13142 19372
rect 13170 19320 13176 19372
rect 13228 19320 13234 19372
rect 13265 19363 13323 19369
rect 13265 19329 13277 19363
rect 13311 19360 13323 19363
rect 13354 19360 13360 19372
rect 13311 19332 13360 19360
rect 13311 19329 13323 19332
rect 13265 19323 13323 19329
rect 13354 19320 13360 19332
rect 13412 19360 13418 19372
rect 13906 19360 13912 19372
rect 13412 19332 13912 19360
rect 13412 19320 13418 19332
rect 13906 19320 13912 19332
rect 13964 19320 13970 19372
rect 14001 19363 14059 19369
rect 14001 19329 14013 19363
rect 14047 19329 14059 19363
rect 14001 19323 14059 19329
rect 5828 19264 6684 19292
rect 6840 19264 7052 19292
rect 2777 19227 2835 19233
rect 2777 19193 2789 19227
rect 2823 19193 2835 19227
rect 2777 19187 2835 19193
rect 6181 19227 6239 19233
rect 6181 19193 6193 19227
rect 6227 19224 6239 19227
rect 6840 19224 6868 19264
rect 7098 19252 7104 19304
rect 7156 19292 7162 19304
rect 7469 19295 7527 19301
rect 7469 19292 7481 19295
rect 7156 19264 7481 19292
rect 7156 19252 7162 19264
rect 7469 19261 7481 19264
rect 7515 19261 7527 19295
rect 7469 19255 7527 19261
rect 8205 19295 8263 19301
rect 8205 19261 8217 19295
rect 8251 19261 8263 19295
rect 8205 19255 8263 19261
rect 6227 19196 6868 19224
rect 6227 19193 6239 19196
rect 6181 19187 6239 19193
rect 7006 19184 7012 19236
rect 7064 19224 7070 19236
rect 8220 19224 8248 19255
rect 10042 19252 10048 19304
rect 10100 19292 10106 19304
rect 11698 19301 11704 19304
rect 10689 19295 10747 19301
rect 10689 19292 10701 19295
rect 10100 19264 10701 19292
rect 10100 19252 10106 19264
rect 10689 19261 10701 19264
rect 10735 19261 10747 19295
rect 10689 19255 10747 19261
rect 11676 19295 11704 19301
rect 11676 19261 11688 19295
rect 11676 19255 11704 19261
rect 11698 19252 11704 19255
rect 11756 19252 11762 19304
rect 11885 19295 11943 19301
rect 11885 19261 11897 19295
rect 11931 19261 11943 19295
rect 11885 19255 11943 19261
rect 12161 19295 12219 19301
rect 12161 19261 12173 19295
rect 12207 19292 12219 19295
rect 12434 19292 12440 19304
rect 12207 19264 12440 19292
rect 12207 19261 12219 19264
rect 12161 19255 12219 19261
rect 7064 19196 8248 19224
rect 10229 19227 10287 19233
rect 7064 19184 7070 19196
rect 10229 19193 10241 19227
rect 10275 19224 10287 19227
rect 10410 19224 10416 19236
rect 10275 19196 10416 19224
rect 10275 19193 10287 19196
rect 10229 19187 10287 19193
rect 10410 19184 10416 19196
rect 10468 19184 10474 19236
rect 11238 19184 11244 19236
rect 11296 19224 11302 19236
rect 11900 19224 11928 19255
rect 12434 19252 12440 19264
rect 12492 19252 12498 19304
rect 12713 19295 12771 19301
rect 12713 19261 12725 19295
rect 12759 19292 12771 19295
rect 13446 19292 13452 19304
rect 12759 19264 13452 19292
rect 12759 19261 12771 19264
rect 12713 19255 12771 19261
rect 13446 19252 13452 19264
rect 13504 19252 13510 19304
rect 14016 19292 14044 19323
rect 14182 19320 14188 19372
rect 14240 19320 14246 19372
rect 14844 19360 14872 19391
rect 14384 19332 14872 19360
rect 14384 19292 14412 19332
rect 14918 19320 14924 19372
rect 14976 19360 14982 19372
rect 15120 19369 15148 19400
rect 15289 19397 15301 19400
rect 15335 19397 15347 19431
rect 15488 19428 15516 19468
rect 15565 19465 15577 19499
rect 15611 19496 15623 19499
rect 15930 19496 15936 19508
rect 15611 19468 15936 19496
rect 15611 19465 15623 19468
rect 15565 19459 15623 19465
rect 15930 19456 15936 19468
rect 15988 19456 15994 19508
rect 16666 19456 16672 19508
rect 16724 19456 16730 19508
rect 19518 19496 19524 19508
rect 16868 19468 19524 19496
rect 16868 19428 16896 19468
rect 19518 19456 19524 19468
rect 19576 19456 19582 19508
rect 19610 19456 19616 19508
rect 19668 19496 19674 19508
rect 19981 19499 20039 19505
rect 19981 19496 19993 19499
rect 19668 19468 19993 19496
rect 19668 19456 19674 19468
rect 19981 19465 19993 19468
rect 20027 19496 20039 19499
rect 20809 19499 20867 19505
rect 20027 19468 20760 19496
rect 20027 19465 20039 19468
rect 19981 19459 20039 19465
rect 15488 19400 16896 19428
rect 16945 19431 17003 19437
rect 15289 19391 15347 19397
rect 16945 19397 16957 19431
rect 16991 19428 17003 19431
rect 18601 19431 18659 19437
rect 18601 19428 18613 19431
rect 16991 19400 18613 19428
rect 16991 19397 17003 19400
rect 16945 19391 17003 19397
rect 18601 19397 18613 19400
rect 18647 19397 18659 19431
rect 18601 19391 18659 19397
rect 15013 19363 15071 19369
rect 15013 19360 15025 19363
rect 14976 19332 15025 19360
rect 14976 19320 14982 19332
rect 15013 19329 15025 19332
rect 15059 19329 15071 19363
rect 15013 19323 15071 19329
rect 15105 19363 15163 19369
rect 15105 19329 15117 19363
rect 15151 19329 15163 19363
rect 15105 19323 15163 19329
rect 15197 19363 15255 19369
rect 15197 19329 15209 19363
rect 15243 19329 15255 19363
rect 15197 19323 15255 19329
rect 14016 19264 14412 19292
rect 14461 19295 14519 19301
rect 14461 19261 14473 19295
rect 14507 19292 14519 19295
rect 14642 19292 14648 19304
rect 14507 19264 14648 19292
rect 14507 19261 14519 19264
rect 14461 19255 14519 19261
rect 11296 19196 11928 19224
rect 11296 19184 11302 19196
rect 12342 19184 12348 19236
rect 12400 19224 12406 19236
rect 14476 19224 14504 19255
rect 14642 19252 14648 19264
rect 14700 19252 14706 19304
rect 14734 19252 14740 19304
rect 14792 19292 14798 19304
rect 14829 19295 14887 19301
rect 14829 19292 14841 19295
rect 14792 19264 14841 19292
rect 14792 19252 14798 19264
rect 14829 19261 14841 19264
rect 14875 19261 14887 19295
rect 15212 19292 15240 19323
rect 15378 19320 15384 19372
rect 15436 19320 15442 19372
rect 15473 19363 15531 19369
rect 15473 19329 15485 19363
rect 15519 19329 15531 19363
rect 15473 19323 15531 19329
rect 14829 19255 14887 19261
rect 15120 19264 15240 19292
rect 15120 19224 15148 19264
rect 15286 19252 15292 19304
rect 15344 19292 15350 19304
rect 15488 19292 15516 19323
rect 15654 19320 15660 19372
rect 15712 19320 15718 19372
rect 15746 19320 15752 19372
rect 15804 19360 15810 19372
rect 16758 19360 16764 19372
rect 15804 19332 16764 19360
rect 15804 19320 15810 19332
rect 16758 19320 16764 19332
rect 16816 19320 16822 19372
rect 16850 19320 16856 19372
rect 16908 19320 16914 19372
rect 17034 19320 17040 19372
rect 17092 19320 17098 19372
rect 17155 19363 17213 19369
rect 17155 19360 17167 19363
rect 17144 19329 17167 19360
rect 17201 19329 17213 19363
rect 17144 19323 17213 19329
rect 17313 19363 17371 19369
rect 17313 19329 17325 19363
rect 17359 19360 17371 19363
rect 17770 19360 17776 19372
rect 17359 19332 17776 19360
rect 17359 19329 17371 19332
rect 17313 19323 17371 19329
rect 15344 19264 15516 19292
rect 16776 19292 16804 19320
rect 17144 19292 17172 19323
rect 17770 19320 17776 19332
rect 17828 19320 17834 19372
rect 18046 19320 18052 19372
rect 18104 19360 18110 19372
rect 18509 19363 18567 19369
rect 18509 19360 18521 19363
rect 18104 19332 18521 19360
rect 18104 19320 18110 19332
rect 18509 19329 18521 19332
rect 18555 19329 18567 19363
rect 18509 19323 18567 19329
rect 16776 19264 17172 19292
rect 15344 19252 15350 19264
rect 12400 19196 15148 19224
rect 12400 19184 12406 19196
rect 8938 19116 8944 19168
rect 8996 19156 9002 19168
rect 9490 19156 9496 19168
rect 8996 19128 9496 19156
rect 8996 19116 9002 19128
rect 9490 19116 9496 19128
rect 9548 19156 9554 19168
rect 9585 19159 9643 19165
rect 9585 19156 9597 19159
rect 9548 19128 9597 19156
rect 9548 19116 9554 19128
rect 9585 19125 9597 19128
rect 9631 19125 9643 19159
rect 9585 19119 9643 19125
rect 11146 19116 11152 19168
rect 11204 19156 11210 19168
rect 11517 19159 11575 19165
rect 11517 19156 11529 19159
rect 11204 19128 11529 19156
rect 11204 19116 11210 19128
rect 11517 19125 11529 19128
rect 11563 19125 11575 19159
rect 11517 19119 11575 19125
rect 13538 19116 13544 19168
rect 13596 19116 13602 19168
rect 14826 19116 14832 19168
rect 14884 19156 14890 19168
rect 15396 19156 15424 19264
rect 14884 19128 15424 19156
rect 18524 19156 18552 19323
rect 18690 19320 18696 19372
rect 18748 19320 18754 19372
rect 18966 19320 18972 19372
rect 19024 19320 19030 19372
rect 19797 19363 19855 19369
rect 19797 19329 19809 19363
rect 19843 19360 19855 19363
rect 19978 19360 19984 19372
rect 19843 19332 19984 19360
rect 19843 19329 19855 19332
rect 19797 19323 19855 19329
rect 19978 19320 19984 19332
rect 20036 19320 20042 19372
rect 20070 19320 20076 19372
rect 20128 19320 20134 19372
rect 20180 19369 20208 19468
rect 20165 19363 20223 19369
rect 20165 19329 20177 19363
rect 20211 19329 20223 19363
rect 20165 19323 20223 19329
rect 20349 19363 20407 19369
rect 20349 19329 20361 19363
rect 20395 19360 20407 19363
rect 20441 19363 20499 19369
rect 20441 19360 20453 19363
rect 20395 19332 20453 19360
rect 20395 19329 20407 19332
rect 20349 19323 20407 19329
rect 20441 19329 20453 19332
rect 20487 19329 20499 19363
rect 20441 19323 20499 19329
rect 20088 19292 20116 19320
rect 20364 19292 20392 19323
rect 20622 19320 20628 19372
rect 20680 19320 20686 19372
rect 20088 19264 20392 19292
rect 20732 19292 20760 19468
rect 20809 19465 20821 19499
rect 20855 19496 20867 19499
rect 21082 19496 21088 19508
rect 20855 19468 21088 19496
rect 20855 19465 20867 19468
rect 20809 19459 20867 19465
rect 21082 19456 21088 19468
rect 21140 19456 21146 19508
rect 23842 19456 23848 19508
rect 23900 19496 23906 19508
rect 24397 19499 24455 19505
rect 24397 19496 24409 19499
rect 23900 19468 24409 19496
rect 23900 19456 23906 19468
rect 24397 19465 24409 19468
rect 24443 19465 24455 19499
rect 24397 19459 24455 19465
rect 22925 19431 22983 19437
rect 22925 19397 22937 19431
rect 22971 19397 22983 19431
rect 22925 19391 22983 19397
rect 23141 19431 23199 19437
rect 23141 19397 23153 19431
rect 23187 19428 23199 19431
rect 23382 19428 23388 19440
rect 23187 19400 23388 19428
rect 23187 19397 23199 19400
rect 23141 19391 23199 19397
rect 20898 19320 20904 19372
rect 20956 19320 20962 19372
rect 22940 19360 22968 19391
rect 23382 19388 23388 19400
rect 23440 19388 23446 19440
rect 23566 19388 23572 19440
rect 23624 19428 23630 19440
rect 23624 19400 24348 19428
rect 23624 19388 23630 19400
rect 23658 19360 23664 19372
rect 22940 19332 23664 19360
rect 23658 19320 23664 19332
rect 23716 19320 23722 19372
rect 23750 19320 23756 19372
rect 23808 19320 23814 19372
rect 24026 19320 24032 19372
rect 24084 19320 24090 19372
rect 24320 19369 24348 19400
rect 24305 19363 24363 19369
rect 24305 19329 24317 19363
rect 24351 19329 24363 19363
rect 24305 19323 24363 19329
rect 25041 19363 25099 19369
rect 25041 19329 25053 19363
rect 25087 19360 25099 19363
rect 25222 19360 25228 19372
rect 25087 19332 25228 19360
rect 25087 19329 25099 19332
rect 25041 19323 25099 19329
rect 25222 19320 25228 19332
rect 25280 19320 25286 19372
rect 21634 19292 21640 19304
rect 20732 19264 21640 19292
rect 21634 19252 21640 19264
rect 21692 19252 21698 19304
rect 24213 19295 24271 19301
rect 24213 19261 24225 19295
rect 24259 19292 24271 19295
rect 24394 19292 24400 19304
rect 24259 19264 24400 19292
rect 24259 19261 24271 19264
rect 24213 19255 24271 19261
rect 24394 19252 24400 19264
rect 24452 19252 24458 19304
rect 24946 19252 24952 19304
rect 25004 19252 25010 19304
rect 18690 19184 18696 19236
rect 18748 19224 18754 19236
rect 19613 19227 19671 19233
rect 19613 19224 19625 19227
rect 18748 19196 19625 19224
rect 18748 19184 18754 19196
rect 19613 19193 19625 19196
rect 19659 19193 19671 19227
rect 19613 19187 19671 19193
rect 21450 19184 21456 19236
rect 21508 19224 21514 19236
rect 24673 19227 24731 19233
rect 24673 19224 24685 19227
rect 21508 19196 24685 19224
rect 21508 19184 21514 19196
rect 24673 19193 24685 19196
rect 24719 19193 24731 19227
rect 24673 19187 24731 19193
rect 18874 19156 18880 19168
rect 18524 19128 18880 19156
rect 14884 19116 14890 19128
rect 18874 19116 18880 19128
rect 18932 19116 18938 19168
rect 20254 19116 20260 19168
rect 20312 19116 20318 19168
rect 21910 19116 21916 19168
rect 21968 19156 21974 19168
rect 23106 19156 23112 19168
rect 21968 19128 23112 19156
rect 21968 19116 21974 19128
rect 23106 19116 23112 19128
rect 23164 19116 23170 19168
rect 23293 19159 23351 19165
rect 23293 19125 23305 19159
rect 23339 19156 23351 19159
rect 23566 19156 23572 19168
rect 23339 19128 23572 19156
rect 23339 19125 23351 19128
rect 23293 19119 23351 19125
rect 23566 19116 23572 19128
rect 23624 19116 23630 19168
rect 1104 19066 27876 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 27876 19066
rect 1104 18992 27876 19014
rect 5258 18912 5264 18964
rect 5316 18952 5322 18964
rect 8662 18952 8668 18964
rect 5316 18924 8668 18952
rect 5316 18912 5322 18924
rect 8662 18912 8668 18924
rect 8720 18912 8726 18964
rect 9769 18955 9827 18961
rect 9769 18921 9781 18955
rect 9815 18952 9827 18955
rect 9858 18952 9864 18964
rect 9815 18924 9864 18952
rect 9815 18921 9827 18924
rect 9769 18915 9827 18921
rect 9858 18912 9864 18924
rect 9916 18912 9922 18964
rect 10410 18912 10416 18964
rect 10468 18912 10474 18964
rect 11238 18952 11244 18964
rect 10520 18924 11244 18952
rect 10134 18844 10140 18896
rect 10192 18884 10198 18896
rect 10520 18884 10548 18924
rect 11238 18912 11244 18924
rect 11296 18912 11302 18964
rect 12342 18912 12348 18964
rect 12400 18912 12406 18964
rect 13170 18912 13176 18964
rect 13228 18912 13234 18964
rect 14829 18955 14887 18961
rect 14829 18921 14841 18955
rect 14875 18921 14887 18955
rect 14829 18915 14887 18921
rect 10192 18856 10548 18884
rect 10192 18844 10198 18856
rect 10686 18844 10692 18896
rect 10744 18884 10750 18896
rect 10965 18887 11023 18893
rect 10965 18884 10977 18887
rect 10744 18856 10977 18884
rect 10744 18844 10750 18856
rect 10965 18853 10977 18856
rect 11011 18853 11023 18887
rect 11885 18887 11943 18893
rect 11885 18884 11897 18887
rect 10965 18847 11023 18853
rect 11532 18856 11897 18884
rect 3878 18776 3884 18828
rect 3936 18776 3942 18828
rect 10152 18816 10180 18844
rect 10229 18819 10287 18825
rect 10229 18816 10241 18819
rect 10152 18788 10241 18816
rect 10229 18785 10241 18788
rect 10275 18785 10287 18819
rect 11146 18816 11152 18828
rect 10229 18779 10287 18785
rect 10888 18788 11152 18816
rect 5445 18751 5503 18757
rect 5445 18717 5457 18751
rect 5491 18748 5503 18751
rect 5994 18748 6000 18760
rect 5491 18720 6000 18748
rect 5491 18717 5503 18720
rect 5445 18711 5503 18717
rect 5994 18708 6000 18720
rect 6052 18708 6058 18760
rect 9217 18751 9275 18757
rect 9217 18717 9229 18751
rect 9263 18748 9275 18751
rect 9674 18748 9680 18760
rect 9263 18720 9680 18748
rect 9263 18717 9275 18720
rect 9217 18711 9275 18717
rect 9674 18708 9680 18720
rect 9732 18708 9738 18760
rect 9950 18708 9956 18760
rect 10008 18708 10014 18760
rect 10042 18708 10048 18760
rect 10100 18708 10106 18760
rect 10137 18751 10195 18757
rect 10137 18717 10149 18751
rect 10183 18717 10195 18751
rect 10137 18711 10195 18717
rect 10594 18751 10652 18757
rect 10594 18717 10606 18751
rect 10640 18748 10652 18751
rect 10888 18748 10916 18788
rect 11146 18776 11152 18788
rect 11204 18776 11210 18828
rect 11532 18825 11560 18856
rect 11885 18853 11897 18856
rect 11931 18853 11943 18887
rect 14844 18884 14872 18915
rect 21634 18912 21640 18964
rect 21692 18912 21698 18964
rect 22830 18912 22836 18964
rect 22888 18952 22894 18964
rect 23017 18955 23075 18961
rect 23017 18952 23029 18955
rect 22888 18924 23029 18952
rect 22888 18912 22894 18924
rect 23017 18921 23029 18924
rect 23063 18921 23075 18955
rect 23017 18915 23075 18921
rect 23106 18912 23112 18964
rect 23164 18952 23170 18964
rect 23750 18952 23756 18964
rect 23164 18924 23756 18952
rect 23164 18912 23170 18924
rect 23750 18912 23756 18924
rect 23808 18912 23814 18964
rect 15286 18884 15292 18896
rect 11885 18847 11943 18853
rect 12176 18856 15292 18884
rect 11517 18819 11575 18825
rect 11517 18785 11529 18819
rect 11563 18785 11575 18819
rect 11517 18779 11575 18785
rect 12176 18760 12204 18856
rect 15286 18844 15292 18856
rect 15344 18844 15350 18896
rect 12989 18819 13047 18825
rect 12989 18785 13001 18819
rect 13035 18816 13047 18819
rect 13354 18816 13360 18828
rect 13035 18788 13360 18816
rect 13035 18785 13047 18788
rect 12989 18779 13047 18785
rect 13354 18776 13360 18788
rect 13412 18776 13418 18828
rect 14642 18776 14648 18828
rect 14700 18816 14706 18828
rect 16114 18816 16120 18828
rect 14700 18788 16120 18816
rect 14700 18776 14706 18788
rect 16114 18776 16120 18788
rect 16172 18776 16178 18828
rect 17972 18788 18460 18816
rect 10640 18720 10916 18748
rect 11057 18751 11115 18757
rect 10640 18717 10652 18720
rect 10594 18711 10652 18717
rect 11057 18717 11069 18751
rect 11103 18748 11115 18751
rect 11103 18720 11284 18748
rect 11103 18717 11115 18720
rect 11057 18711 11115 18717
rect 4148 18683 4206 18689
rect 4148 18649 4160 18683
rect 4194 18680 4206 18683
rect 4798 18680 4804 18692
rect 4194 18652 4804 18680
rect 4194 18649 4206 18652
rect 4148 18643 4206 18649
rect 4798 18640 4804 18652
rect 4856 18640 4862 18692
rect 8294 18640 8300 18692
rect 8352 18680 8358 18692
rect 10060 18680 10088 18708
rect 8352 18652 9076 18680
rect 8352 18640 8358 18652
rect 9048 18624 9076 18652
rect 9692 18652 10088 18680
rect 10152 18680 10180 18711
rect 10318 18680 10324 18692
rect 10152 18652 10324 18680
rect 9692 18624 9720 18652
rect 10318 18640 10324 18652
rect 10376 18680 10382 18692
rect 11149 18683 11207 18689
rect 11149 18680 11161 18683
rect 10376 18652 11161 18680
rect 10376 18640 10382 18652
rect 11149 18649 11161 18652
rect 11195 18649 11207 18683
rect 11149 18643 11207 18649
rect 5261 18615 5319 18621
rect 5261 18581 5273 18615
rect 5307 18612 5319 18615
rect 5718 18612 5724 18624
rect 5307 18584 5724 18612
rect 5307 18581 5319 18584
rect 5261 18575 5319 18581
rect 5718 18572 5724 18584
rect 5776 18572 5782 18624
rect 6638 18572 6644 18624
rect 6696 18612 6702 18624
rect 6733 18615 6791 18621
rect 6733 18612 6745 18615
rect 6696 18584 6745 18612
rect 6696 18572 6702 18584
rect 6733 18581 6745 18584
rect 6779 18612 6791 18615
rect 7006 18612 7012 18624
rect 6779 18584 7012 18612
rect 6779 18581 6791 18584
rect 6733 18575 6791 18581
rect 7006 18572 7012 18584
rect 7064 18572 7070 18624
rect 7098 18572 7104 18624
rect 7156 18612 7162 18624
rect 8938 18612 8944 18624
rect 7156 18584 8944 18612
rect 7156 18572 7162 18584
rect 8938 18572 8944 18584
rect 8996 18572 9002 18624
rect 9030 18572 9036 18624
rect 9088 18572 9094 18624
rect 9674 18572 9680 18624
rect 9732 18572 9738 18624
rect 10597 18615 10655 18621
rect 10597 18581 10609 18615
rect 10643 18612 10655 18615
rect 10962 18612 10968 18624
rect 10643 18584 10968 18612
rect 10643 18581 10655 18584
rect 10597 18575 10655 18581
rect 10962 18572 10968 18584
rect 11020 18572 11026 18624
rect 11256 18612 11284 18720
rect 11606 18708 11612 18760
rect 11664 18708 11670 18760
rect 11698 18708 11704 18760
rect 11756 18748 11762 18760
rect 12069 18751 12127 18757
rect 12069 18748 12081 18751
rect 11756 18720 12081 18748
rect 11756 18708 11762 18720
rect 12069 18717 12081 18720
rect 12115 18717 12127 18751
rect 12069 18711 12127 18717
rect 12158 18708 12164 18760
rect 12216 18708 12222 18760
rect 13262 18708 13268 18760
rect 13320 18708 13326 18760
rect 14734 18748 14740 18760
rect 14200 18720 14740 18748
rect 11974 18640 11980 18692
rect 12032 18680 12038 18692
rect 12434 18680 12440 18692
rect 12032 18652 12440 18680
rect 12032 18640 12038 18652
rect 12434 18640 12440 18652
rect 12492 18680 12498 18692
rect 12529 18683 12587 18689
rect 12529 18680 12541 18683
rect 12492 18652 12541 18680
rect 12492 18640 12498 18652
rect 12529 18649 12541 18652
rect 12575 18680 12587 18683
rect 14200 18680 14228 18720
rect 14734 18708 14740 18720
rect 14792 18708 14798 18760
rect 15194 18708 15200 18760
rect 15252 18748 15258 18760
rect 15289 18751 15347 18757
rect 15289 18748 15301 18751
rect 15252 18720 15301 18748
rect 15252 18708 15258 18720
rect 15289 18717 15301 18720
rect 15335 18748 15347 18751
rect 15470 18748 15476 18760
rect 15335 18720 15476 18748
rect 15335 18717 15347 18720
rect 15289 18711 15347 18717
rect 15470 18708 15476 18720
rect 15528 18708 15534 18760
rect 17972 18757 18000 18788
rect 18432 18760 18460 18788
rect 18616 18788 21496 18816
rect 17957 18751 18015 18757
rect 17957 18717 17969 18751
rect 18003 18717 18015 18751
rect 17957 18711 18015 18717
rect 18049 18751 18107 18757
rect 18049 18717 18061 18751
rect 18095 18717 18107 18751
rect 18049 18711 18107 18717
rect 18233 18751 18291 18757
rect 18233 18717 18245 18751
rect 18279 18717 18291 18751
rect 18233 18711 18291 18717
rect 12575 18652 14228 18680
rect 12575 18649 12587 18652
rect 12529 18643 12587 18649
rect 14550 18640 14556 18692
rect 14608 18680 14614 18692
rect 14645 18683 14703 18689
rect 14645 18680 14657 18683
rect 14608 18652 14657 18680
rect 14608 18640 14614 18652
rect 14645 18649 14657 18652
rect 14691 18649 14703 18683
rect 14645 18643 14703 18649
rect 14861 18683 14919 18689
rect 14861 18649 14873 18683
rect 14907 18680 14919 18683
rect 15378 18680 15384 18692
rect 14907 18652 15384 18680
rect 14907 18649 14919 18652
rect 14861 18643 14919 18649
rect 15378 18640 15384 18652
rect 15436 18640 15442 18692
rect 11793 18615 11851 18621
rect 11793 18612 11805 18615
rect 11256 18584 11805 18612
rect 11793 18581 11805 18584
rect 11839 18581 11851 18615
rect 11793 18575 11851 18581
rect 12618 18572 12624 18624
rect 12676 18612 12682 18624
rect 12713 18615 12771 18621
rect 12713 18612 12725 18615
rect 12676 18584 12725 18612
rect 12676 18572 12682 18584
rect 12713 18581 12725 18584
rect 12759 18581 12771 18615
rect 12713 18575 12771 18581
rect 15013 18615 15071 18621
rect 15013 18581 15025 18615
rect 15059 18612 15071 18615
rect 15746 18612 15752 18624
rect 15059 18584 15752 18612
rect 15059 18581 15071 18584
rect 15013 18575 15071 18581
rect 15746 18572 15752 18584
rect 15804 18572 15810 18624
rect 17034 18572 17040 18624
rect 17092 18612 17098 18624
rect 17773 18615 17831 18621
rect 17773 18612 17785 18615
rect 17092 18584 17785 18612
rect 17092 18572 17098 18584
rect 17773 18581 17785 18584
rect 17819 18581 17831 18615
rect 18064 18612 18092 18711
rect 18248 18680 18276 18711
rect 18322 18708 18328 18760
rect 18380 18708 18386 18760
rect 18414 18708 18420 18760
rect 18472 18708 18478 18760
rect 18616 18757 18644 18788
rect 21468 18760 21496 18788
rect 18601 18751 18659 18757
rect 18601 18717 18613 18751
rect 18647 18717 18659 18751
rect 18601 18711 18659 18717
rect 18509 18683 18567 18689
rect 18509 18680 18521 18683
rect 18248 18652 18521 18680
rect 18509 18649 18521 18652
rect 18555 18649 18567 18683
rect 18509 18643 18567 18649
rect 18616 18612 18644 18711
rect 18690 18708 18696 18760
rect 18748 18708 18754 18760
rect 18874 18708 18880 18760
rect 18932 18708 18938 18760
rect 21450 18708 21456 18760
rect 21508 18708 21514 18760
rect 21726 18708 21732 18760
rect 21784 18748 21790 18760
rect 24670 18748 24676 18760
rect 21784 18720 24676 18748
rect 21784 18708 21790 18720
rect 24670 18708 24676 18720
rect 24728 18708 24734 18760
rect 19886 18640 19892 18692
rect 19944 18680 19950 18692
rect 20073 18683 20131 18689
rect 20073 18680 20085 18683
rect 19944 18652 20085 18680
rect 19944 18640 19950 18652
rect 20073 18649 20085 18652
rect 20119 18649 20131 18683
rect 20073 18643 20131 18649
rect 20257 18683 20315 18689
rect 20257 18649 20269 18683
rect 20303 18680 20315 18683
rect 20622 18680 20628 18692
rect 20303 18652 20628 18680
rect 20303 18649 20315 18652
rect 20257 18643 20315 18649
rect 20622 18640 20628 18652
rect 20680 18640 20686 18692
rect 22646 18640 22652 18692
rect 22704 18640 22710 18692
rect 22830 18640 22836 18692
rect 22888 18640 22894 18692
rect 23382 18640 23388 18692
rect 23440 18680 23446 18692
rect 23842 18680 23848 18692
rect 23440 18652 23848 18680
rect 23440 18640 23446 18652
rect 23842 18640 23848 18652
rect 23900 18640 23906 18692
rect 18064 18584 18644 18612
rect 18877 18615 18935 18621
rect 17773 18575 17831 18581
rect 18877 18581 18889 18615
rect 18923 18612 18935 18615
rect 19058 18612 19064 18624
rect 18923 18584 19064 18612
rect 18923 18581 18935 18584
rect 18877 18575 18935 18581
rect 19058 18572 19064 18584
rect 19116 18572 19122 18624
rect 21269 18615 21327 18621
rect 21269 18581 21281 18615
rect 21315 18612 21327 18615
rect 21450 18612 21456 18624
rect 21315 18584 21456 18612
rect 21315 18581 21327 18584
rect 21269 18575 21327 18581
rect 21450 18572 21456 18584
rect 21508 18572 21514 18624
rect 23566 18572 23572 18624
rect 23624 18612 23630 18624
rect 24026 18612 24032 18624
rect 23624 18584 24032 18612
rect 23624 18572 23630 18584
rect 24026 18572 24032 18584
rect 24084 18572 24090 18624
rect 1104 18522 27876 18544
rect 1104 18470 4874 18522
rect 4926 18470 4938 18522
rect 4990 18470 5002 18522
rect 5054 18470 5066 18522
rect 5118 18470 5130 18522
rect 5182 18470 27876 18522
rect 1104 18448 27876 18470
rect 4798 18368 4804 18420
rect 4856 18368 4862 18420
rect 4890 18368 4896 18420
rect 4948 18408 4954 18420
rect 5994 18408 6000 18420
rect 4948 18380 6000 18408
rect 4948 18368 4954 18380
rect 5994 18368 6000 18380
rect 6052 18368 6058 18420
rect 6178 18368 6184 18420
rect 6236 18408 6242 18420
rect 6533 18411 6591 18417
rect 6533 18408 6545 18411
rect 6236 18380 6545 18408
rect 6236 18368 6242 18380
rect 6533 18377 6545 18380
rect 6579 18408 6591 18411
rect 6579 18380 7144 18408
rect 6579 18377 6591 18380
rect 6533 18371 6591 18377
rect 6638 18340 6644 18352
rect 2332 18312 6644 18340
rect 2332 18284 2360 18312
rect 2225 18275 2283 18281
rect 2225 18241 2237 18275
rect 2271 18272 2283 18275
rect 2314 18272 2320 18284
rect 2271 18244 2320 18272
rect 2271 18241 2283 18244
rect 2225 18235 2283 18241
rect 2314 18232 2320 18244
rect 2372 18232 2378 18284
rect 2492 18275 2550 18281
rect 2492 18241 2504 18275
rect 2538 18272 2550 18275
rect 2866 18272 2872 18284
rect 2538 18244 2872 18272
rect 2538 18241 2550 18244
rect 2492 18235 2550 18241
rect 2866 18232 2872 18244
rect 2924 18232 2930 18284
rect 3050 18232 3056 18284
rect 3108 18272 3114 18284
rect 3697 18275 3755 18281
rect 3697 18272 3709 18275
rect 3108 18244 3709 18272
rect 3108 18232 3114 18244
rect 3697 18241 3709 18244
rect 3743 18241 3755 18275
rect 3697 18235 3755 18241
rect 3881 18275 3939 18281
rect 3881 18241 3893 18275
rect 3927 18241 3939 18275
rect 3881 18235 3939 18241
rect 3896 18204 3924 18235
rect 3970 18232 3976 18284
rect 4028 18272 4034 18284
rect 4065 18275 4123 18281
rect 4065 18272 4077 18275
rect 4028 18244 4077 18272
rect 4028 18232 4034 18244
rect 4065 18241 4077 18244
rect 4111 18241 4123 18275
rect 4065 18235 4123 18241
rect 4157 18275 4215 18281
rect 4157 18241 4169 18275
rect 4203 18241 4215 18275
rect 4157 18235 4215 18241
rect 4341 18275 4399 18281
rect 4341 18241 4353 18275
rect 4387 18272 4399 18275
rect 4890 18272 4896 18284
rect 4387 18244 4896 18272
rect 4387 18241 4399 18244
rect 4341 18235 4399 18241
rect 4172 18204 4200 18235
rect 3620 18176 4200 18204
rect 3620 18080 3648 18176
rect 3878 18096 3884 18148
rect 3936 18136 3942 18148
rect 4356 18136 4384 18235
rect 4890 18232 4896 18244
rect 4948 18232 4954 18284
rect 4985 18275 5043 18281
rect 4985 18241 4997 18275
rect 5031 18241 5043 18275
rect 4985 18235 5043 18241
rect 5077 18275 5135 18281
rect 5077 18241 5089 18275
rect 5123 18241 5135 18275
rect 5077 18235 5135 18241
rect 3936 18108 4384 18136
rect 3936 18096 3942 18108
rect 3602 18028 3608 18080
rect 3660 18028 3666 18080
rect 4154 18028 4160 18080
rect 4212 18068 4218 18080
rect 4249 18071 4307 18077
rect 4249 18068 4261 18071
rect 4212 18040 4261 18068
rect 4212 18028 4218 18040
rect 4249 18037 4261 18040
rect 4295 18037 4307 18071
rect 5000 18068 5028 18235
rect 5092 18136 5120 18235
rect 5166 18232 5172 18284
rect 5224 18232 5230 18284
rect 5258 18232 5264 18284
rect 5316 18281 5322 18284
rect 5552 18281 5580 18312
rect 6638 18300 6644 18312
rect 6696 18300 6702 18352
rect 6733 18343 6791 18349
rect 6733 18309 6745 18343
rect 6779 18340 6791 18343
rect 7009 18343 7067 18349
rect 7009 18340 7021 18343
rect 6779 18312 7021 18340
rect 6779 18309 6791 18312
rect 6733 18303 6791 18309
rect 7009 18309 7021 18312
rect 7055 18309 7067 18343
rect 7009 18303 7067 18309
rect 7116 18340 7144 18380
rect 9766 18368 9772 18420
rect 9824 18408 9830 18420
rect 9953 18411 10011 18417
rect 9953 18408 9965 18411
rect 9824 18380 9965 18408
rect 9824 18368 9830 18380
rect 9953 18377 9965 18380
rect 9999 18377 10011 18411
rect 9953 18371 10011 18377
rect 10318 18368 10324 18420
rect 10376 18368 10382 18420
rect 11514 18368 11520 18420
rect 11572 18408 11578 18420
rect 12342 18408 12348 18420
rect 11572 18380 12348 18408
rect 11572 18368 11578 18380
rect 12342 18368 12348 18380
rect 12400 18368 12406 18420
rect 19518 18368 19524 18420
rect 19576 18368 19582 18420
rect 20254 18368 20260 18420
rect 20312 18368 20318 18420
rect 24489 18411 24547 18417
rect 24489 18408 24501 18411
rect 20456 18380 24501 18408
rect 9401 18343 9459 18349
rect 9401 18340 9413 18343
rect 7116 18312 9413 18340
rect 5316 18275 5345 18281
rect 5333 18241 5345 18275
rect 5316 18235 5345 18241
rect 5537 18275 5595 18281
rect 5537 18241 5549 18275
rect 5583 18241 5595 18275
rect 5537 18235 5595 18241
rect 5316 18232 5322 18235
rect 5445 18207 5503 18213
rect 5445 18173 5457 18207
rect 5491 18204 5503 18207
rect 5718 18204 5724 18216
rect 5491 18176 5724 18204
rect 5491 18173 5503 18176
rect 5445 18167 5503 18173
rect 5718 18164 5724 18176
rect 5776 18204 5782 18216
rect 6748 18204 6776 18303
rect 7116 18281 7144 18312
rect 9401 18309 9413 18312
rect 9447 18340 9459 18343
rect 9447 18312 9904 18340
rect 9447 18309 9459 18312
rect 9401 18303 9459 18309
rect 7466 18281 7472 18284
rect 6825 18275 6883 18281
rect 6825 18241 6837 18275
rect 6871 18241 6883 18275
rect 6825 18235 6883 18241
rect 7101 18275 7159 18281
rect 7101 18241 7113 18275
rect 7147 18241 7159 18275
rect 7101 18235 7159 18241
rect 7460 18235 7472 18281
rect 5776 18176 6776 18204
rect 5776 18164 5782 18176
rect 5534 18136 5540 18148
rect 5092 18108 5540 18136
rect 5534 18096 5540 18108
rect 5592 18096 5598 18148
rect 5994 18096 6000 18148
rect 6052 18136 6058 18148
rect 6365 18139 6423 18145
rect 6365 18136 6377 18139
rect 6052 18108 6377 18136
rect 6052 18096 6058 18108
rect 6365 18105 6377 18108
rect 6411 18136 6423 18139
rect 6638 18136 6644 18148
rect 6411 18108 6644 18136
rect 6411 18105 6423 18108
rect 6365 18099 6423 18105
rect 6638 18096 6644 18108
rect 6696 18096 6702 18148
rect 6840 18136 6868 18235
rect 7466 18232 7472 18235
rect 7524 18232 7530 18284
rect 9306 18232 9312 18284
rect 9364 18272 9370 18284
rect 9876 18281 9904 18312
rect 9585 18275 9643 18281
rect 9585 18272 9597 18275
rect 9364 18244 9597 18272
rect 9364 18232 9370 18244
rect 9585 18241 9597 18244
rect 9631 18241 9643 18275
rect 9585 18235 9643 18241
rect 9861 18275 9919 18281
rect 9861 18241 9873 18275
rect 9907 18241 9919 18275
rect 9861 18235 9919 18241
rect 10042 18232 10048 18284
rect 10100 18232 10106 18284
rect 10229 18275 10287 18281
rect 10229 18241 10241 18275
rect 10275 18241 10287 18275
rect 10229 18235 10287 18241
rect 10413 18275 10471 18281
rect 10413 18241 10425 18275
rect 10459 18272 10471 18275
rect 11146 18272 11152 18284
rect 10459 18244 11152 18272
rect 10459 18241 10471 18244
rect 10413 18235 10471 18241
rect 7006 18164 7012 18216
rect 7064 18204 7070 18216
rect 7193 18207 7251 18213
rect 7193 18204 7205 18207
rect 7064 18176 7205 18204
rect 7064 18164 7070 18176
rect 7193 18173 7205 18176
rect 7239 18173 7251 18207
rect 7193 18167 7251 18173
rect 9217 18207 9275 18213
rect 9217 18173 9229 18207
rect 9263 18173 9275 18207
rect 9217 18167 9275 18173
rect 8573 18139 8631 18145
rect 6748 18108 7052 18136
rect 6086 18068 6092 18080
rect 5000 18040 6092 18068
rect 4249 18031 4307 18037
rect 6086 18028 6092 18040
rect 6144 18028 6150 18080
rect 6546 18028 6552 18080
rect 6604 18068 6610 18080
rect 6748 18068 6776 18108
rect 6604 18040 6776 18068
rect 6825 18071 6883 18077
rect 6604 18028 6610 18040
rect 6825 18037 6837 18071
rect 6871 18068 6883 18071
rect 6914 18068 6920 18080
rect 6871 18040 6920 18068
rect 6871 18037 6883 18040
rect 6825 18031 6883 18037
rect 6914 18028 6920 18040
rect 6972 18028 6978 18080
rect 7024 18068 7052 18108
rect 8573 18105 8585 18139
rect 8619 18136 8631 18139
rect 9232 18136 9260 18167
rect 9490 18164 9496 18216
rect 9548 18204 9554 18216
rect 9769 18207 9827 18213
rect 9769 18204 9781 18207
rect 9548 18176 9781 18204
rect 9548 18164 9554 18176
rect 9769 18173 9781 18176
rect 9815 18204 9827 18207
rect 10244 18204 10272 18235
rect 9815 18176 10272 18204
rect 9815 18173 9827 18176
rect 9769 18167 9827 18173
rect 10428 18136 10456 18235
rect 11146 18232 11152 18244
rect 11204 18232 11210 18284
rect 11885 18275 11943 18281
rect 11885 18241 11897 18275
rect 11931 18241 11943 18275
rect 11885 18235 11943 18241
rect 11900 18204 11928 18235
rect 11974 18232 11980 18284
rect 12032 18232 12038 18284
rect 12066 18232 12072 18284
rect 12124 18272 12130 18284
rect 12161 18275 12219 18281
rect 12161 18272 12173 18275
rect 12124 18244 12173 18272
rect 12124 18232 12130 18244
rect 12161 18241 12173 18244
rect 12207 18241 12219 18275
rect 12161 18235 12219 18241
rect 12263 18275 12321 18281
rect 12263 18241 12275 18275
rect 12309 18272 12321 18275
rect 12360 18272 12388 18368
rect 20456 18352 20484 18380
rect 24489 18377 24501 18380
rect 24535 18377 24547 18411
rect 24489 18371 24547 18377
rect 24670 18368 24676 18420
rect 24728 18368 24734 18420
rect 14093 18343 14151 18349
rect 14093 18309 14105 18343
rect 14139 18340 14151 18343
rect 14737 18343 14795 18349
rect 14737 18340 14749 18343
rect 14139 18312 14749 18340
rect 14139 18309 14151 18312
rect 14093 18303 14151 18309
rect 14737 18309 14749 18312
rect 14783 18340 14795 18343
rect 15010 18340 15016 18352
rect 14783 18312 15016 18340
rect 14783 18309 14795 18312
rect 14737 18303 14795 18309
rect 15010 18300 15016 18312
rect 15068 18300 15074 18352
rect 19058 18300 19064 18352
rect 19116 18300 19122 18352
rect 20438 18300 20444 18352
rect 20496 18300 20502 18352
rect 21637 18343 21695 18349
rect 21637 18309 21649 18343
rect 21683 18340 21695 18343
rect 21910 18340 21916 18352
rect 21683 18312 21916 18340
rect 21683 18309 21695 18312
rect 21637 18303 21695 18309
rect 21910 18300 21916 18312
rect 21968 18300 21974 18352
rect 23382 18300 23388 18352
rect 23440 18300 23446 18352
rect 25133 18343 25191 18349
rect 25133 18340 25145 18343
rect 24412 18312 25145 18340
rect 24412 18284 24440 18312
rect 25133 18309 25145 18312
rect 25179 18309 25191 18343
rect 25133 18303 25191 18309
rect 12309 18244 12388 18272
rect 12309 18241 12321 18244
rect 12263 18235 12321 18241
rect 16758 18232 16764 18284
rect 16816 18272 16822 18284
rect 16925 18275 16983 18281
rect 16925 18272 16937 18275
rect 16816 18244 16937 18272
rect 16816 18232 16822 18244
rect 16925 18241 16937 18244
rect 16971 18241 16983 18275
rect 16925 18235 16983 18241
rect 18782 18232 18788 18284
rect 18840 18272 18846 18284
rect 18877 18275 18935 18281
rect 18877 18272 18889 18275
rect 18840 18244 18889 18272
rect 18840 18232 18846 18244
rect 18877 18241 18889 18244
rect 18923 18241 18935 18275
rect 18877 18235 18935 18241
rect 19153 18275 19211 18281
rect 19153 18241 19165 18275
rect 19199 18241 19211 18275
rect 19153 18235 19211 18241
rect 19245 18275 19303 18281
rect 19245 18241 19257 18275
rect 19291 18272 19303 18275
rect 20070 18272 20076 18284
rect 19291 18244 20076 18272
rect 19291 18241 19303 18244
rect 19245 18235 19303 18241
rect 12986 18204 12992 18216
rect 11900 18176 12992 18204
rect 12986 18164 12992 18176
rect 13044 18164 13050 18216
rect 16298 18204 16304 18216
rect 16040 18176 16304 18204
rect 8619 18108 10456 18136
rect 8619 18105 8631 18108
rect 8573 18099 8631 18105
rect 8588 18068 8616 18099
rect 7024 18040 8616 18068
rect 8662 18028 8668 18080
rect 8720 18028 8726 18080
rect 10502 18028 10508 18080
rect 10560 18068 10566 18080
rect 11701 18071 11759 18077
rect 11701 18068 11713 18071
rect 10560 18040 11713 18068
rect 10560 18028 10566 18040
rect 11701 18037 11713 18040
rect 11747 18037 11759 18071
rect 11701 18031 11759 18037
rect 12621 18071 12679 18077
rect 12621 18037 12633 18071
rect 12667 18068 12679 18071
rect 12710 18068 12716 18080
rect 12667 18040 12716 18068
rect 12667 18037 12679 18040
rect 12621 18031 12679 18037
rect 12710 18028 12716 18040
rect 12768 18028 12774 18080
rect 15470 18028 15476 18080
rect 15528 18068 15534 18080
rect 16040 18077 16068 18176
rect 16298 18164 16304 18176
rect 16356 18204 16362 18216
rect 16669 18207 16727 18213
rect 16669 18204 16681 18207
rect 16356 18176 16681 18204
rect 16356 18164 16362 18176
rect 16669 18173 16681 18176
rect 16715 18173 16727 18207
rect 16669 18167 16727 18173
rect 16025 18071 16083 18077
rect 16025 18068 16037 18071
rect 15528 18040 16037 18068
rect 15528 18028 15534 18040
rect 16025 18037 16037 18040
rect 16071 18037 16083 18071
rect 16684 18068 16712 18167
rect 18046 18164 18052 18216
rect 18104 18204 18110 18216
rect 18141 18207 18199 18213
rect 18141 18204 18153 18207
rect 18104 18176 18153 18204
rect 18104 18164 18110 18176
rect 18141 18173 18153 18176
rect 18187 18173 18199 18207
rect 18141 18167 18199 18173
rect 18693 18207 18751 18213
rect 18693 18173 18705 18207
rect 18739 18173 18751 18207
rect 18693 18167 18751 18173
rect 17678 18096 17684 18148
rect 17736 18136 17742 18148
rect 18708 18136 18736 18167
rect 17736 18108 18736 18136
rect 19168 18136 19196 18235
rect 20070 18232 20076 18244
rect 20128 18232 20134 18284
rect 20165 18275 20223 18281
rect 20165 18241 20177 18275
rect 20211 18241 20223 18275
rect 21818 18272 21824 18284
rect 21298 18244 21824 18272
rect 20165 18235 20223 18241
rect 19334 18164 19340 18216
rect 19392 18204 19398 18216
rect 19794 18204 19800 18216
rect 19392 18176 19800 18204
rect 19392 18164 19398 18176
rect 19794 18164 19800 18176
rect 19852 18164 19858 18216
rect 19886 18164 19892 18216
rect 19944 18204 19950 18216
rect 20180 18204 20208 18235
rect 21818 18232 21824 18244
rect 21876 18232 21882 18284
rect 22370 18232 22376 18284
rect 22428 18232 22434 18284
rect 22830 18232 22836 18284
rect 22888 18232 22894 18284
rect 23566 18232 23572 18284
rect 23624 18232 23630 18284
rect 23750 18232 23756 18284
rect 23808 18232 23814 18284
rect 23842 18232 23848 18284
rect 23900 18232 23906 18284
rect 24394 18232 24400 18284
rect 24452 18232 24458 18284
rect 24581 18275 24639 18281
rect 24581 18241 24593 18275
rect 24627 18241 24639 18275
rect 24581 18235 24639 18241
rect 24857 18275 24915 18281
rect 24857 18241 24869 18275
rect 24903 18272 24915 18275
rect 24946 18272 24952 18284
rect 24903 18244 24952 18272
rect 24903 18241 24915 18244
rect 24857 18235 24915 18241
rect 19944 18176 20208 18204
rect 19944 18164 19950 18176
rect 20806 18164 20812 18216
rect 20864 18164 20870 18216
rect 23658 18164 23664 18216
rect 23716 18164 23722 18216
rect 24596 18204 24624 18235
rect 24946 18232 24952 18244
rect 25004 18272 25010 18284
rect 25409 18275 25467 18281
rect 25409 18272 25421 18275
rect 25004 18244 25421 18272
rect 25004 18232 25010 18244
rect 25409 18241 25421 18244
rect 25455 18241 25467 18275
rect 25409 18235 25467 18241
rect 25590 18232 25596 18284
rect 25648 18232 25654 18284
rect 25038 18204 25044 18216
rect 24596 18176 25044 18204
rect 25038 18164 25044 18176
rect 25096 18164 25102 18216
rect 25225 18139 25283 18145
rect 25225 18136 25237 18139
rect 19168 18108 23612 18136
rect 17736 18096 17742 18108
rect 17954 18068 17960 18080
rect 16684 18040 17960 18068
rect 16025 18031 16083 18037
rect 17954 18028 17960 18040
rect 18012 18028 18018 18080
rect 18064 18077 18092 18108
rect 18049 18071 18107 18077
rect 18049 18037 18061 18071
rect 18095 18037 18107 18071
rect 18049 18031 18107 18037
rect 19426 18028 19432 18080
rect 19484 18028 19490 18080
rect 19981 18071 20039 18077
rect 19981 18037 19993 18071
rect 20027 18068 20039 18071
rect 20441 18071 20499 18077
rect 20441 18068 20453 18071
rect 20027 18040 20453 18068
rect 20027 18037 20039 18040
rect 19981 18031 20039 18037
rect 20441 18037 20453 18040
rect 20487 18037 20499 18071
rect 23584 18068 23612 18108
rect 23768 18108 25237 18136
rect 23768 18068 23796 18108
rect 25225 18105 25237 18108
rect 25271 18105 25283 18139
rect 25225 18099 25283 18105
rect 23584 18040 23796 18068
rect 24029 18071 24087 18077
rect 20441 18031 20499 18037
rect 24029 18037 24041 18071
rect 24075 18068 24087 18071
rect 24578 18068 24584 18080
rect 24075 18040 24584 18068
rect 24075 18037 24087 18040
rect 24029 18031 24087 18037
rect 24578 18028 24584 18040
rect 24636 18028 24642 18080
rect 25133 18071 25191 18077
rect 25133 18037 25145 18071
rect 25179 18068 25191 18071
rect 25590 18068 25596 18080
rect 25179 18040 25596 18068
rect 25179 18037 25191 18040
rect 25133 18031 25191 18037
rect 25590 18028 25596 18040
rect 25648 18028 25654 18080
rect 1104 17978 27876 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 27876 17978
rect 1104 17904 27876 17926
rect 2777 17867 2835 17873
rect 2777 17833 2789 17867
rect 2823 17864 2835 17867
rect 2866 17864 2872 17876
rect 2823 17836 2872 17864
rect 2823 17833 2835 17836
rect 2777 17827 2835 17833
rect 2866 17824 2872 17836
rect 2924 17824 2930 17876
rect 5258 17864 5264 17876
rect 4540 17836 5264 17864
rect 4062 17728 4068 17740
rect 2976 17700 4068 17728
rect 2976 17669 3004 17700
rect 4062 17688 4068 17700
rect 4120 17688 4126 17740
rect 2961 17663 3019 17669
rect 2961 17629 2973 17663
rect 3007 17629 3019 17663
rect 2961 17623 3019 17629
rect 3050 17620 3056 17672
rect 3108 17620 3114 17672
rect 3421 17663 3479 17669
rect 3421 17629 3433 17663
rect 3467 17660 3479 17663
rect 3602 17660 3608 17672
rect 3467 17632 3608 17660
rect 3467 17629 3479 17632
rect 3421 17623 3479 17629
rect 3602 17620 3608 17632
rect 3660 17660 3666 17672
rect 4154 17660 4160 17672
rect 3660 17632 4160 17660
rect 3660 17620 3666 17632
rect 4154 17620 4160 17632
rect 4212 17620 4218 17672
rect 2314 17552 2320 17604
rect 2372 17592 2378 17604
rect 3145 17595 3203 17601
rect 3145 17592 3157 17595
rect 2372 17564 3157 17592
rect 2372 17552 2378 17564
rect 3145 17561 3157 17564
rect 3191 17561 3203 17595
rect 3145 17555 3203 17561
rect 3283 17595 3341 17601
rect 3283 17561 3295 17595
rect 3329 17592 3341 17595
rect 4540 17592 4568 17836
rect 5258 17824 5264 17836
rect 5316 17824 5322 17876
rect 5534 17824 5540 17876
rect 5592 17824 5598 17876
rect 6086 17824 6092 17876
rect 6144 17824 6150 17876
rect 6730 17824 6736 17876
rect 6788 17864 6794 17876
rect 7098 17864 7104 17876
rect 6788 17836 7104 17864
rect 6788 17824 6794 17836
rect 7098 17824 7104 17836
rect 7156 17824 7162 17876
rect 7377 17867 7435 17873
rect 7377 17833 7389 17867
rect 7423 17864 7435 17867
rect 7466 17864 7472 17876
rect 7423 17836 7472 17864
rect 7423 17833 7435 17836
rect 7377 17827 7435 17833
rect 7466 17824 7472 17836
rect 7524 17824 7530 17876
rect 9677 17867 9735 17873
rect 9677 17833 9689 17867
rect 9723 17864 9735 17867
rect 9950 17864 9956 17876
rect 9723 17836 9956 17864
rect 9723 17833 9735 17836
rect 9677 17827 9735 17833
rect 9950 17824 9956 17836
rect 10008 17824 10014 17876
rect 10321 17867 10379 17873
rect 10321 17833 10333 17867
rect 10367 17864 10379 17867
rect 10686 17864 10692 17876
rect 10367 17836 10692 17864
rect 10367 17833 10379 17836
rect 10321 17827 10379 17833
rect 10686 17824 10692 17836
rect 10744 17824 10750 17876
rect 11149 17867 11207 17873
rect 11149 17833 11161 17867
rect 11195 17833 11207 17867
rect 11149 17827 11207 17833
rect 4893 17799 4951 17805
rect 4893 17765 4905 17799
rect 4939 17796 4951 17799
rect 9401 17799 9459 17805
rect 4939 17768 9260 17796
rect 4939 17765 4951 17768
rect 4893 17759 4951 17765
rect 5166 17728 5172 17740
rect 3329 17564 4568 17592
rect 4632 17700 5172 17728
rect 3329 17561 3341 17564
rect 3283 17555 3341 17561
rect 3160 17524 3188 17555
rect 4632 17524 4660 17700
rect 5166 17688 5172 17700
rect 5224 17728 5230 17740
rect 6733 17731 6791 17737
rect 5224 17700 6316 17728
rect 5224 17688 5230 17700
rect 4709 17663 4767 17669
rect 4709 17629 4721 17663
rect 4755 17629 4767 17663
rect 4709 17623 4767 17629
rect 4724 17592 4752 17623
rect 4798 17620 4804 17672
rect 4856 17660 4862 17672
rect 4893 17663 4951 17669
rect 4893 17660 4905 17663
rect 4856 17632 4905 17660
rect 4856 17620 4862 17632
rect 4893 17629 4905 17632
rect 4939 17629 4951 17663
rect 5997 17663 6055 17669
rect 5997 17660 6009 17663
rect 4893 17623 4951 17629
rect 5736 17632 6009 17660
rect 5736 17604 5764 17632
rect 5997 17629 6009 17632
rect 6043 17629 6055 17663
rect 5997 17623 6055 17629
rect 6178 17620 6184 17672
rect 6236 17620 6242 17672
rect 5258 17592 5264 17604
rect 4724 17564 5264 17592
rect 5258 17552 5264 17564
rect 5316 17552 5322 17604
rect 5718 17552 5724 17604
rect 5776 17552 5782 17604
rect 5905 17595 5963 17601
rect 5905 17561 5917 17595
rect 5951 17592 5963 17595
rect 6196 17592 6224 17620
rect 5951 17564 6224 17592
rect 6288 17592 6316 17700
rect 6733 17697 6745 17731
rect 6779 17728 6791 17731
rect 8021 17731 8079 17737
rect 6779 17700 7604 17728
rect 6779 17697 6791 17700
rect 6733 17691 6791 17697
rect 6638 17620 6644 17672
rect 6696 17620 6702 17672
rect 6825 17663 6883 17669
rect 6825 17629 6837 17663
rect 6871 17660 6883 17663
rect 6914 17660 6920 17672
rect 6871 17632 6920 17660
rect 6871 17629 6883 17632
rect 6825 17623 6883 17629
rect 6914 17620 6920 17632
rect 6972 17620 6978 17672
rect 7576 17669 7604 17700
rect 8021 17697 8033 17731
rect 8067 17728 8079 17731
rect 8662 17728 8668 17740
rect 8067 17700 8668 17728
rect 8067 17697 8079 17700
rect 8021 17691 8079 17697
rect 8662 17688 8668 17700
rect 8720 17688 8726 17740
rect 9232 17728 9260 17768
rect 9401 17765 9413 17799
rect 9447 17796 9459 17799
rect 10042 17796 10048 17808
rect 9447 17768 10048 17796
rect 9447 17765 9459 17768
rect 9401 17759 9459 17765
rect 10042 17756 10048 17768
rect 10100 17756 10106 17808
rect 10226 17756 10232 17808
rect 10284 17796 10290 17808
rect 10781 17799 10839 17805
rect 10781 17796 10793 17799
rect 10284 17768 10793 17796
rect 10284 17756 10290 17768
rect 10781 17765 10793 17768
rect 10827 17765 10839 17799
rect 11164 17796 11192 17827
rect 11606 17824 11612 17876
rect 11664 17864 11670 17876
rect 11793 17867 11851 17873
rect 11793 17864 11805 17867
rect 11664 17836 11805 17864
rect 11664 17824 11670 17836
rect 11793 17833 11805 17836
rect 11839 17833 11851 17867
rect 11793 17827 11851 17833
rect 12986 17824 12992 17876
rect 13044 17824 13050 17876
rect 13449 17867 13507 17873
rect 13449 17833 13461 17867
rect 13495 17864 13507 17867
rect 13538 17864 13544 17876
rect 13495 17836 13544 17864
rect 13495 17833 13507 17836
rect 13449 17827 13507 17833
rect 13538 17824 13544 17836
rect 13596 17824 13602 17876
rect 16022 17864 16028 17876
rect 15488 17836 16028 17864
rect 12618 17796 12624 17808
rect 11164 17768 12624 17796
rect 10781 17759 10839 17765
rect 12618 17756 12624 17768
rect 12676 17756 12682 17808
rect 15286 17756 15292 17808
rect 15344 17796 15350 17808
rect 15488 17805 15516 17836
rect 16022 17824 16028 17836
rect 16080 17824 16086 17876
rect 16758 17824 16764 17876
rect 16816 17824 16822 17876
rect 18049 17867 18107 17873
rect 18049 17833 18061 17867
rect 18095 17833 18107 17867
rect 18049 17827 18107 17833
rect 18325 17867 18383 17873
rect 18325 17833 18337 17867
rect 18371 17864 18383 17867
rect 18414 17864 18420 17876
rect 18371 17836 18420 17864
rect 18371 17833 18383 17836
rect 18325 17827 18383 17833
rect 15473 17799 15531 17805
rect 15473 17796 15485 17799
rect 15344 17768 15485 17796
rect 15344 17756 15350 17768
rect 15473 17765 15485 17768
rect 15519 17765 15531 17799
rect 18064 17796 18092 17827
rect 18414 17824 18420 17836
rect 18472 17824 18478 17876
rect 20070 17824 20076 17876
rect 20128 17864 20134 17876
rect 20165 17867 20223 17873
rect 20165 17864 20177 17867
rect 20128 17836 20177 17864
rect 20128 17824 20134 17836
rect 20165 17833 20177 17836
rect 20211 17833 20223 17867
rect 20165 17827 20223 17833
rect 22830 17824 22836 17876
rect 22888 17824 22894 17876
rect 23017 17867 23075 17873
rect 23017 17833 23029 17867
rect 23063 17864 23075 17867
rect 23658 17864 23664 17876
rect 23063 17836 23664 17864
rect 23063 17833 23075 17836
rect 23017 17827 23075 17833
rect 23658 17824 23664 17836
rect 23716 17824 23722 17876
rect 24394 17824 24400 17876
rect 24452 17824 24458 17876
rect 24578 17824 24584 17876
rect 24636 17824 24642 17876
rect 25038 17824 25044 17876
rect 25096 17864 25102 17876
rect 25225 17867 25283 17873
rect 25225 17864 25237 17867
rect 25096 17836 25237 17864
rect 25096 17824 25102 17836
rect 25225 17833 25237 17836
rect 25271 17833 25283 17867
rect 25225 17827 25283 17833
rect 19242 17796 19248 17808
rect 15473 17759 15531 17765
rect 15764 17768 16344 17796
rect 9232 17700 9536 17728
rect 7561 17663 7619 17669
rect 7561 17629 7573 17663
rect 7607 17629 7619 17663
rect 7561 17623 7619 17629
rect 7650 17620 7656 17672
rect 7708 17620 7714 17672
rect 8938 17620 8944 17672
rect 8996 17660 9002 17672
rect 9217 17663 9275 17669
rect 9217 17660 9229 17663
rect 8996 17632 9229 17660
rect 8996 17620 9002 17632
rect 9217 17629 9229 17632
rect 9263 17629 9275 17663
rect 9217 17623 9275 17629
rect 9306 17620 9312 17672
rect 9364 17660 9370 17672
rect 9401 17663 9459 17669
rect 9401 17660 9413 17663
rect 9364 17632 9413 17660
rect 9364 17620 9370 17632
rect 9401 17629 9413 17632
rect 9447 17629 9459 17663
rect 9508 17660 9536 17700
rect 9582 17688 9588 17740
rect 9640 17688 9646 17740
rect 9769 17731 9827 17737
rect 9769 17697 9781 17731
rect 9815 17728 9827 17731
rect 9953 17731 10011 17737
rect 9953 17728 9965 17731
rect 9815 17700 9965 17728
rect 9815 17697 9827 17700
rect 9769 17691 9827 17697
rect 9953 17697 9965 17700
rect 9999 17697 10011 17731
rect 11057 17731 11115 17737
rect 11057 17728 11069 17731
rect 9953 17691 10011 17697
rect 10152 17700 11069 17728
rect 9674 17660 9680 17672
rect 9508 17632 9680 17660
rect 9401 17623 9459 17629
rect 9674 17620 9680 17632
rect 9732 17620 9738 17672
rect 9861 17663 9919 17669
rect 9861 17629 9873 17663
rect 9907 17660 9919 17663
rect 10152 17660 10180 17700
rect 11057 17697 11069 17700
rect 11103 17728 11115 17731
rect 11238 17728 11244 17740
rect 11103 17700 11244 17728
rect 11103 17697 11115 17700
rect 11057 17691 11115 17697
rect 11238 17688 11244 17700
rect 11296 17688 11302 17740
rect 12894 17728 12900 17740
rect 12406 17700 12900 17728
rect 9907 17632 10180 17660
rect 10229 17663 10287 17669
rect 9907 17629 9919 17632
rect 9861 17623 9919 17629
rect 10229 17629 10241 17663
rect 10275 17629 10287 17663
rect 10229 17623 10287 17629
rect 10413 17663 10471 17669
rect 10413 17629 10425 17663
rect 10459 17629 10471 17663
rect 10413 17623 10471 17629
rect 7668 17592 7696 17620
rect 6288 17564 7696 17592
rect 7745 17595 7803 17601
rect 5951 17561 5963 17564
rect 5905 17555 5963 17561
rect 7745 17561 7757 17595
rect 7791 17561 7803 17595
rect 7745 17555 7803 17561
rect 3160 17496 4660 17524
rect 4706 17484 4712 17536
rect 4764 17524 4770 17536
rect 5736 17524 5764 17552
rect 4764 17496 5764 17524
rect 7760 17524 7788 17555
rect 7834 17552 7840 17604
rect 7892 17601 7898 17604
rect 7892 17595 7921 17601
rect 7909 17561 7921 17595
rect 7892 17555 7921 17561
rect 7892 17552 7898 17555
rect 9490 17552 9496 17604
rect 9548 17592 9554 17604
rect 10244 17592 10272 17623
rect 9548 17564 10272 17592
rect 10428 17592 10456 17623
rect 10502 17620 10508 17672
rect 10560 17660 10566 17672
rect 10626 17663 10684 17669
rect 10626 17660 10638 17663
rect 10560 17632 10638 17660
rect 10560 17620 10566 17632
rect 10626 17629 10638 17632
rect 10672 17629 10684 17663
rect 10626 17623 10684 17629
rect 11149 17663 11207 17669
rect 11149 17629 11161 17663
rect 11195 17629 11207 17663
rect 11149 17623 11207 17629
rect 11977 17663 12035 17669
rect 11977 17629 11989 17663
rect 12023 17660 12035 17663
rect 12158 17660 12164 17672
rect 12023 17632 12164 17660
rect 12023 17629 12035 17632
rect 11977 17623 12035 17629
rect 11164 17592 11192 17623
rect 12158 17620 12164 17632
rect 12216 17660 12222 17672
rect 12406 17660 12434 17700
rect 12894 17688 12900 17700
rect 12952 17688 12958 17740
rect 14274 17688 14280 17740
rect 14332 17728 14338 17740
rect 15764 17728 15792 17768
rect 14332 17700 15792 17728
rect 14332 17688 14338 17700
rect 15838 17688 15844 17740
rect 15896 17688 15902 17740
rect 12216 17632 12434 17660
rect 12216 17620 12222 17632
rect 12710 17620 12716 17672
rect 12768 17620 12774 17672
rect 13170 17620 13176 17672
rect 13228 17620 13234 17672
rect 13541 17663 13599 17669
rect 13541 17629 13553 17663
rect 13587 17629 13599 17663
rect 13541 17623 13599 17629
rect 10428 17564 11192 17592
rect 9548 17552 9554 17564
rect 9030 17524 9036 17536
rect 7760 17496 9036 17524
rect 4764 17484 4770 17496
rect 9030 17484 9036 17496
rect 9088 17484 9094 17536
rect 9398 17484 9404 17536
rect 9456 17524 9462 17536
rect 10428 17524 10456 17564
rect 11698 17552 11704 17604
rect 11756 17552 11762 17604
rect 11885 17595 11943 17601
rect 11885 17561 11897 17595
rect 11931 17592 11943 17595
rect 13078 17592 13084 17604
rect 11931 17564 13084 17592
rect 11931 17561 11943 17564
rect 11885 17555 11943 17561
rect 13078 17552 13084 17564
rect 13136 17552 13142 17604
rect 9456 17496 10456 17524
rect 10597 17527 10655 17533
rect 9456 17484 9462 17496
rect 10597 17493 10609 17527
rect 10643 17524 10655 17527
rect 10870 17524 10876 17536
rect 10643 17496 10876 17524
rect 10643 17493 10655 17496
rect 10597 17487 10655 17493
rect 10870 17484 10876 17496
rect 10928 17524 10934 17536
rect 13262 17524 13268 17536
rect 10928 17496 13268 17524
rect 10928 17484 10934 17496
rect 13262 17484 13268 17496
rect 13320 17524 13326 17536
rect 13556 17524 13584 17623
rect 13906 17620 13912 17672
rect 13964 17660 13970 17672
rect 14093 17663 14151 17669
rect 14093 17660 14105 17663
rect 13964 17632 14105 17660
rect 13964 17620 13970 17632
rect 14093 17629 14105 17632
rect 14139 17629 14151 17663
rect 14093 17623 14151 17629
rect 14369 17663 14427 17669
rect 14369 17629 14381 17663
rect 14415 17660 14427 17663
rect 14734 17660 14740 17672
rect 14415 17632 14740 17660
rect 14415 17629 14427 17632
rect 14369 17623 14427 17629
rect 14734 17620 14740 17632
rect 14792 17620 14798 17672
rect 15194 17620 15200 17672
rect 15252 17660 15258 17672
rect 16117 17663 16175 17669
rect 16117 17660 16129 17663
rect 15252 17632 16129 17660
rect 15252 17620 15258 17632
rect 16117 17629 16129 17632
rect 16163 17660 16175 17663
rect 16206 17660 16212 17672
rect 16163 17632 16212 17660
rect 16163 17629 16175 17632
rect 16117 17623 16175 17629
rect 16206 17620 16212 17632
rect 16264 17620 16270 17672
rect 16316 17660 16344 17768
rect 16960 17768 18092 17796
rect 18156 17768 19248 17796
rect 16960 17669 16988 17768
rect 17405 17731 17463 17737
rect 17405 17697 17417 17731
rect 17451 17728 17463 17731
rect 18046 17728 18052 17740
rect 17451 17700 18052 17728
rect 17451 17697 17463 17700
rect 17405 17691 17463 17697
rect 18046 17688 18052 17700
rect 18104 17688 18110 17740
rect 18156 17737 18184 17768
rect 19242 17756 19248 17768
rect 19300 17756 19306 17808
rect 18141 17731 18199 17737
rect 18141 17697 18153 17731
rect 18187 17697 18199 17731
rect 18690 17728 18696 17740
rect 18141 17691 18199 17697
rect 18248 17700 18696 17728
rect 16945 17663 17003 17669
rect 16316 17632 16436 17660
rect 16298 17592 16304 17604
rect 15488 17564 16304 17592
rect 15488 17524 15516 17564
rect 16298 17552 16304 17564
rect 16356 17552 16362 17604
rect 16408 17592 16436 17632
rect 16945 17629 16957 17663
rect 16991 17629 17003 17663
rect 16945 17623 17003 17629
rect 17034 17620 17040 17672
rect 17092 17620 17098 17672
rect 17126 17620 17132 17672
rect 17184 17620 17190 17672
rect 17247 17663 17305 17669
rect 17247 17629 17259 17663
rect 17293 17660 17305 17663
rect 17586 17660 17592 17672
rect 17293 17632 17592 17660
rect 17293 17629 17305 17632
rect 17247 17623 17305 17629
rect 17262 17592 17290 17623
rect 17586 17620 17592 17632
rect 17644 17620 17650 17672
rect 17678 17620 17684 17672
rect 17736 17660 17742 17672
rect 17773 17663 17831 17669
rect 17773 17660 17785 17663
rect 17736 17632 17785 17660
rect 17736 17620 17742 17632
rect 17773 17629 17785 17632
rect 17819 17629 17831 17663
rect 17773 17623 17831 17629
rect 17862 17620 17868 17672
rect 17920 17620 17926 17672
rect 18248 17669 18276 17700
rect 18690 17688 18696 17700
rect 18748 17688 18754 17740
rect 17957 17663 18015 17669
rect 17957 17629 17969 17663
rect 18003 17629 18015 17663
rect 17957 17623 18015 17629
rect 18233 17663 18291 17669
rect 18233 17629 18245 17663
rect 18279 17629 18291 17663
rect 18233 17623 18291 17629
rect 18417 17663 18475 17669
rect 18417 17629 18429 17663
rect 18463 17660 18475 17663
rect 19886 17660 19892 17672
rect 18463 17632 19892 17660
rect 18463 17629 18475 17632
rect 18417 17623 18475 17629
rect 16408 17564 17290 17592
rect 17402 17552 17408 17604
rect 17460 17592 17466 17604
rect 17972 17592 18000 17623
rect 19886 17620 19892 17632
rect 19944 17620 19950 17672
rect 20165 17663 20223 17669
rect 20165 17629 20177 17663
rect 20211 17660 20223 17663
rect 20438 17660 20444 17672
rect 20211 17632 20444 17660
rect 20211 17629 20223 17632
rect 20165 17623 20223 17629
rect 20438 17620 20444 17632
rect 20496 17620 20502 17672
rect 22646 17620 22652 17672
rect 22704 17620 22710 17672
rect 22833 17663 22891 17669
rect 22833 17629 22845 17663
rect 22879 17660 22891 17663
rect 23014 17660 23020 17672
rect 22879 17632 23020 17660
rect 22879 17629 22891 17632
rect 22833 17623 22891 17629
rect 23014 17620 23020 17632
rect 23072 17620 23078 17672
rect 24578 17620 24584 17672
rect 24636 17620 24642 17672
rect 24854 17620 24860 17672
rect 24912 17660 24918 17672
rect 24949 17663 25007 17669
rect 24949 17660 24961 17663
rect 24912 17632 24961 17660
rect 24912 17620 24918 17632
rect 24949 17629 24961 17632
rect 24995 17660 25007 17663
rect 25041 17663 25099 17669
rect 25041 17660 25053 17663
rect 24995 17632 25053 17660
rect 24995 17629 25007 17632
rect 24949 17623 25007 17629
rect 25041 17629 25053 17632
rect 25087 17629 25099 17663
rect 25041 17623 25099 17629
rect 25501 17663 25559 17669
rect 25501 17629 25513 17663
rect 25547 17629 25559 17663
rect 25501 17623 25559 17629
rect 17460 17564 18000 17592
rect 20073 17595 20131 17601
rect 17460 17552 17466 17564
rect 20073 17561 20085 17595
rect 20119 17592 20131 17595
rect 20254 17592 20260 17604
rect 20119 17564 20260 17592
rect 20119 17561 20131 17564
rect 20073 17555 20131 17561
rect 20254 17552 20260 17564
rect 20312 17552 20318 17604
rect 22664 17592 22692 17620
rect 23198 17592 23204 17604
rect 22664 17564 23204 17592
rect 23198 17552 23204 17564
rect 23256 17552 23262 17604
rect 23290 17552 23296 17604
rect 23348 17592 23354 17604
rect 24596 17592 24624 17620
rect 25409 17595 25467 17601
rect 25409 17592 25421 17595
rect 23348 17564 24440 17592
rect 24596 17564 25421 17592
rect 23348 17552 23354 17564
rect 13320 17496 15516 17524
rect 13320 17484 13326 17496
rect 15562 17484 15568 17536
rect 15620 17524 15626 17536
rect 16114 17524 16120 17536
rect 15620 17496 16120 17524
rect 15620 17484 15626 17496
rect 16114 17484 16120 17496
rect 16172 17484 16178 17536
rect 16316 17524 16344 17552
rect 17589 17527 17647 17533
rect 17589 17524 17601 17527
rect 16316 17496 17601 17524
rect 17589 17493 17601 17496
rect 17635 17493 17647 17527
rect 17589 17487 17647 17493
rect 22186 17484 22192 17536
rect 22244 17524 22250 17536
rect 23658 17524 23664 17536
rect 22244 17496 23664 17524
rect 22244 17484 22250 17496
rect 23658 17484 23664 17496
rect 23716 17484 23722 17536
rect 24412 17524 24440 17564
rect 25409 17561 25421 17564
rect 25455 17561 25467 17595
rect 25409 17555 25467 17561
rect 24581 17527 24639 17533
rect 24581 17524 24593 17527
rect 24412 17496 24593 17524
rect 24581 17493 24593 17496
rect 24627 17524 24639 17527
rect 25516 17524 25544 17623
rect 25774 17524 25780 17536
rect 24627 17496 25780 17524
rect 24627 17493 24639 17496
rect 24581 17487 24639 17493
rect 25774 17484 25780 17496
rect 25832 17484 25838 17536
rect 1104 17434 27876 17456
rect 1104 17382 4874 17434
rect 4926 17382 4938 17434
rect 4990 17382 5002 17434
rect 5054 17382 5066 17434
rect 5118 17382 5130 17434
rect 5182 17382 27876 17434
rect 1104 17360 27876 17382
rect 3973 17323 4031 17329
rect 3973 17289 3985 17323
rect 4019 17320 4031 17323
rect 4154 17320 4160 17332
rect 4019 17292 4160 17320
rect 4019 17289 4031 17292
rect 3973 17283 4031 17289
rect 4154 17280 4160 17292
rect 4212 17280 4218 17332
rect 4798 17280 4804 17332
rect 4856 17320 4862 17332
rect 4893 17323 4951 17329
rect 4893 17320 4905 17323
rect 4856 17292 4905 17320
rect 4856 17280 4862 17292
rect 4893 17289 4905 17292
rect 4939 17289 4951 17323
rect 6733 17323 6791 17329
rect 6733 17320 6745 17323
rect 4893 17283 4951 17289
rect 5092 17292 6745 17320
rect 3804 17224 4568 17252
rect 1664 17187 1722 17193
rect 1664 17153 1676 17187
rect 1710 17184 1722 17187
rect 1946 17184 1952 17196
rect 1710 17156 1952 17184
rect 1710 17153 1722 17156
rect 1664 17147 1722 17153
rect 1946 17144 1952 17156
rect 2004 17144 2010 17196
rect 3804 17193 3832 17224
rect 3789 17187 3847 17193
rect 3789 17153 3801 17187
rect 3835 17153 3847 17187
rect 3789 17147 3847 17153
rect 1397 17119 1455 17125
rect 1397 17085 1409 17119
rect 1443 17085 1455 17119
rect 3234 17116 3240 17128
rect 1397 17079 1455 17085
rect 2792 17088 3240 17116
rect 1412 16980 1440 17079
rect 2792 17057 2820 17088
rect 3234 17076 3240 17088
rect 3292 17116 3298 17128
rect 3421 17119 3479 17125
rect 3421 17116 3433 17119
rect 3292 17088 3433 17116
rect 3292 17076 3298 17088
rect 3421 17085 3433 17088
rect 3467 17116 3479 17119
rect 3804 17116 3832 17147
rect 4062 17144 4068 17196
rect 4120 17144 4126 17196
rect 4433 17187 4491 17193
rect 4433 17153 4445 17187
rect 4479 17153 4491 17187
rect 4433 17147 4491 17153
rect 3467 17088 3832 17116
rect 3467 17085 3479 17088
rect 3421 17079 3479 17085
rect 2777 17051 2835 17057
rect 2777 17017 2789 17051
rect 2823 17017 2835 17051
rect 4448 17048 4476 17147
rect 4540 17125 4568 17224
rect 4706 17144 4712 17196
rect 4764 17144 4770 17196
rect 4798 17144 4804 17196
rect 4856 17184 4862 17196
rect 5092 17193 5120 17292
rect 6733 17289 6745 17292
rect 6779 17289 6791 17323
rect 8110 17320 8116 17332
rect 6733 17283 6791 17289
rect 7208 17292 8116 17320
rect 4985 17187 5043 17193
rect 4985 17184 4997 17187
rect 4856 17156 4997 17184
rect 4856 17144 4862 17156
rect 4985 17153 4997 17156
rect 5031 17153 5043 17187
rect 4985 17147 5043 17153
rect 5077 17187 5135 17193
rect 5077 17153 5089 17187
rect 5123 17153 5135 17187
rect 5077 17147 5135 17153
rect 4525 17119 4583 17125
rect 4525 17085 4537 17119
rect 4571 17085 4583 17119
rect 4525 17079 4583 17085
rect 4614 17076 4620 17128
rect 4672 17116 4678 17128
rect 5092 17116 5120 17147
rect 5258 17144 5264 17196
rect 5316 17144 5322 17196
rect 5442 17144 5448 17196
rect 5500 17184 5506 17196
rect 5537 17187 5595 17193
rect 5537 17184 5549 17187
rect 5500 17156 5549 17184
rect 5500 17144 5506 17156
rect 5537 17153 5549 17156
rect 5583 17153 5595 17187
rect 5721 17187 5779 17193
rect 5721 17184 5733 17187
rect 5537 17147 5595 17153
rect 5644 17156 5733 17184
rect 4672 17088 5120 17116
rect 4672 17076 4678 17088
rect 5644 17048 5672 17156
rect 5721 17153 5733 17156
rect 5767 17153 5779 17187
rect 5721 17147 5779 17153
rect 6178 17144 6184 17196
rect 6236 17184 6242 17196
rect 6365 17187 6423 17193
rect 6365 17184 6377 17187
rect 6236 17156 6377 17184
rect 6236 17144 6242 17156
rect 6365 17153 6377 17156
rect 6411 17184 6423 17187
rect 6546 17184 6552 17196
rect 6411 17156 6552 17184
rect 6411 17153 6423 17156
rect 6365 17147 6423 17153
rect 6546 17144 6552 17156
rect 6604 17144 6610 17196
rect 6457 17119 6515 17125
rect 6457 17085 6469 17119
rect 6503 17085 6515 17119
rect 6748 17116 6776 17283
rect 7208 17193 7236 17292
rect 8110 17280 8116 17292
rect 8168 17280 8174 17332
rect 9030 17280 9036 17332
rect 9088 17320 9094 17332
rect 10134 17320 10140 17332
rect 9088 17292 10140 17320
rect 9088 17280 9094 17292
rect 10134 17280 10140 17292
rect 10192 17280 10198 17332
rect 10505 17323 10563 17329
rect 10505 17289 10517 17323
rect 10551 17320 10563 17323
rect 10686 17320 10692 17332
rect 10551 17292 10692 17320
rect 10551 17289 10563 17292
rect 10505 17283 10563 17289
rect 10686 17280 10692 17292
rect 10744 17280 10750 17332
rect 11517 17323 11575 17329
rect 11517 17289 11529 17323
rect 11563 17320 11575 17323
rect 11790 17320 11796 17332
rect 11563 17292 11796 17320
rect 11563 17289 11575 17292
rect 11517 17283 11575 17289
rect 11790 17280 11796 17292
rect 11848 17280 11854 17332
rect 14734 17280 14740 17332
rect 14792 17280 14798 17332
rect 14918 17280 14924 17332
rect 14976 17320 14982 17332
rect 16393 17323 16451 17329
rect 14976 17292 15792 17320
rect 14976 17280 14982 17292
rect 8021 17255 8079 17261
rect 8021 17252 8033 17255
rect 7300 17224 8033 17252
rect 7300 17193 7328 17224
rect 8021 17221 8033 17224
rect 8067 17252 8079 17255
rect 8573 17255 8631 17261
rect 8573 17252 8585 17255
rect 8067 17224 8585 17252
rect 8067 17221 8079 17224
rect 8021 17215 8079 17221
rect 8573 17221 8585 17224
rect 8619 17221 8631 17255
rect 8573 17215 8631 17221
rect 9306 17212 9312 17264
rect 9364 17252 9370 17264
rect 9364 17224 10364 17252
rect 9364 17212 9370 17224
rect 7193 17187 7251 17193
rect 7193 17153 7205 17187
rect 7239 17153 7251 17187
rect 7193 17147 7251 17153
rect 7285 17187 7343 17193
rect 7285 17153 7297 17187
rect 7331 17153 7343 17187
rect 7285 17147 7343 17153
rect 7469 17187 7527 17193
rect 7469 17153 7481 17187
rect 7515 17153 7527 17187
rect 7469 17147 7527 17153
rect 7561 17187 7619 17193
rect 7561 17153 7573 17187
rect 7607 17184 7619 17187
rect 7837 17187 7895 17193
rect 7837 17184 7849 17187
rect 7607 17156 7849 17184
rect 7607 17153 7619 17156
rect 7561 17147 7619 17153
rect 7837 17153 7849 17156
rect 7883 17153 7895 17187
rect 7837 17147 7895 17153
rect 7484 17116 7512 17147
rect 6748 17088 7512 17116
rect 7852 17116 7880 17147
rect 8110 17144 8116 17196
rect 8168 17144 8174 17196
rect 8478 17144 8484 17196
rect 8536 17144 8542 17196
rect 8665 17187 8723 17193
rect 8665 17153 8677 17187
rect 8711 17184 8723 17187
rect 9398 17184 9404 17196
rect 8711 17156 9404 17184
rect 8711 17153 8723 17156
rect 8665 17147 8723 17153
rect 9398 17144 9404 17156
rect 9456 17144 9462 17196
rect 10042 17144 10048 17196
rect 10100 17144 10106 17196
rect 10137 17187 10195 17193
rect 10137 17153 10149 17187
rect 10183 17153 10195 17187
rect 10137 17147 10195 17153
rect 9582 17116 9588 17128
rect 7852 17088 9588 17116
rect 6457 17079 6515 17085
rect 2777 17011 2835 17017
rect 3988 17020 5672 17048
rect 3988 16992 4016 17020
rect 5718 17008 5724 17060
rect 5776 17048 5782 17060
rect 6472 17048 6500 17079
rect 9582 17076 9588 17088
rect 9640 17076 9646 17128
rect 10152 17116 10180 17147
rect 9968 17088 10180 17116
rect 6546 17048 6552 17060
rect 5776 17020 6408 17048
rect 6472 17020 6552 17048
rect 5776 17008 5782 17020
rect 6380 16992 6408 17020
rect 6546 17008 6552 17020
rect 6604 17008 6610 17060
rect 9968 16992 9996 17088
rect 10226 17076 10232 17128
rect 10284 17076 10290 17128
rect 2406 16980 2412 16992
rect 1412 16952 2412 16980
rect 2406 16940 2412 16952
rect 2464 16940 2470 16992
rect 2866 16940 2872 16992
rect 2924 16940 2930 16992
rect 3602 16940 3608 16992
rect 3660 16940 3666 16992
rect 3970 16940 3976 16992
rect 4028 16940 4034 16992
rect 4062 16940 4068 16992
rect 4120 16980 4126 16992
rect 4433 16983 4491 16989
rect 4433 16980 4445 16983
rect 4120 16952 4445 16980
rect 4120 16940 4126 16952
rect 4433 16949 4445 16952
rect 4479 16949 4491 16983
rect 4433 16943 4491 16949
rect 5442 16940 5448 16992
rect 5500 16940 5506 16992
rect 5629 16983 5687 16989
rect 5629 16949 5641 16983
rect 5675 16980 5687 16983
rect 5810 16980 5816 16992
rect 5675 16952 5816 16980
rect 5675 16949 5687 16952
rect 5629 16943 5687 16949
rect 5810 16940 5816 16952
rect 5868 16940 5874 16992
rect 6362 16940 6368 16992
rect 6420 16940 6426 16992
rect 6454 16940 6460 16992
rect 6512 16980 6518 16992
rect 7009 16983 7067 16989
rect 7009 16980 7021 16983
rect 6512 16952 7021 16980
rect 6512 16940 6518 16952
rect 7009 16949 7021 16952
rect 7055 16949 7067 16983
rect 7009 16943 7067 16949
rect 7650 16940 7656 16992
rect 7708 16940 7714 16992
rect 9950 16940 9956 16992
rect 10008 16940 10014 16992
rect 10226 16940 10232 16992
rect 10284 16940 10290 16992
rect 10336 16980 10364 17224
rect 11330 17212 11336 17264
rect 11388 17252 11394 17264
rect 11885 17255 11943 17261
rect 11885 17252 11897 17255
rect 11388 17224 11897 17252
rect 11388 17212 11394 17224
rect 11885 17221 11897 17224
rect 11931 17221 11943 17255
rect 15473 17255 15531 17261
rect 15473 17252 15485 17255
rect 11885 17215 11943 17221
rect 14936 17224 15485 17252
rect 11146 17144 11152 17196
rect 11204 17184 11210 17196
rect 11701 17187 11759 17193
rect 11701 17184 11713 17187
rect 11204 17156 11713 17184
rect 11204 17144 11210 17156
rect 11701 17153 11713 17156
rect 11747 17153 11759 17187
rect 11701 17147 11759 17153
rect 11793 17187 11851 17193
rect 11793 17153 11805 17187
rect 11839 17153 11851 17187
rect 11793 17147 11851 17153
rect 13653 17187 13711 17193
rect 13653 17153 13665 17187
rect 13699 17184 13711 17187
rect 13814 17184 13820 17196
rect 13699 17156 13820 17184
rect 13699 17153 13711 17156
rect 13653 17147 13711 17153
rect 11808 17116 11836 17147
rect 13814 17144 13820 17156
rect 13872 17144 13878 17196
rect 14936 17193 14964 17224
rect 15473 17221 15485 17224
rect 15519 17221 15531 17255
rect 15764 17252 15792 17292
rect 16393 17289 16405 17323
rect 16439 17320 16451 17323
rect 17402 17320 17408 17332
rect 16439 17292 17408 17320
rect 16439 17289 16451 17292
rect 16393 17283 16451 17289
rect 17402 17280 17408 17292
rect 17460 17280 17466 17332
rect 17586 17280 17592 17332
rect 17644 17280 17650 17332
rect 17865 17323 17923 17329
rect 17865 17289 17877 17323
rect 17911 17289 17923 17323
rect 17865 17283 17923 17289
rect 15764 17224 15884 17252
rect 15473 17215 15531 17221
rect 14921 17187 14979 17193
rect 14921 17153 14933 17187
rect 14967 17153 14979 17187
rect 14921 17147 14979 17153
rect 15013 17187 15071 17193
rect 15013 17153 15025 17187
rect 15059 17153 15071 17187
rect 15013 17147 15071 17153
rect 11808 17088 12572 17116
rect 11606 17008 11612 17060
rect 11664 17048 11670 17060
rect 12066 17048 12072 17060
rect 11664 17020 12072 17048
rect 11664 17008 11670 17020
rect 12066 17008 12072 17020
rect 12124 17008 12130 17060
rect 12434 16980 12440 16992
rect 10336 16952 12440 16980
rect 12434 16940 12440 16952
rect 12492 16940 12498 16992
rect 12544 16989 12572 17088
rect 13906 17076 13912 17128
rect 13964 17076 13970 17128
rect 15028 17116 15056 17147
rect 15102 17144 15108 17196
rect 15160 17144 15166 17196
rect 15243 17187 15301 17193
rect 15243 17153 15255 17187
rect 15289 17184 15301 17187
rect 15654 17184 15660 17196
rect 15289 17156 15660 17184
rect 15289 17153 15301 17156
rect 15243 17147 15301 17153
rect 15654 17144 15660 17156
rect 15712 17144 15718 17196
rect 15746 17144 15752 17196
rect 15804 17144 15810 17196
rect 15856 17193 15884 17224
rect 16666 17212 16672 17264
rect 16724 17212 16730 17264
rect 17126 17212 17132 17264
rect 17184 17252 17190 17264
rect 17604 17252 17632 17280
rect 17880 17252 17908 17283
rect 18046 17280 18052 17332
rect 18104 17320 18110 17332
rect 19337 17323 19395 17329
rect 19337 17320 19349 17323
rect 18104 17292 19349 17320
rect 18104 17280 18110 17292
rect 19337 17289 19349 17292
rect 19383 17289 19395 17323
rect 19337 17283 19395 17289
rect 20806 17280 20812 17332
rect 20864 17320 20870 17332
rect 21177 17323 21235 17329
rect 21177 17320 21189 17323
rect 20864 17292 21189 17320
rect 20864 17280 20870 17292
rect 21177 17289 21189 17292
rect 21223 17289 21235 17323
rect 21177 17283 21235 17289
rect 21818 17280 21824 17332
rect 21876 17280 21882 17332
rect 22005 17323 22063 17329
rect 22005 17289 22017 17323
rect 22051 17320 22063 17323
rect 22186 17320 22192 17332
rect 22051 17292 22192 17320
rect 22051 17289 22063 17292
rect 22005 17283 22063 17289
rect 22186 17280 22192 17292
rect 22244 17280 22250 17332
rect 22278 17280 22284 17332
rect 22336 17320 22342 17332
rect 22336 17292 22508 17320
rect 22336 17280 22342 17292
rect 18202 17255 18260 17261
rect 18202 17252 18214 17255
rect 17184 17224 17448 17252
rect 17604 17224 17724 17252
rect 17880 17224 18214 17252
rect 17184 17212 17190 17224
rect 15841 17187 15899 17193
rect 15841 17153 15853 17187
rect 15887 17153 15899 17187
rect 15841 17147 15899 17153
rect 16022 17144 16028 17196
rect 16080 17144 16086 17196
rect 16298 17144 16304 17196
rect 16356 17144 16362 17196
rect 16485 17187 16543 17193
rect 16485 17153 16497 17187
rect 16531 17182 16543 17187
rect 16853 17187 16911 17193
rect 16853 17184 16865 17187
rect 16592 17182 16865 17184
rect 16531 17156 16865 17182
rect 16531 17154 16620 17156
rect 16531 17153 16543 17154
rect 16485 17147 16543 17153
rect 16853 17153 16865 17156
rect 16899 17153 16911 17187
rect 16853 17147 16911 17153
rect 17313 17187 17371 17193
rect 17313 17153 17325 17187
rect 17359 17153 17371 17187
rect 17420 17190 17448 17224
rect 17494 17190 17500 17196
rect 17420 17162 17500 17190
rect 17313 17147 17371 17153
rect 15028 17088 15148 17116
rect 15120 17048 15148 17088
rect 15378 17076 15384 17128
rect 15436 17076 15442 17128
rect 15473 17119 15531 17125
rect 15473 17085 15485 17119
rect 15519 17116 15531 17119
rect 15562 17116 15568 17128
rect 15519 17088 15568 17116
rect 15519 17085 15531 17088
rect 15473 17079 15531 17085
rect 15562 17076 15568 17088
rect 15620 17076 15626 17128
rect 15764 17116 15792 17144
rect 16500 17116 16528 17147
rect 15764 17088 16528 17116
rect 17037 17119 17095 17125
rect 17037 17085 17049 17119
rect 17083 17085 17095 17119
rect 17037 17079 17095 17085
rect 15120 17020 15976 17048
rect 12529 16983 12587 16989
rect 12529 16949 12541 16983
rect 12575 16980 12587 16983
rect 12802 16980 12808 16992
rect 12575 16952 12808 16980
rect 12575 16949 12587 16952
rect 12529 16943 12587 16949
rect 12802 16940 12808 16952
rect 12860 16940 12866 16992
rect 15657 16983 15715 16989
rect 15657 16949 15669 16983
rect 15703 16980 15715 16983
rect 15841 16983 15899 16989
rect 15841 16980 15853 16983
rect 15703 16952 15853 16980
rect 15703 16949 15715 16952
rect 15657 16943 15715 16949
rect 15841 16949 15853 16952
rect 15887 16949 15899 16983
rect 15948 16980 15976 17020
rect 16298 17008 16304 17060
rect 16356 17048 16362 17060
rect 17052 17048 17080 17079
rect 16356 17020 17080 17048
rect 17328 17048 17356 17147
rect 17494 17144 17500 17162
rect 17552 17144 17558 17196
rect 17696 17193 17724 17224
rect 18202 17221 18214 17224
rect 18248 17221 18260 17255
rect 21545 17255 21603 17261
rect 18202 17215 18260 17221
rect 20456 17224 21404 17252
rect 20456 17196 20484 17224
rect 17589 17187 17647 17193
rect 17589 17153 17601 17187
rect 17635 17153 17647 17187
rect 17589 17147 17647 17153
rect 17681 17187 17739 17193
rect 17681 17153 17693 17187
rect 17727 17184 17739 17187
rect 17862 17184 17868 17196
rect 17727 17156 17868 17184
rect 17727 17153 17739 17156
rect 17681 17147 17739 17153
rect 17600 17116 17628 17147
rect 17862 17144 17868 17156
rect 17920 17144 17926 17196
rect 17954 17144 17960 17196
rect 18012 17144 18018 17196
rect 18046 17144 18052 17196
rect 18104 17144 18110 17196
rect 20438 17144 20444 17196
rect 20496 17144 20502 17196
rect 20599 17187 20657 17193
rect 20599 17153 20611 17187
rect 20645 17184 20657 17187
rect 20645 17153 20668 17184
rect 20599 17147 20668 17153
rect 18064 17116 18092 17144
rect 17600 17088 18092 17116
rect 17954 17048 17960 17060
rect 17328 17020 17960 17048
rect 16356 17008 16362 17020
rect 17954 17008 17960 17020
rect 18012 17008 18018 17060
rect 19426 16980 19432 16992
rect 15948 16952 19432 16980
rect 15841 16943 15899 16949
rect 19426 16940 19432 16952
rect 19484 16940 19490 16992
rect 20640 16980 20668 17147
rect 20714 17144 20720 17196
rect 20772 17144 20778 17196
rect 20809 17187 20867 17193
rect 20809 17153 20821 17187
rect 20855 17153 20867 17187
rect 20809 17147 20867 17153
rect 20824 17116 20852 17147
rect 20898 17144 20904 17196
rect 20956 17144 20962 17196
rect 21174 17144 21180 17196
rect 21232 17144 21238 17196
rect 21376 17193 21404 17224
rect 21545 17221 21557 17255
rect 21591 17252 21603 17255
rect 22480 17252 22508 17292
rect 22830 17280 22836 17332
rect 22888 17320 22894 17332
rect 22925 17323 22983 17329
rect 22925 17320 22937 17323
rect 22888 17292 22937 17320
rect 22888 17280 22894 17292
rect 22925 17289 22937 17292
rect 22971 17289 22983 17323
rect 22925 17283 22983 17289
rect 23198 17280 23204 17332
rect 23256 17280 23262 17332
rect 23308 17292 23612 17320
rect 23308 17252 23336 17292
rect 23584 17261 23612 17292
rect 24946 17280 24952 17332
rect 25004 17320 25010 17332
rect 25041 17323 25099 17329
rect 25041 17320 25053 17323
rect 25004 17292 25053 17320
rect 25004 17280 25010 17292
rect 25041 17289 25053 17292
rect 25087 17289 25099 17323
rect 25041 17283 25099 17289
rect 25209 17323 25267 17329
rect 25209 17289 25221 17323
rect 25255 17320 25267 17323
rect 25314 17320 25320 17332
rect 25255 17292 25320 17320
rect 25255 17289 25267 17292
rect 25209 17283 25267 17289
rect 25314 17280 25320 17292
rect 25372 17320 25378 17332
rect 26418 17320 26424 17332
rect 25372 17292 26424 17320
rect 25372 17280 25378 17292
rect 26418 17280 26424 17292
rect 26476 17280 26482 17332
rect 21591 17224 22416 17252
rect 21591 17221 21603 17224
rect 21545 17215 21603 17221
rect 22388 17196 22416 17224
rect 22480 17224 23336 17252
rect 23369 17255 23427 17261
rect 21361 17187 21419 17193
rect 21361 17153 21373 17187
rect 21407 17153 21419 17187
rect 21361 17147 21419 17153
rect 21453 17187 21511 17193
rect 21453 17153 21465 17187
rect 21499 17153 21511 17187
rect 21453 17147 21511 17153
rect 20990 17116 20996 17128
rect 20824 17088 20996 17116
rect 20990 17076 20996 17088
rect 21048 17116 21054 17128
rect 21468 17116 21496 17147
rect 21634 17144 21640 17196
rect 21692 17144 21698 17196
rect 22002 17187 22060 17193
rect 22002 17153 22014 17187
rect 22048 17153 22060 17187
rect 22002 17147 22060 17153
rect 21048 17088 21496 17116
rect 22017 17116 22045 17147
rect 22370 17144 22376 17196
rect 22428 17144 22434 17196
rect 22480 17193 22508 17224
rect 23369 17221 23381 17255
rect 23415 17252 23427 17255
rect 23569 17255 23627 17261
rect 23415 17224 23520 17252
rect 23415 17221 23427 17224
rect 23369 17215 23427 17221
rect 22465 17187 22523 17193
rect 22465 17153 22477 17187
rect 22511 17184 22523 17187
rect 22557 17187 22615 17193
rect 22557 17184 22569 17187
rect 22511 17156 22569 17184
rect 22511 17153 22523 17156
rect 22465 17147 22523 17153
rect 22557 17153 22569 17156
rect 22603 17153 22615 17187
rect 22557 17147 22615 17153
rect 22925 17187 22983 17193
rect 22925 17153 22937 17187
rect 22971 17184 22983 17187
rect 23492 17184 23520 17224
rect 23569 17221 23581 17255
rect 23615 17221 23627 17255
rect 23569 17215 23627 17221
rect 25409 17255 25467 17261
rect 25409 17221 25421 17255
rect 25455 17221 25467 17255
rect 25409 17215 25467 17221
rect 23658 17184 23664 17196
rect 22971 17156 23060 17184
rect 22971 17153 22983 17156
rect 22925 17147 22983 17153
rect 23032 17116 23060 17156
rect 23492 17156 23664 17184
rect 22017 17088 23060 17116
rect 21048 17076 21054 17088
rect 21085 17051 21143 17057
rect 21085 17017 21097 17051
rect 21131 17048 21143 17051
rect 23032 17048 23060 17088
rect 23109 17119 23167 17125
rect 23109 17085 23121 17119
rect 23155 17116 23167 17119
rect 23492 17116 23520 17156
rect 23658 17144 23664 17156
rect 23716 17144 23722 17196
rect 24578 17144 24584 17196
rect 24636 17184 24642 17196
rect 24765 17187 24823 17193
rect 24765 17184 24777 17187
rect 24636 17156 24777 17184
rect 24636 17144 24642 17156
rect 24765 17153 24777 17156
rect 24811 17153 24823 17187
rect 24765 17147 24823 17153
rect 24854 17144 24860 17196
rect 24912 17184 24918 17196
rect 24949 17187 25007 17193
rect 24949 17184 24961 17187
rect 24912 17156 24961 17184
rect 24912 17144 24918 17156
rect 24949 17153 24961 17156
rect 24995 17153 25007 17187
rect 25424 17184 25452 17215
rect 25498 17184 25504 17196
rect 25424 17156 25504 17184
rect 24949 17147 25007 17153
rect 25498 17144 25504 17156
rect 25556 17144 25562 17196
rect 25685 17187 25743 17193
rect 25685 17153 25697 17187
rect 25731 17153 25743 17187
rect 25685 17147 25743 17153
rect 23155 17088 23520 17116
rect 23155 17085 23167 17088
rect 23109 17079 23167 17085
rect 24857 17051 24915 17057
rect 21131 17020 22094 17048
rect 23032 17020 23428 17048
rect 21131 17017 21143 17020
rect 21085 17011 21143 17017
rect 21174 16980 21180 16992
rect 20640 16952 21180 16980
rect 21174 16940 21180 16952
rect 21232 16940 21238 16992
rect 22066 16980 22094 17020
rect 23400 16992 23428 17020
rect 24857 17017 24869 17051
rect 24903 17048 24915 17051
rect 25700 17048 25728 17147
rect 25774 17144 25780 17196
rect 25832 17144 25838 17196
rect 25866 17144 25872 17196
rect 25924 17184 25930 17196
rect 26053 17187 26111 17193
rect 26053 17184 26065 17187
rect 25924 17156 26065 17184
rect 25924 17144 25930 17156
rect 26053 17153 26065 17156
rect 26099 17153 26111 17187
rect 26053 17147 26111 17153
rect 24903 17020 25728 17048
rect 25792 17048 25820 17144
rect 25869 17051 25927 17057
rect 25869 17048 25881 17051
rect 25792 17020 25881 17048
rect 24903 17017 24915 17020
rect 24857 17011 24915 17017
rect 22830 16980 22836 16992
rect 22066 16952 22836 16980
rect 22830 16940 22836 16952
rect 22888 16940 22894 16992
rect 23382 16940 23388 16992
rect 23440 16940 23446 16992
rect 25240 16989 25268 17020
rect 25869 17017 25881 17020
rect 25915 17017 25927 17051
rect 25869 17011 25927 17017
rect 25225 16983 25283 16989
rect 25225 16949 25237 16983
rect 25271 16949 25283 16983
rect 25225 16943 25283 16949
rect 25501 16983 25559 16989
rect 25501 16949 25513 16983
rect 25547 16980 25559 16983
rect 25590 16980 25596 16992
rect 25547 16952 25596 16980
rect 25547 16949 25559 16952
rect 25501 16943 25559 16949
rect 25590 16940 25596 16952
rect 25648 16940 25654 16992
rect 1104 16890 27876 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 27876 16890
rect 1104 16816 27876 16838
rect 1946 16736 1952 16788
rect 2004 16736 2010 16788
rect 4798 16776 4804 16788
rect 3988 16748 4804 16776
rect 2590 16668 2596 16720
rect 2648 16708 2654 16720
rect 2866 16708 2872 16720
rect 2648 16680 2872 16708
rect 2648 16668 2654 16680
rect 2866 16668 2872 16680
rect 2924 16668 2930 16720
rect 2958 16668 2964 16720
rect 3016 16668 3022 16720
rect 2976 16640 3004 16668
rect 2332 16612 2728 16640
rect 2133 16575 2191 16581
rect 2133 16541 2145 16575
rect 2179 16572 2191 16575
rect 2332 16572 2360 16612
rect 2179 16544 2360 16572
rect 2179 16541 2191 16544
rect 2133 16535 2191 16541
rect 2590 16532 2596 16584
rect 2648 16532 2654 16584
rect 2700 16572 2728 16612
rect 2884 16612 3004 16640
rect 3329 16643 3387 16649
rect 2884 16581 2912 16612
rect 3329 16609 3341 16643
rect 3375 16640 3387 16643
rect 3988 16640 4016 16748
rect 4798 16736 4804 16748
rect 4856 16736 4862 16788
rect 6362 16736 6368 16788
rect 6420 16776 6426 16788
rect 6549 16779 6607 16785
rect 6549 16776 6561 16779
rect 6420 16748 6561 16776
rect 6420 16736 6426 16748
rect 6549 16745 6561 16748
rect 6595 16745 6607 16779
rect 6549 16739 6607 16745
rect 9582 16736 9588 16788
rect 9640 16736 9646 16788
rect 10042 16736 10048 16788
rect 10100 16776 10106 16788
rect 10594 16776 10600 16788
rect 10100 16748 10600 16776
rect 10100 16736 10106 16748
rect 10594 16736 10600 16748
rect 10652 16736 10658 16788
rect 11054 16736 11060 16788
rect 11112 16736 11118 16788
rect 12161 16779 12219 16785
rect 12161 16745 12173 16779
rect 12207 16776 12219 16779
rect 13078 16776 13084 16788
rect 12207 16748 13084 16776
rect 12207 16745 12219 16748
rect 12161 16739 12219 16745
rect 13078 16736 13084 16748
rect 13136 16736 13142 16788
rect 13906 16736 13912 16788
rect 13964 16776 13970 16788
rect 15470 16776 15476 16788
rect 13964 16748 15476 16776
rect 13964 16736 13970 16748
rect 4430 16668 4436 16720
rect 4488 16708 4494 16720
rect 5258 16708 5264 16720
rect 4488 16680 5264 16708
rect 4488 16668 4494 16680
rect 5258 16668 5264 16680
rect 5316 16668 5322 16720
rect 8570 16668 8576 16720
rect 8628 16708 8634 16720
rect 9490 16708 9496 16720
rect 8628 16680 9496 16708
rect 8628 16668 8634 16680
rect 9490 16668 9496 16680
rect 9548 16708 9554 16720
rect 10413 16711 10471 16717
rect 10413 16708 10425 16711
rect 9548 16680 10425 16708
rect 9548 16668 9554 16680
rect 5442 16640 5448 16652
rect 3375 16612 4016 16640
rect 4080 16612 5448 16640
rect 3375 16609 3387 16612
rect 3329 16603 3387 16609
rect 2777 16575 2835 16581
rect 2777 16572 2789 16575
rect 2700 16544 2789 16572
rect 2777 16541 2789 16544
rect 2823 16541 2835 16575
rect 2777 16535 2835 16541
rect 2869 16575 2927 16581
rect 2869 16541 2881 16575
rect 2915 16541 2927 16575
rect 2869 16535 2927 16541
rect 3145 16575 3203 16581
rect 3145 16541 3157 16575
rect 3191 16572 3203 16575
rect 3878 16572 3884 16584
rect 3191 16544 3884 16572
rect 3191 16541 3203 16544
rect 3145 16535 3203 16541
rect 3878 16532 3884 16544
rect 3936 16532 3942 16584
rect 3970 16532 3976 16584
rect 4028 16532 4034 16584
rect 4080 16581 4108 16612
rect 5442 16600 5448 16612
rect 5500 16600 5506 16652
rect 6641 16643 6699 16649
rect 6641 16640 6653 16643
rect 5828 16612 6653 16640
rect 5828 16584 5856 16612
rect 6641 16609 6653 16612
rect 6687 16609 6699 16643
rect 6641 16603 6699 16609
rect 9033 16643 9091 16649
rect 9033 16609 9045 16643
rect 9079 16640 9091 16643
rect 9769 16643 9827 16649
rect 9079 16612 9444 16640
rect 9079 16609 9091 16612
rect 9033 16603 9091 16609
rect 9416 16584 9444 16612
rect 9769 16609 9781 16643
rect 9815 16640 9827 16643
rect 9950 16640 9956 16652
rect 9815 16612 9956 16640
rect 9815 16609 9827 16612
rect 9769 16603 9827 16609
rect 9950 16600 9956 16612
rect 10008 16600 10014 16652
rect 10244 16649 10272 16680
rect 10413 16677 10425 16680
rect 10459 16677 10471 16711
rect 10612 16708 10640 16736
rect 12345 16711 12403 16717
rect 10612 16680 12020 16708
rect 10413 16671 10471 16677
rect 11992 16652 12020 16680
rect 12345 16677 12357 16711
rect 12391 16708 12403 16711
rect 12391 16680 12480 16708
rect 12391 16677 12403 16680
rect 12345 16671 12403 16677
rect 10229 16643 10287 16649
rect 10229 16609 10241 16643
rect 10275 16609 10287 16643
rect 10229 16603 10287 16609
rect 11514 16600 11520 16652
rect 11572 16640 11578 16652
rect 11609 16643 11667 16649
rect 11609 16640 11621 16643
rect 11572 16612 11621 16640
rect 11572 16600 11578 16612
rect 11609 16609 11621 16612
rect 11655 16609 11667 16643
rect 11609 16603 11667 16609
rect 11974 16600 11980 16652
rect 12032 16600 12038 16652
rect 4065 16575 4123 16581
rect 4065 16541 4077 16575
rect 4111 16541 4123 16575
rect 4065 16535 4123 16541
rect 4430 16532 4436 16584
rect 4488 16532 4494 16584
rect 4614 16532 4620 16584
rect 4672 16532 4678 16584
rect 5810 16532 5816 16584
rect 5868 16532 5874 16584
rect 5905 16575 5963 16581
rect 5905 16541 5917 16575
rect 5951 16572 5963 16575
rect 5994 16572 6000 16584
rect 5951 16544 6000 16572
rect 5951 16541 5963 16544
rect 5905 16535 5963 16541
rect 5994 16532 6000 16544
rect 6052 16572 6058 16584
rect 6454 16572 6460 16584
rect 6052 16544 6460 16572
rect 6052 16532 6058 16544
rect 6454 16532 6460 16544
rect 6512 16532 6518 16584
rect 6546 16532 6552 16584
rect 6604 16532 6610 16584
rect 6822 16532 6828 16584
rect 6880 16572 6886 16584
rect 7650 16572 7656 16584
rect 6880 16544 7656 16572
rect 6880 16532 6886 16544
rect 7650 16532 7656 16544
rect 7708 16532 7714 16584
rect 8846 16532 8852 16584
rect 8904 16572 8910 16584
rect 8941 16575 8999 16581
rect 8941 16572 8953 16575
rect 8904 16544 8953 16572
rect 8904 16532 8910 16544
rect 8941 16541 8953 16544
rect 8987 16541 8999 16575
rect 8941 16535 8999 16541
rect 9125 16575 9183 16581
rect 9125 16541 9137 16575
rect 9171 16541 9183 16575
rect 9125 16535 9183 16541
rect 2225 16507 2283 16513
rect 2225 16473 2237 16507
rect 2271 16473 2283 16507
rect 2225 16467 2283 16473
rect 2240 16436 2268 16467
rect 2314 16464 2320 16516
rect 2372 16464 2378 16516
rect 2498 16513 2504 16516
rect 2455 16507 2504 16513
rect 2455 16473 2467 16507
rect 2501 16473 2504 16507
rect 2455 16467 2504 16473
rect 2498 16464 2504 16467
rect 2556 16464 2562 16516
rect 3602 16504 3608 16516
rect 2746 16476 3608 16504
rect 2746 16436 2774 16476
rect 3602 16464 3608 16476
rect 3660 16464 3666 16516
rect 6178 16464 6184 16516
rect 6236 16464 6242 16516
rect 6273 16507 6331 16513
rect 6273 16473 6285 16507
rect 6319 16473 6331 16507
rect 9140 16504 9168 16535
rect 9398 16532 9404 16584
rect 9456 16572 9462 16584
rect 9861 16575 9919 16581
rect 9861 16572 9873 16575
rect 9456 16544 9873 16572
rect 9456 16532 9462 16544
rect 9861 16541 9873 16544
rect 9907 16541 9919 16575
rect 9861 16535 9919 16541
rect 10597 16575 10655 16581
rect 10597 16541 10609 16575
rect 10643 16572 10655 16575
rect 11425 16575 11483 16581
rect 11425 16572 11437 16575
rect 10643 16544 11437 16572
rect 10643 16541 10655 16544
rect 10597 16535 10655 16541
rect 11425 16541 11437 16544
rect 11471 16572 11483 16575
rect 11882 16572 11888 16584
rect 11471 16544 11888 16572
rect 11471 16541 11483 16544
rect 11425 16535 11483 16541
rect 11882 16532 11888 16544
rect 11940 16532 11946 16584
rect 12158 16532 12164 16584
rect 12216 16532 12222 16584
rect 12452 16581 12480 16680
rect 13446 16600 13452 16652
rect 13504 16640 13510 16652
rect 14274 16640 14280 16652
rect 13504 16612 14280 16640
rect 13504 16600 13510 16612
rect 14274 16600 14280 16612
rect 14332 16600 14338 16652
rect 14476 16649 14504 16748
rect 15470 16736 15476 16748
rect 15528 16736 15534 16788
rect 17954 16736 17960 16788
rect 18012 16776 18018 16788
rect 18049 16779 18107 16785
rect 18049 16776 18061 16779
rect 18012 16748 18061 16776
rect 18012 16736 18018 16748
rect 18049 16745 18061 16748
rect 18095 16745 18107 16779
rect 18049 16739 18107 16745
rect 19978 16736 19984 16788
rect 20036 16776 20042 16788
rect 20073 16779 20131 16785
rect 20073 16776 20085 16779
rect 20036 16748 20085 16776
rect 20036 16736 20042 16748
rect 20073 16745 20085 16748
rect 20119 16745 20131 16779
rect 20073 16739 20131 16745
rect 20438 16736 20444 16788
rect 20496 16776 20502 16788
rect 20533 16779 20591 16785
rect 20533 16776 20545 16779
rect 20496 16748 20545 16776
rect 20496 16736 20502 16748
rect 20533 16745 20545 16748
rect 20579 16745 20591 16779
rect 20533 16739 20591 16745
rect 20990 16736 20996 16788
rect 21048 16736 21054 16788
rect 21082 16736 21088 16788
rect 21140 16776 21146 16788
rect 21177 16779 21235 16785
rect 21177 16776 21189 16779
rect 21140 16748 21189 16776
rect 21140 16736 21146 16748
rect 21177 16745 21189 16748
rect 21223 16745 21235 16779
rect 21177 16739 21235 16745
rect 23385 16779 23443 16785
rect 23385 16745 23397 16779
rect 23431 16776 23443 16779
rect 23566 16776 23572 16788
rect 23431 16748 23572 16776
rect 23431 16745 23443 16748
rect 23385 16739 23443 16745
rect 23566 16736 23572 16748
rect 23624 16736 23630 16788
rect 17126 16668 17132 16720
rect 17184 16708 17190 16720
rect 19889 16711 19947 16717
rect 17184 16680 18736 16708
rect 17184 16668 17190 16680
rect 14461 16643 14519 16649
rect 14461 16609 14473 16643
rect 14507 16609 14519 16643
rect 14461 16603 14519 16609
rect 17218 16600 17224 16652
rect 17276 16600 17282 16652
rect 18708 16649 18736 16680
rect 19889 16677 19901 16711
rect 19935 16708 19947 16711
rect 19935 16680 20852 16708
rect 19935 16677 19947 16680
rect 19889 16671 19947 16677
rect 17681 16643 17739 16649
rect 17681 16609 17693 16643
rect 17727 16640 17739 16643
rect 18509 16643 18567 16649
rect 18509 16640 18521 16643
rect 17727 16612 18521 16640
rect 17727 16609 17739 16612
rect 17681 16603 17739 16609
rect 18509 16609 18521 16612
rect 18555 16609 18567 16643
rect 18509 16603 18567 16609
rect 18693 16643 18751 16649
rect 18693 16609 18705 16643
rect 18739 16640 18751 16643
rect 19150 16640 19156 16652
rect 18739 16612 19156 16640
rect 18739 16609 18751 16612
rect 18693 16603 18751 16609
rect 19150 16600 19156 16612
rect 19208 16600 19214 16652
rect 19659 16643 19717 16649
rect 19659 16609 19671 16643
rect 19705 16640 19717 16643
rect 20257 16643 20315 16649
rect 20257 16640 20269 16643
rect 19705 16612 20269 16640
rect 19705 16609 19717 16612
rect 19659 16603 19717 16609
rect 20257 16609 20269 16612
rect 20303 16640 20315 16643
rect 20714 16640 20720 16652
rect 20303 16612 20720 16640
rect 20303 16609 20315 16612
rect 20257 16603 20315 16609
rect 20714 16600 20720 16612
rect 20772 16600 20778 16652
rect 20824 16640 20852 16680
rect 20898 16668 20904 16720
rect 20956 16708 20962 16720
rect 21545 16711 21603 16717
rect 21545 16708 21557 16711
rect 20956 16680 21557 16708
rect 20956 16668 20962 16680
rect 21545 16677 21557 16680
rect 21591 16708 21603 16711
rect 21634 16708 21640 16720
rect 21591 16680 21640 16708
rect 21591 16677 21603 16680
rect 21545 16671 21603 16677
rect 21634 16668 21640 16680
rect 21692 16668 21698 16720
rect 21174 16640 21180 16652
rect 20824 16612 21180 16640
rect 21174 16600 21180 16612
rect 21232 16600 21238 16652
rect 21269 16643 21327 16649
rect 21269 16609 21281 16643
rect 21315 16640 21327 16643
rect 21453 16643 21511 16649
rect 21453 16640 21465 16643
rect 21315 16612 21465 16640
rect 21315 16609 21327 16612
rect 21269 16603 21327 16609
rect 21453 16609 21465 16612
rect 21499 16609 21511 16643
rect 21453 16603 21511 16609
rect 23201 16643 23259 16649
rect 23201 16609 23213 16643
rect 23247 16640 23259 16643
rect 23569 16643 23627 16649
rect 23569 16640 23581 16643
rect 23247 16612 23581 16640
rect 23247 16609 23259 16612
rect 23201 16603 23259 16609
rect 23569 16609 23581 16612
rect 23615 16609 23627 16643
rect 23569 16603 23627 16609
rect 12437 16575 12495 16581
rect 12437 16541 12449 16575
rect 12483 16541 12495 16575
rect 12437 16535 12495 16541
rect 12802 16532 12808 16584
rect 12860 16572 12866 16584
rect 12989 16575 13047 16581
rect 12989 16572 13001 16575
rect 12860 16544 13001 16572
rect 12860 16532 12866 16544
rect 12989 16541 13001 16544
rect 13035 16541 13047 16575
rect 12989 16535 13047 16541
rect 14093 16575 14151 16581
rect 14093 16541 14105 16575
rect 14139 16572 14151 16575
rect 14366 16572 14372 16584
rect 14139 16544 14372 16572
rect 14139 16541 14151 16544
rect 14093 16535 14151 16541
rect 14366 16532 14372 16544
rect 14424 16532 14430 16584
rect 15562 16532 15568 16584
rect 15620 16572 15626 16584
rect 17313 16575 17371 16581
rect 17313 16572 17325 16575
rect 15620 16544 17325 16572
rect 15620 16532 15626 16544
rect 17313 16541 17325 16544
rect 17359 16572 17371 16575
rect 18046 16572 18052 16584
rect 17359 16544 18052 16572
rect 17359 16541 17371 16544
rect 17313 16535 17371 16541
rect 18046 16532 18052 16544
rect 18104 16532 18110 16584
rect 19521 16575 19579 16581
rect 19521 16541 19533 16575
rect 19567 16572 19579 16575
rect 19797 16575 19855 16581
rect 19567 16544 19748 16572
rect 19567 16541 19579 16544
rect 19521 16535 19579 16541
rect 19720 16516 19748 16544
rect 19797 16541 19809 16575
rect 19843 16541 19855 16575
rect 19797 16535 19855 16541
rect 9674 16504 9680 16516
rect 9140 16476 9680 16504
rect 6273 16467 6331 16473
rect 2240 16408 2774 16436
rect 4246 16396 4252 16448
rect 4304 16396 4310 16448
rect 4522 16396 4528 16448
rect 4580 16396 4586 16448
rect 5626 16396 5632 16448
rect 5684 16396 5690 16448
rect 6288 16436 6316 16467
rect 9674 16464 9680 16476
rect 9732 16504 9738 16516
rect 10137 16507 10195 16513
rect 10137 16504 10149 16507
rect 9732 16476 10149 16504
rect 9732 16464 9738 16476
rect 10137 16473 10149 16476
rect 10183 16473 10195 16507
rect 10137 16467 10195 16473
rect 10686 16464 10692 16516
rect 10744 16504 10750 16516
rect 10781 16507 10839 16513
rect 10781 16504 10793 16507
rect 10744 16476 10793 16504
rect 10744 16464 10750 16476
rect 10781 16473 10793 16476
rect 10827 16473 10839 16507
rect 10781 16467 10839 16473
rect 11241 16507 11299 16513
rect 11241 16473 11253 16507
rect 11287 16504 11299 16507
rect 11287 16476 11560 16504
rect 11287 16473 11299 16476
rect 11241 16467 11299 16473
rect 6365 16439 6423 16445
rect 6365 16436 6377 16439
rect 6288 16408 6377 16436
rect 6365 16405 6377 16408
rect 6411 16405 6423 16439
rect 6365 16399 6423 16405
rect 8938 16396 8944 16448
rect 8996 16436 9002 16448
rect 11333 16439 11391 16445
rect 11333 16436 11345 16439
rect 8996 16408 11345 16436
rect 8996 16396 9002 16408
rect 11333 16405 11345 16408
rect 11379 16405 11391 16439
rect 11532 16436 11560 16476
rect 11698 16464 11704 16516
rect 11756 16464 11762 16516
rect 14734 16513 14740 16516
rect 14728 16467 14740 16513
rect 14734 16464 14740 16467
rect 14792 16464 14798 16516
rect 19702 16464 19708 16516
rect 19760 16464 19766 16516
rect 19812 16504 19840 16535
rect 19978 16532 19984 16584
rect 20036 16532 20042 16584
rect 20346 16532 20352 16584
rect 20404 16572 20410 16584
rect 21284 16572 21312 16603
rect 20404 16544 21312 16572
rect 20404 16532 20410 16544
rect 21358 16532 21364 16584
rect 21416 16532 21422 16584
rect 21637 16575 21695 16581
rect 21637 16541 21649 16575
rect 21683 16541 21695 16575
rect 21637 16535 21695 16541
rect 21729 16575 21787 16581
rect 21729 16541 21741 16575
rect 21775 16572 21787 16575
rect 21910 16572 21916 16584
rect 21775 16544 21916 16572
rect 21775 16541 21787 16544
rect 21729 16535 21787 16541
rect 20073 16507 20131 16513
rect 20073 16504 20085 16507
rect 19812 16476 20085 16504
rect 20073 16473 20085 16476
rect 20119 16504 20131 16507
rect 20254 16504 20260 16516
rect 20119 16476 20260 16504
rect 20119 16473 20131 16476
rect 20073 16467 20131 16473
rect 20254 16464 20260 16476
rect 20312 16504 20318 16516
rect 21652 16504 21680 16535
rect 20312 16476 21680 16504
rect 20312 16464 20318 16476
rect 12529 16439 12587 16445
rect 12529 16436 12541 16439
rect 11532 16408 12541 16436
rect 11333 16399 11391 16405
rect 12529 16405 12541 16408
rect 12575 16405 12587 16439
rect 12529 16399 12587 16405
rect 13262 16396 13268 16448
rect 13320 16436 13326 16448
rect 13633 16439 13691 16445
rect 13633 16436 13645 16439
rect 13320 16408 13645 16436
rect 13320 16396 13326 16408
rect 13633 16405 13645 16408
rect 13679 16405 13691 16439
rect 13633 16399 13691 16405
rect 14274 16396 14280 16448
rect 14332 16396 14338 16448
rect 15654 16396 15660 16448
rect 15712 16436 15718 16448
rect 15841 16439 15899 16445
rect 15841 16436 15853 16439
rect 15712 16408 15853 16436
rect 15712 16396 15718 16408
rect 15841 16405 15853 16408
rect 15887 16405 15899 16439
rect 15841 16399 15899 16405
rect 18417 16439 18475 16445
rect 18417 16405 18429 16439
rect 18463 16436 18475 16439
rect 19242 16436 19248 16448
rect 18463 16408 19248 16436
rect 18463 16405 18475 16408
rect 18417 16399 18475 16405
rect 19242 16396 19248 16408
rect 19300 16396 19306 16448
rect 19720 16436 19748 16464
rect 20346 16436 20352 16448
rect 19720 16408 20352 16436
rect 20346 16396 20352 16408
rect 20404 16396 20410 16448
rect 20714 16396 20720 16448
rect 20772 16436 20778 16448
rect 21744 16436 21772 16535
rect 21910 16532 21916 16544
rect 21968 16532 21974 16584
rect 23106 16532 23112 16584
rect 23164 16532 23170 16584
rect 23753 16575 23811 16581
rect 23753 16541 23765 16575
rect 23799 16541 23811 16575
rect 23753 16535 23811 16541
rect 22830 16464 22836 16516
rect 22888 16504 22894 16516
rect 23768 16504 23796 16535
rect 24026 16532 24032 16584
rect 24084 16532 24090 16584
rect 22888 16476 23796 16504
rect 22888 16464 22894 16476
rect 20772 16408 21772 16436
rect 20772 16396 20778 16408
rect 23382 16396 23388 16448
rect 23440 16436 23446 16448
rect 23937 16439 23995 16445
rect 23937 16436 23949 16439
rect 23440 16408 23949 16436
rect 23440 16396 23446 16408
rect 23937 16405 23949 16408
rect 23983 16436 23995 16439
rect 25130 16436 25136 16448
rect 23983 16408 25136 16436
rect 23983 16405 23995 16408
rect 23937 16399 23995 16405
rect 25130 16396 25136 16408
rect 25188 16396 25194 16448
rect 1104 16346 27876 16368
rect 1104 16294 4874 16346
rect 4926 16294 4938 16346
rect 4990 16294 5002 16346
rect 5054 16294 5066 16346
rect 5118 16294 5130 16346
rect 5182 16294 27876 16346
rect 1104 16272 27876 16294
rect 2314 16192 2320 16244
rect 2372 16232 2378 16244
rect 2498 16232 2504 16244
rect 2372 16204 2504 16232
rect 2372 16192 2378 16204
rect 2498 16192 2504 16204
rect 2556 16232 2562 16244
rect 7834 16232 7840 16244
rect 2556 16204 7840 16232
rect 2556 16192 2562 16204
rect 7834 16192 7840 16204
rect 7892 16192 7898 16244
rect 9953 16235 10011 16241
rect 9953 16201 9965 16235
rect 9999 16201 10011 16235
rect 11698 16232 11704 16244
rect 9953 16195 10011 16201
rect 10244 16204 11704 16232
rect 3970 16124 3976 16176
rect 4028 16164 4034 16176
rect 4028 16136 4476 16164
rect 4028 16124 4034 16136
rect 4246 16056 4252 16108
rect 4304 16056 4310 16108
rect 4448 16105 4476 16136
rect 4798 16124 4804 16176
rect 4856 16164 4862 16176
rect 9968 16164 9996 16195
rect 10244 16176 10272 16204
rect 11698 16192 11704 16204
rect 11756 16192 11762 16244
rect 12526 16192 12532 16244
rect 12584 16192 12590 16244
rect 13173 16235 13231 16241
rect 13173 16201 13185 16235
rect 13219 16232 13231 16235
rect 13219 16204 13759 16232
rect 13219 16201 13231 16204
rect 13173 16195 13231 16201
rect 10226 16164 10232 16176
rect 4856 16136 5304 16164
rect 4856 16124 4862 16136
rect 4433 16099 4491 16105
rect 4433 16065 4445 16099
rect 4479 16065 4491 16099
rect 4433 16059 4491 16065
rect 4522 16056 4528 16108
rect 4580 16096 4586 16108
rect 4706 16096 4712 16108
rect 4580 16068 4712 16096
rect 4580 16056 4586 16068
rect 4706 16056 4712 16068
rect 4764 16096 4770 16108
rect 5276 16105 5304 16136
rect 5828 16136 6224 16164
rect 4893 16099 4951 16105
rect 4893 16096 4905 16099
rect 4764 16068 4905 16096
rect 4764 16056 4770 16068
rect 4893 16065 4905 16068
rect 4939 16065 4951 16099
rect 4893 16059 4951 16065
rect 5261 16099 5319 16105
rect 5261 16065 5273 16099
rect 5307 16065 5319 16099
rect 5261 16059 5319 16065
rect 5718 16056 5724 16108
rect 5776 16096 5782 16108
rect 5828 16105 5856 16136
rect 5813 16099 5871 16105
rect 5813 16096 5825 16099
rect 5776 16068 5825 16096
rect 5776 16056 5782 16068
rect 5813 16065 5825 16068
rect 5859 16065 5871 16099
rect 5813 16059 5871 16065
rect 5902 16056 5908 16108
rect 5960 16096 5966 16108
rect 6196 16105 6224 16136
rect 8128 16136 9996 16164
rect 10060 16136 10232 16164
rect 8128 16108 8156 16136
rect 5997 16099 6055 16105
rect 5997 16096 6009 16099
rect 5960 16068 6009 16096
rect 5960 16056 5966 16068
rect 5997 16065 6009 16068
rect 6043 16065 6055 16099
rect 5997 16059 6055 16065
rect 6181 16099 6239 16105
rect 6181 16065 6193 16099
rect 6227 16096 6239 16099
rect 6822 16096 6828 16108
rect 6227 16068 6828 16096
rect 6227 16065 6239 16068
rect 6181 16059 6239 16065
rect 6822 16056 6828 16068
rect 6880 16056 6886 16108
rect 7469 16099 7527 16105
rect 7469 16065 7481 16099
rect 7515 16065 7527 16099
rect 7469 16059 7527 16065
rect 4264 16028 4292 16056
rect 4614 16028 4620 16040
rect 4264 16000 4620 16028
rect 4614 15988 4620 16000
rect 4672 15988 4678 16040
rect 7484 16028 7512 16059
rect 7650 16056 7656 16108
rect 7708 16056 7714 16108
rect 7742 16056 7748 16108
rect 7800 16056 7806 16108
rect 8021 16099 8079 16105
rect 8021 16065 8033 16099
rect 8067 16096 8079 16099
rect 8110 16096 8116 16108
rect 8067 16068 8116 16096
rect 8067 16065 8079 16068
rect 8021 16059 8079 16065
rect 8110 16056 8116 16068
rect 8168 16056 8174 16108
rect 8205 16099 8263 16105
rect 8205 16065 8217 16099
rect 8251 16096 8263 16099
rect 8386 16096 8392 16108
rect 8251 16068 8392 16096
rect 8251 16065 8263 16068
rect 8205 16059 8263 16065
rect 8386 16056 8392 16068
rect 8444 16056 8450 16108
rect 8478 16056 8484 16108
rect 8536 16096 8542 16108
rect 8956 16105 8984 16136
rect 8665 16099 8723 16105
rect 8665 16096 8677 16099
rect 8536 16068 8677 16096
rect 8536 16056 8542 16068
rect 8665 16065 8677 16068
rect 8711 16096 8723 16099
rect 8757 16099 8815 16105
rect 8757 16096 8769 16099
rect 8711 16068 8769 16096
rect 8711 16065 8723 16068
rect 8665 16059 8723 16065
rect 8757 16065 8769 16068
rect 8803 16065 8815 16099
rect 8757 16059 8815 16065
rect 8941 16099 8999 16105
rect 8941 16065 8953 16099
rect 8987 16065 8999 16099
rect 8941 16059 8999 16065
rect 9950 16056 9956 16108
rect 10008 16096 10014 16108
rect 10060 16096 10088 16136
rect 10226 16124 10232 16136
rect 10284 16124 10290 16176
rect 10321 16167 10379 16173
rect 10321 16133 10333 16167
rect 10367 16164 10379 16167
rect 10778 16164 10784 16176
rect 10367 16136 10784 16164
rect 10367 16133 10379 16136
rect 10321 16127 10379 16133
rect 10778 16124 10784 16136
rect 10836 16124 10842 16176
rect 10870 16124 10876 16176
rect 10928 16124 10934 16176
rect 11054 16124 11060 16176
rect 11112 16164 11118 16176
rect 13446 16173 13452 16176
rect 12161 16167 12219 16173
rect 12161 16164 12173 16167
rect 11112 16136 12173 16164
rect 11112 16124 11118 16136
rect 12161 16133 12173 16136
rect 12207 16133 12219 16167
rect 12161 16127 12219 16133
rect 12377 16167 12435 16173
rect 12377 16133 12389 16167
rect 12423 16164 12435 16167
rect 13423 16167 13452 16173
rect 12423 16136 12940 16164
rect 12423 16133 12435 16136
rect 12377 16127 12435 16133
rect 10008 16068 10088 16096
rect 10132 16099 10190 16105
rect 10008 16056 10014 16068
rect 10132 16065 10144 16099
rect 10178 16065 10190 16099
rect 10132 16059 10190 16065
rect 5460 16000 8524 16028
rect 5460 15972 5488 16000
rect 4065 15963 4123 15969
rect 4065 15929 4077 15963
rect 4111 15960 4123 15963
rect 5442 15960 5448 15972
rect 4111 15932 5448 15960
rect 4111 15929 4123 15932
rect 4065 15923 4123 15929
rect 5442 15920 5448 15932
rect 5500 15920 5506 15972
rect 6178 15852 6184 15904
rect 6236 15852 6242 15904
rect 7190 15852 7196 15904
rect 7248 15892 7254 15904
rect 7285 15895 7343 15901
rect 7285 15892 7297 15895
rect 7248 15864 7297 15892
rect 7248 15852 7254 15864
rect 7285 15861 7297 15864
rect 7331 15861 7343 15895
rect 7285 15855 7343 15861
rect 8021 15895 8079 15901
rect 8021 15861 8033 15895
rect 8067 15892 8079 15895
rect 8110 15892 8116 15904
rect 8067 15864 8116 15892
rect 8067 15861 8079 15864
rect 8021 15855 8079 15861
rect 8110 15852 8116 15864
rect 8168 15852 8174 15904
rect 8294 15852 8300 15904
rect 8352 15852 8358 15904
rect 8496 15901 8524 16000
rect 8570 15988 8576 16040
rect 8628 15988 8634 16040
rect 8846 15988 8852 16040
rect 8904 16028 8910 16040
rect 9125 16031 9183 16037
rect 9125 16028 9137 16031
rect 8904 16000 9137 16028
rect 8904 15988 8910 16000
rect 9125 15997 9137 16000
rect 9171 15997 9183 16031
rect 10147 16028 10175 16059
rect 10410 16056 10416 16108
rect 10468 16105 10474 16108
rect 10468 16099 10507 16105
rect 10495 16065 10507 16099
rect 10468 16059 10507 16065
rect 10468 16056 10474 16059
rect 10594 16056 10600 16108
rect 10652 16056 10658 16108
rect 10686 16056 10692 16108
rect 10744 16096 10750 16108
rect 11793 16099 11851 16105
rect 11793 16096 11805 16099
rect 10744 16068 11805 16096
rect 10744 16056 10750 16068
rect 11793 16065 11805 16068
rect 11839 16065 11851 16099
rect 11793 16059 11851 16065
rect 10147 16000 10492 16028
rect 9125 15991 9183 15997
rect 10464 15960 10492 16000
rect 10689 15963 10747 15969
rect 10689 15960 10701 15963
rect 10464 15932 10701 15960
rect 10689 15929 10701 15932
rect 10735 15929 10747 15963
rect 11241 15963 11299 15969
rect 11241 15960 11253 15963
rect 10689 15923 10747 15929
rect 10796 15932 11253 15960
rect 8481 15895 8539 15901
rect 8481 15861 8493 15895
rect 8527 15892 8539 15895
rect 9858 15892 9864 15904
rect 8527 15864 9864 15892
rect 8527 15861 8539 15864
rect 8481 15855 8539 15861
rect 9858 15852 9864 15864
rect 9916 15852 9922 15904
rect 10410 15852 10416 15904
rect 10468 15892 10474 15904
rect 10594 15892 10600 15904
rect 10468 15864 10600 15892
rect 10468 15852 10474 15864
rect 10594 15852 10600 15864
rect 10652 15892 10658 15904
rect 10796 15892 10824 15932
rect 11241 15929 11253 15932
rect 11287 15960 11299 15963
rect 11330 15960 11336 15972
rect 11287 15932 11336 15960
rect 11287 15929 11299 15932
rect 11241 15923 11299 15929
rect 11330 15920 11336 15932
rect 11388 15920 11394 15972
rect 11808 15960 11836 16059
rect 11882 16056 11888 16108
rect 11940 16096 11946 16108
rect 11977 16099 12035 16105
rect 11977 16096 11989 16099
rect 11940 16068 11989 16096
rect 11940 16056 11946 16068
rect 11977 16065 11989 16068
rect 12023 16065 12035 16099
rect 12802 16096 12808 16108
rect 11977 16059 12035 16065
rect 12406 16068 12808 16096
rect 12406 15960 12434 16068
rect 12802 16056 12808 16068
rect 12860 16056 12866 16108
rect 12912 16040 12940 16136
rect 13423 16133 13435 16167
rect 13423 16127 13452 16133
rect 13446 16124 13452 16127
rect 13504 16124 13510 16176
rect 13731 16164 13759 16204
rect 13814 16192 13820 16244
rect 13872 16232 13878 16244
rect 13909 16235 13967 16241
rect 13909 16232 13921 16235
rect 13872 16204 13921 16232
rect 13872 16192 13878 16204
rect 13909 16201 13921 16204
rect 13955 16201 13967 16235
rect 13909 16195 13967 16201
rect 14918 16192 14924 16244
rect 14976 16232 14982 16244
rect 15013 16235 15071 16241
rect 15013 16232 15025 16235
rect 14976 16204 15025 16232
rect 14976 16192 14982 16204
rect 15013 16201 15025 16204
rect 15059 16201 15071 16235
rect 15013 16195 15071 16201
rect 15194 16192 15200 16244
rect 15252 16192 15258 16244
rect 19150 16192 19156 16244
rect 19208 16232 19214 16244
rect 21818 16232 21824 16244
rect 19208 16204 21824 16232
rect 19208 16192 19214 16204
rect 21818 16192 21824 16204
rect 21876 16192 21882 16244
rect 15381 16167 15439 16173
rect 13731 16136 14044 16164
rect 13262 16056 13268 16108
rect 13320 16056 13326 16108
rect 13538 16056 13544 16108
rect 13596 16056 13602 16108
rect 14016 16105 14044 16136
rect 15381 16133 15393 16167
rect 15427 16164 15439 16167
rect 17678 16164 17684 16176
rect 15427 16136 17684 16164
rect 15427 16133 15439 16136
rect 15381 16127 15439 16133
rect 17678 16124 17684 16136
rect 17736 16124 17742 16176
rect 24946 16124 24952 16176
rect 25004 16164 25010 16176
rect 25222 16164 25228 16176
rect 25004 16136 25228 16164
rect 25004 16124 25010 16136
rect 25222 16124 25228 16136
rect 25280 16164 25286 16176
rect 25280 16136 25360 16164
rect 25280 16124 25286 16136
rect 13633 16099 13691 16105
rect 13633 16065 13645 16099
rect 13679 16065 13691 16099
rect 13633 16059 13691 16065
rect 13725 16099 13783 16105
rect 13725 16065 13737 16099
rect 13771 16094 13783 16099
rect 14001 16099 14059 16105
rect 13771 16066 13860 16094
rect 13771 16065 13783 16066
rect 13725 16059 13783 16065
rect 12894 15988 12900 16040
rect 12952 15988 12958 16040
rect 11808 15932 12434 15960
rect 10652 15864 10824 15892
rect 10873 15895 10931 15901
rect 10652 15852 10658 15864
rect 10873 15861 10885 15895
rect 10919 15892 10931 15895
rect 11146 15892 11152 15904
rect 10919 15864 11152 15892
rect 10919 15861 10931 15864
rect 10873 15855 10931 15861
rect 11146 15852 11152 15864
rect 11204 15852 11210 15904
rect 11790 15852 11796 15904
rect 11848 15852 11854 15904
rect 12360 15901 12388 15932
rect 12345 15895 12403 15901
rect 12345 15861 12357 15895
rect 12391 15861 12403 15895
rect 13648 15892 13676 16059
rect 13832 16058 13860 16066
rect 14001 16065 14013 16099
rect 14047 16065 14059 16099
rect 14001 16059 14059 16065
rect 14185 16099 14243 16105
rect 14185 16065 14197 16099
rect 14231 16096 14243 16099
rect 14274 16096 14280 16108
rect 14231 16068 14280 16096
rect 14231 16065 14243 16068
rect 14185 16059 14243 16065
rect 13832 16030 13952 16058
rect 13924 16028 13952 16030
rect 14093 16031 14151 16037
rect 14093 16028 14105 16031
rect 13924 16000 14105 16028
rect 14093 15997 14105 16000
rect 14139 15997 14151 16031
rect 14093 15991 14151 15997
rect 13722 15920 13728 15972
rect 13780 15960 13786 15972
rect 14200 15960 14228 16059
rect 14274 16056 14280 16068
rect 14332 16056 14338 16108
rect 15102 16056 15108 16108
rect 15160 16096 15166 16108
rect 15838 16096 15844 16108
rect 15160 16068 15844 16096
rect 15160 16056 15166 16068
rect 15838 16056 15844 16068
rect 15896 16056 15902 16108
rect 16850 16056 16856 16108
rect 16908 16056 16914 16108
rect 16945 16099 17003 16105
rect 16945 16065 16957 16099
rect 16991 16096 17003 16099
rect 17218 16096 17224 16108
rect 16991 16068 17224 16096
rect 16991 16065 17003 16068
rect 16945 16059 17003 16065
rect 14829 16031 14887 16037
rect 14829 15997 14841 16031
rect 14875 16028 14887 16031
rect 15010 16028 15016 16040
rect 14875 16000 15016 16028
rect 14875 15997 14887 16000
rect 14829 15991 14887 15997
rect 15010 15988 15016 16000
rect 15068 16028 15074 16040
rect 16960 16028 16988 16059
rect 17218 16056 17224 16068
rect 17276 16056 17282 16108
rect 24578 16056 24584 16108
rect 24636 16096 24642 16108
rect 24765 16099 24823 16105
rect 24765 16096 24777 16099
rect 24636 16068 24777 16096
rect 24636 16056 24642 16068
rect 24765 16065 24777 16068
rect 24811 16065 24823 16099
rect 24765 16059 24823 16065
rect 24854 16056 24860 16108
rect 24912 16056 24918 16108
rect 25332 16105 25360 16136
rect 25041 16099 25099 16105
rect 25041 16065 25053 16099
rect 25087 16065 25099 16099
rect 25041 16059 25099 16065
rect 25317 16099 25375 16105
rect 25317 16065 25329 16099
rect 25363 16065 25375 16099
rect 25317 16059 25375 16065
rect 15068 16000 16988 16028
rect 15068 15988 15074 16000
rect 17126 15988 17132 16040
rect 17184 15988 17190 16040
rect 25056 16028 25084 16059
rect 25498 16056 25504 16108
rect 25556 16056 25562 16108
rect 25409 16031 25467 16037
rect 25409 16028 25421 16031
rect 25056 16000 25421 16028
rect 25409 15997 25421 16000
rect 25455 15997 25467 16031
rect 25409 15991 25467 15997
rect 16390 15960 16396 15972
rect 13780 15932 16396 15960
rect 13780 15920 13786 15932
rect 16390 15920 16396 15932
rect 16448 15920 16454 15972
rect 17770 15960 17776 15972
rect 16960 15932 17776 15960
rect 16960 15892 16988 15932
rect 17770 15920 17776 15932
rect 17828 15920 17834 15972
rect 13648 15864 16988 15892
rect 17037 15895 17095 15901
rect 12345 15855 12403 15861
rect 17037 15861 17049 15895
rect 17083 15892 17095 15895
rect 17402 15892 17408 15904
rect 17083 15864 17408 15892
rect 17083 15861 17095 15864
rect 17037 15855 17095 15861
rect 17402 15852 17408 15864
rect 17460 15852 17466 15904
rect 25225 15895 25283 15901
rect 25225 15861 25237 15895
rect 25271 15892 25283 15895
rect 25314 15892 25320 15904
rect 25271 15864 25320 15892
rect 25271 15861 25283 15864
rect 25225 15855 25283 15861
rect 25314 15852 25320 15864
rect 25372 15852 25378 15904
rect 1104 15802 27876 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 27876 15802
rect 1104 15728 27876 15750
rect 7742 15648 7748 15700
rect 7800 15688 7806 15700
rect 8113 15691 8171 15697
rect 8113 15688 8125 15691
rect 7800 15660 8125 15688
rect 7800 15648 7806 15660
rect 8113 15657 8125 15660
rect 8159 15657 8171 15691
rect 8113 15651 8171 15657
rect 11698 15648 11704 15700
rect 11756 15688 11762 15700
rect 17129 15691 17187 15697
rect 11756 15660 15148 15688
rect 11756 15648 11762 15660
rect 4157 15623 4215 15629
rect 4157 15589 4169 15623
rect 4203 15620 4215 15623
rect 4203 15592 5028 15620
rect 4203 15589 4215 15592
rect 4157 15583 4215 15589
rect 4341 15555 4399 15561
rect 4341 15521 4353 15555
rect 4387 15552 4399 15555
rect 4614 15552 4620 15564
rect 4387 15524 4620 15552
rect 4387 15521 4399 15524
rect 4341 15515 4399 15521
rect 4614 15512 4620 15524
rect 4672 15512 4678 15564
rect 1949 15487 2007 15493
rect 1949 15453 1961 15487
rect 1995 15484 2007 15487
rect 2774 15484 2780 15496
rect 1995 15456 2780 15484
rect 1995 15453 2007 15456
rect 1949 15447 2007 15453
rect 2774 15444 2780 15456
rect 2832 15444 2838 15496
rect 3970 15484 3976 15496
rect 3344 15456 3976 15484
rect 2216 15419 2274 15425
rect 2216 15385 2228 15419
rect 2262 15416 2274 15419
rect 2498 15416 2504 15428
rect 2262 15388 2504 15416
rect 2262 15385 2274 15388
rect 2216 15379 2274 15385
rect 2498 15376 2504 15388
rect 2556 15376 2562 15428
rect 2774 15308 2780 15360
rect 2832 15348 2838 15360
rect 3344 15357 3372 15456
rect 3970 15444 3976 15456
rect 4028 15484 4034 15496
rect 4433 15487 4491 15493
rect 4433 15484 4445 15487
rect 4028 15456 4445 15484
rect 4028 15444 4034 15456
rect 4433 15453 4445 15456
rect 4479 15453 4491 15487
rect 4433 15447 4491 15453
rect 4706 15444 4712 15496
rect 4764 15444 4770 15496
rect 4801 15487 4859 15493
rect 4801 15453 4813 15487
rect 4847 15453 4859 15487
rect 5000 15484 5028 15592
rect 7650 15580 7656 15632
rect 7708 15620 7714 15632
rect 11790 15620 11796 15632
rect 7708 15592 11796 15620
rect 7708 15580 7714 15592
rect 11790 15580 11796 15592
rect 11848 15580 11854 15632
rect 6178 15512 6184 15564
rect 6236 15512 6242 15564
rect 8110 15512 8116 15564
rect 8168 15552 8174 15564
rect 8168 15524 8340 15552
rect 8168 15512 8174 15524
rect 5077 15487 5135 15493
rect 5077 15484 5089 15487
rect 5000 15456 5089 15484
rect 4801 15447 4859 15453
rect 5077 15453 5089 15456
rect 5123 15484 5135 15487
rect 5123 15456 6040 15484
rect 5123 15453 5135 15456
rect 5077 15447 5135 15453
rect 4724 15416 4752 15444
rect 4632 15388 4752 15416
rect 4816 15416 4844 15447
rect 5718 15416 5724 15428
rect 4816 15388 5724 15416
rect 4632 15357 4660 15388
rect 5718 15376 5724 15388
rect 5776 15376 5782 15428
rect 6012 15416 6040 15456
rect 6086 15444 6092 15496
rect 6144 15484 6150 15496
rect 6546 15484 6552 15496
rect 6144 15456 6552 15484
rect 6144 15444 6150 15456
rect 6546 15444 6552 15456
rect 6604 15444 6610 15496
rect 8018 15444 8024 15496
rect 8076 15444 8082 15496
rect 8312 15493 8340 15524
rect 11974 15512 11980 15564
rect 12032 15552 12038 15564
rect 13814 15552 13820 15564
rect 12032 15524 13820 15552
rect 12032 15512 12038 15524
rect 13814 15512 13820 15524
rect 13872 15512 13878 15564
rect 8205 15487 8263 15493
rect 8205 15453 8217 15487
rect 8251 15453 8263 15487
rect 8205 15447 8263 15453
rect 8297 15487 8355 15493
rect 8297 15453 8309 15487
rect 8343 15453 8355 15487
rect 8297 15447 8355 15453
rect 7650 15416 7656 15428
rect 6012 15388 7656 15416
rect 7650 15376 7656 15388
rect 7708 15376 7714 15428
rect 8220 15416 8248 15447
rect 8386 15444 8392 15496
rect 8444 15444 8450 15496
rect 8478 15444 8484 15496
rect 8536 15444 8542 15496
rect 12526 15444 12532 15496
rect 12584 15484 12590 15496
rect 13081 15487 13139 15493
rect 13081 15484 13093 15487
rect 12584 15456 13093 15484
rect 12584 15444 12590 15456
rect 13081 15453 13093 15456
rect 13127 15453 13139 15487
rect 13081 15447 13139 15453
rect 15010 15444 15016 15496
rect 15068 15444 15074 15496
rect 15120 15484 15148 15660
rect 17129 15657 17141 15691
rect 17175 15688 17187 15691
rect 17678 15688 17684 15700
rect 17175 15660 17684 15688
rect 17175 15657 17187 15660
rect 17129 15651 17187 15657
rect 17678 15648 17684 15660
rect 17736 15648 17742 15700
rect 20349 15691 20407 15697
rect 20349 15657 20361 15691
rect 20395 15657 20407 15691
rect 20349 15651 20407 15657
rect 15289 15623 15347 15629
rect 15289 15589 15301 15623
rect 15335 15620 15347 15623
rect 15746 15620 15752 15632
rect 15335 15592 15752 15620
rect 15335 15589 15347 15592
rect 15289 15583 15347 15589
rect 15746 15580 15752 15592
rect 15804 15580 15810 15632
rect 18969 15623 19027 15629
rect 18969 15620 18981 15623
rect 17512 15592 18981 15620
rect 15289 15487 15347 15493
rect 15289 15484 15301 15487
rect 15120 15456 15301 15484
rect 15289 15453 15301 15456
rect 15335 15484 15347 15487
rect 15378 15484 15384 15496
rect 15335 15456 15384 15484
rect 15335 15453 15347 15456
rect 15289 15447 15347 15453
rect 15378 15444 15384 15456
rect 15436 15444 15442 15496
rect 15470 15444 15476 15496
rect 15528 15484 15534 15496
rect 15749 15487 15807 15493
rect 15749 15484 15761 15487
rect 15528 15456 15761 15484
rect 15528 15444 15534 15456
rect 15749 15453 15761 15456
rect 15795 15453 15807 15487
rect 15749 15447 15807 15453
rect 17402 15444 17408 15496
rect 17460 15444 17466 15496
rect 17512 15493 17540 15592
rect 18969 15589 18981 15592
rect 19015 15589 19027 15623
rect 18969 15583 19027 15589
rect 19242 15580 19248 15632
rect 19300 15580 19306 15632
rect 19889 15623 19947 15629
rect 19889 15620 19901 15623
rect 19720 15592 19901 15620
rect 17678 15512 17684 15564
rect 17736 15552 17742 15564
rect 19720 15561 19748 15592
rect 19889 15589 19901 15592
rect 19935 15589 19947 15623
rect 19889 15583 19947 15589
rect 18509 15555 18567 15561
rect 18509 15552 18521 15555
rect 17736 15524 18521 15552
rect 17736 15512 17742 15524
rect 18509 15521 18521 15524
rect 18555 15521 18567 15555
rect 19705 15555 19763 15561
rect 19705 15552 19717 15555
rect 18509 15515 18567 15521
rect 18892 15524 19717 15552
rect 17497 15487 17555 15493
rect 17497 15453 17509 15487
rect 17543 15453 17555 15487
rect 17497 15447 17555 15453
rect 17586 15444 17592 15496
rect 17644 15444 17650 15496
rect 18892 15493 18920 15524
rect 19705 15521 19717 15524
rect 19751 15521 19763 15555
rect 20364 15552 20392 15651
rect 20806 15648 20812 15700
rect 20864 15688 20870 15700
rect 21634 15688 21640 15700
rect 20864 15660 21640 15688
rect 20864 15648 20870 15660
rect 21634 15648 21640 15660
rect 21692 15688 21698 15700
rect 21913 15691 21971 15697
rect 21913 15688 21925 15691
rect 21692 15660 21925 15688
rect 21692 15648 21698 15660
rect 21913 15657 21925 15660
rect 21959 15688 21971 15691
rect 22002 15688 22008 15700
rect 21959 15660 22008 15688
rect 21959 15657 21971 15660
rect 21913 15651 21971 15657
rect 22002 15648 22008 15660
rect 22060 15648 22066 15700
rect 24949 15691 25007 15697
rect 24949 15657 24961 15691
rect 24995 15688 25007 15691
rect 25498 15688 25504 15700
rect 24995 15660 25504 15688
rect 24995 15657 25007 15660
rect 24949 15651 25007 15657
rect 25498 15648 25504 15660
rect 25556 15648 25562 15700
rect 20622 15580 20628 15632
rect 20680 15620 20686 15632
rect 25593 15623 25651 15629
rect 25593 15620 25605 15623
rect 20680 15592 25605 15620
rect 20680 15580 20686 15592
rect 25593 15589 25605 15592
rect 25639 15589 25651 15623
rect 25593 15583 25651 15589
rect 20364 15524 20944 15552
rect 19705 15515 19763 15521
rect 17865 15487 17923 15493
rect 17865 15453 17877 15487
rect 17911 15484 17923 15487
rect 17957 15487 18015 15493
rect 17957 15484 17969 15487
rect 17911 15456 17969 15484
rect 17911 15453 17923 15456
rect 17865 15447 17923 15453
rect 17957 15453 17969 15456
rect 18003 15453 18015 15487
rect 17957 15447 18015 15453
rect 18877 15487 18935 15493
rect 18877 15453 18889 15487
rect 18923 15453 18935 15487
rect 18877 15447 18935 15453
rect 19061 15487 19119 15493
rect 19061 15453 19073 15487
rect 19107 15484 19119 15487
rect 19426 15484 19432 15496
rect 19107 15456 19432 15484
rect 19107 15453 19119 15456
rect 19061 15447 19119 15453
rect 19426 15444 19432 15456
rect 19484 15444 19490 15496
rect 19613 15487 19671 15493
rect 19613 15453 19625 15487
rect 19659 15453 19671 15487
rect 19613 15447 19671 15453
rect 20165 15487 20223 15493
rect 20165 15453 20177 15487
rect 20211 15484 20223 15487
rect 20346 15484 20352 15496
rect 20211 15456 20352 15484
rect 20211 15453 20223 15456
rect 20165 15447 20223 15453
rect 8404 15416 8432 15444
rect 8846 15416 8852 15428
rect 8220 15388 8852 15416
rect 8846 15376 8852 15388
rect 8904 15376 8910 15428
rect 11146 15376 11152 15428
rect 11204 15416 11210 15428
rect 15105 15419 15163 15425
rect 15105 15416 15117 15419
rect 11204 15388 15117 15416
rect 11204 15376 11210 15388
rect 15105 15385 15117 15388
rect 15151 15416 15163 15419
rect 15562 15416 15568 15428
rect 15151 15388 15568 15416
rect 15151 15385 15163 15388
rect 15105 15379 15163 15385
rect 15562 15376 15568 15388
rect 15620 15376 15626 15428
rect 16016 15419 16074 15425
rect 16016 15385 16028 15419
rect 16062 15416 16074 15419
rect 17221 15419 17279 15425
rect 17221 15416 17233 15419
rect 16062 15388 17233 15416
rect 16062 15385 16074 15388
rect 16016 15379 16074 15385
rect 17221 15385 17233 15388
rect 17267 15385 17279 15419
rect 17221 15379 17279 15385
rect 17727 15419 17785 15425
rect 17727 15385 17739 15419
rect 17773 15416 17785 15419
rect 19628 15416 19656 15447
rect 20346 15444 20352 15456
rect 20404 15444 20410 15496
rect 20441 15487 20499 15493
rect 20441 15453 20453 15487
rect 20487 15484 20499 15487
rect 20806 15484 20812 15496
rect 20487 15456 20812 15484
rect 20487 15453 20499 15456
rect 20441 15447 20499 15453
rect 20806 15444 20812 15456
rect 20864 15444 20870 15496
rect 20916 15493 20944 15524
rect 24670 15512 24676 15564
rect 24728 15512 24734 15564
rect 25038 15512 25044 15564
rect 25096 15552 25102 15564
rect 26053 15555 26111 15561
rect 25096 15524 26004 15552
rect 25096 15512 25102 15524
rect 20901 15487 20959 15493
rect 20901 15453 20913 15487
rect 20947 15484 20959 15487
rect 21266 15484 21272 15496
rect 20947 15456 21272 15484
rect 20947 15453 20959 15456
rect 20901 15447 20959 15453
rect 21266 15444 21272 15456
rect 21324 15444 21330 15496
rect 21450 15444 21456 15496
rect 21508 15444 21514 15496
rect 21542 15444 21548 15496
rect 21600 15444 21606 15496
rect 21729 15487 21787 15493
rect 21729 15453 21741 15487
rect 21775 15453 21787 15487
rect 21729 15447 21787 15453
rect 21174 15416 21180 15428
rect 17773 15388 17908 15416
rect 19628 15388 21180 15416
rect 17773 15385 17785 15388
rect 17727 15379 17785 15385
rect 17880 15360 17908 15388
rect 21174 15376 21180 15388
rect 21232 15376 21238 15428
rect 3329 15351 3387 15357
rect 3329 15348 3341 15351
rect 2832 15320 3341 15348
rect 2832 15308 2838 15320
rect 3329 15317 3341 15320
rect 3375 15317 3387 15351
rect 3329 15311 3387 15317
rect 4617 15351 4675 15357
rect 4617 15317 4629 15351
rect 4663 15317 4675 15351
rect 4617 15311 4675 15317
rect 4709 15351 4767 15357
rect 4709 15317 4721 15351
rect 4755 15348 4767 15351
rect 4798 15348 4804 15360
rect 4755 15320 4804 15348
rect 4755 15317 4767 15320
rect 4709 15311 4767 15317
rect 4798 15308 4804 15320
rect 4856 15308 4862 15360
rect 4985 15351 5043 15357
rect 4985 15317 4997 15351
rect 5031 15348 5043 15351
rect 5350 15348 5356 15360
rect 5031 15320 5356 15348
rect 5031 15317 5043 15320
rect 4985 15311 5043 15317
rect 5350 15308 5356 15320
rect 5408 15308 5414 15360
rect 5445 15351 5503 15357
rect 5445 15317 5457 15351
rect 5491 15348 5503 15351
rect 5534 15348 5540 15360
rect 5491 15320 5540 15348
rect 5491 15317 5503 15320
rect 5445 15311 5503 15317
rect 5534 15308 5540 15320
rect 5592 15308 5598 15360
rect 8386 15308 8392 15360
rect 8444 15308 8450 15360
rect 13173 15351 13231 15357
rect 13173 15317 13185 15351
rect 13219 15348 13231 15351
rect 13262 15348 13268 15360
rect 13219 15320 13268 15348
rect 13219 15317 13231 15320
rect 13173 15311 13231 15317
rect 13262 15308 13268 15320
rect 13320 15308 13326 15360
rect 13446 15308 13452 15360
rect 13504 15348 13510 15360
rect 14090 15348 14096 15360
rect 13504 15320 14096 15348
rect 13504 15308 13510 15320
rect 14090 15308 14096 15320
rect 14148 15348 14154 15360
rect 15194 15348 15200 15360
rect 14148 15320 15200 15348
rect 14148 15308 14154 15320
rect 15194 15308 15200 15320
rect 15252 15308 15258 15360
rect 15378 15308 15384 15360
rect 15436 15348 15442 15360
rect 15654 15348 15660 15360
rect 15436 15320 15660 15348
rect 15436 15308 15442 15320
rect 15654 15308 15660 15320
rect 15712 15308 15718 15360
rect 16390 15308 16396 15360
rect 16448 15348 16454 15360
rect 17126 15348 17132 15360
rect 16448 15320 17132 15348
rect 16448 15308 16454 15320
rect 17126 15308 17132 15320
rect 17184 15308 17190 15360
rect 17862 15308 17868 15360
rect 17920 15308 17926 15360
rect 20070 15308 20076 15360
rect 20128 15348 20134 15360
rect 20533 15351 20591 15357
rect 20533 15348 20545 15351
rect 20128 15320 20545 15348
rect 20128 15308 20134 15320
rect 20533 15317 20545 15320
rect 20579 15317 20591 15351
rect 20533 15311 20591 15317
rect 20714 15308 20720 15360
rect 20772 15348 20778 15360
rect 21744 15348 21772 15447
rect 22186 15444 22192 15496
rect 22244 15484 22250 15496
rect 22465 15487 22523 15493
rect 22465 15484 22477 15487
rect 22244 15456 22477 15484
rect 22244 15444 22250 15456
rect 22465 15453 22477 15456
rect 22511 15453 22523 15487
rect 22465 15447 22523 15453
rect 20772 15320 21772 15348
rect 23124 15348 23152 15470
rect 23566 15444 23572 15496
rect 23624 15484 23630 15496
rect 23694 15487 23752 15493
rect 23694 15484 23706 15487
rect 23624 15456 23706 15484
rect 23624 15444 23630 15456
rect 23694 15453 23706 15456
rect 23740 15453 23752 15487
rect 23694 15447 23752 15453
rect 24118 15444 24124 15496
rect 24176 15444 24182 15496
rect 24210 15444 24216 15496
rect 24268 15484 24274 15496
rect 24581 15487 24639 15493
rect 24581 15484 24593 15487
rect 24268 15456 24593 15484
rect 24268 15444 24274 15456
rect 24581 15453 24593 15456
rect 24627 15453 24639 15487
rect 24581 15447 24639 15453
rect 25222 15444 25228 15496
rect 25280 15444 25286 15496
rect 25976 15493 26004 15524
rect 26053 15521 26065 15555
rect 26099 15552 26111 15555
rect 26329 15555 26387 15561
rect 26329 15552 26341 15555
rect 26099 15524 26341 15552
rect 26099 15521 26111 15524
rect 26053 15515 26111 15521
rect 26329 15521 26341 15524
rect 26375 15521 26387 15555
rect 26329 15515 26387 15521
rect 25961 15487 26019 15493
rect 25961 15453 25973 15487
rect 26007 15453 26019 15487
rect 25961 15447 26019 15453
rect 26237 15487 26295 15493
rect 26237 15453 26249 15487
rect 26283 15453 26295 15487
rect 26237 15447 26295 15453
rect 23477 15419 23535 15425
rect 23477 15385 23489 15419
rect 23523 15416 23535 15419
rect 24946 15416 24952 15428
rect 23523 15388 24952 15416
rect 23523 15385 23535 15388
rect 23477 15379 23535 15385
rect 24946 15376 24952 15388
rect 25004 15376 25010 15428
rect 25314 15376 25320 15428
rect 25372 15416 25378 15428
rect 26252 15416 26280 15447
rect 26418 15444 26424 15496
rect 26476 15444 26482 15496
rect 25372 15388 26280 15416
rect 25372 15376 25378 15388
rect 23569 15351 23627 15357
rect 23569 15348 23581 15351
rect 23124 15320 23581 15348
rect 20772 15308 20778 15320
rect 23569 15317 23581 15320
rect 23615 15317 23627 15351
rect 23569 15311 23627 15317
rect 23753 15351 23811 15357
rect 23753 15317 23765 15351
rect 23799 15348 23811 15351
rect 24026 15348 24032 15360
rect 23799 15320 24032 15348
rect 23799 15317 23811 15320
rect 23753 15311 23811 15317
rect 24026 15308 24032 15320
rect 24084 15348 24090 15360
rect 24578 15348 24584 15360
rect 24084 15320 24584 15348
rect 24084 15308 24090 15320
rect 24578 15308 24584 15320
rect 24636 15308 24642 15360
rect 25041 15351 25099 15357
rect 25041 15317 25053 15351
rect 25087 15348 25099 15351
rect 25130 15348 25136 15360
rect 25087 15320 25136 15348
rect 25087 15317 25099 15320
rect 25041 15311 25099 15317
rect 25130 15308 25136 15320
rect 25188 15308 25194 15360
rect 1104 15258 27876 15280
rect 1104 15206 4874 15258
rect 4926 15206 4938 15258
rect 4990 15206 5002 15258
rect 5054 15206 5066 15258
rect 5118 15206 5130 15258
rect 5182 15206 27876 15258
rect 1104 15184 27876 15206
rect 2498 15104 2504 15156
rect 2556 15104 2562 15156
rect 3878 15104 3884 15156
rect 3936 15144 3942 15156
rect 4325 15147 4383 15153
rect 4325 15144 4337 15147
rect 3936 15116 4337 15144
rect 3936 15104 3942 15116
rect 4325 15113 4337 15116
rect 4371 15144 4383 15147
rect 4371 15116 5120 15144
rect 4371 15113 4383 15116
rect 4325 15107 4383 15113
rect 2225 15079 2283 15085
rect 2225 15045 2237 15079
rect 2271 15076 2283 15079
rect 2774 15076 2780 15088
rect 2271 15048 2780 15076
rect 2271 15045 2283 15048
rect 2225 15039 2283 15045
rect 2774 15036 2780 15048
rect 2832 15036 2838 15088
rect 4525 15079 4583 15085
rect 3436 15048 4016 15076
rect 1946 14968 1952 15020
rect 2004 14968 2010 15020
rect 2038 14968 2044 15020
rect 2096 15008 2102 15020
rect 2133 15011 2191 15017
rect 2133 15008 2145 15011
rect 2096 14980 2145 15008
rect 2096 14968 2102 14980
rect 2133 14977 2145 14980
rect 2179 14977 2191 15011
rect 2133 14971 2191 14977
rect 2314 14968 2320 15020
rect 2372 14968 2378 15020
rect 3234 14968 3240 15020
rect 3292 14968 3298 15020
rect 3436 15017 3464 15048
rect 3421 15011 3479 15017
rect 3421 14977 3433 15011
rect 3467 14977 3479 15011
rect 3421 14971 3479 14977
rect 3878 14968 3884 15020
rect 3936 14968 3942 15020
rect 3988 15008 4016 15048
rect 4525 15045 4537 15079
rect 4571 15045 4583 15079
rect 4525 15039 4583 15045
rect 5092 15076 5120 15116
rect 8386 15104 8392 15156
rect 8444 15144 8450 15156
rect 8941 15147 8999 15153
rect 8941 15144 8953 15147
rect 8444 15116 8953 15144
rect 8444 15104 8450 15116
rect 8941 15113 8953 15116
rect 8987 15113 8999 15147
rect 9674 15144 9680 15156
rect 8941 15107 8999 15113
rect 9232 15116 9680 15144
rect 5994 15076 6000 15088
rect 5092 15048 6000 15076
rect 4062 15008 4068 15020
rect 3988 14980 4068 15008
rect 4062 14968 4068 14980
rect 4120 15008 4126 15020
rect 4540 15008 4568 15039
rect 4801 15011 4859 15017
rect 4801 15008 4813 15011
rect 4120 14980 4813 15008
rect 4120 14968 4126 14980
rect 4801 14977 4813 14980
rect 4847 14977 4859 15011
rect 4801 14971 4859 14977
rect 4982 14968 4988 15020
rect 5040 14968 5046 15020
rect 5092 15017 5120 15048
rect 5994 15036 6000 15048
rect 6052 15036 6058 15088
rect 7650 15036 7656 15088
rect 7708 15076 7714 15088
rect 9030 15076 9036 15088
rect 7708 15048 9036 15076
rect 7708 15036 7714 15048
rect 9030 15036 9036 15048
rect 9088 15036 9094 15088
rect 5077 15011 5135 15017
rect 5077 14977 5089 15011
rect 5123 14977 5135 15011
rect 5077 14971 5135 14977
rect 5718 14968 5724 15020
rect 5776 14968 5782 15020
rect 5905 15011 5963 15017
rect 5905 14977 5917 15011
rect 5951 15008 5963 15011
rect 6086 15008 6092 15020
rect 5951 14980 6092 15008
rect 5951 14977 5963 14980
rect 5905 14971 5963 14977
rect 6086 14968 6092 14980
rect 6144 14968 6150 15020
rect 7190 14968 7196 15020
rect 7248 14968 7254 15020
rect 7282 14968 7288 15020
rect 7340 15008 7346 15020
rect 9232 15008 9260 15116
rect 9674 15104 9680 15116
rect 9732 15144 9738 15156
rect 10962 15144 10968 15156
rect 9732 15116 10968 15144
rect 9732 15104 9738 15116
rect 10962 15104 10968 15116
rect 11020 15104 11026 15156
rect 11333 15147 11391 15153
rect 11333 15113 11345 15147
rect 11379 15113 11391 15147
rect 11333 15107 11391 15113
rect 10686 15076 10692 15088
rect 9416 15048 10692 15076
rect 9416 15017 9444 15048
rect 10686 15036 10692 15048
rect 10744 15036 10750 15088
rect 11348 15076 11376 15107
rect 11882 15104 11888 15156
rect 11940 15144 11946 15156
rect 12342 15144 12348 15156
rect 11940 15116 12348 15144
rect 11940 15104 11946 15116
rect 12342 15104 12348 15116
rect 12400 15144 12406 15156
rect 14093 15147 14151 15153
rect 14093 15144 14105 15147
rect 12400 15116 14105 15144
rect 12400 15104 12406 15116
rect 14093 15113 14105 15116
rect 14139 15113 14151 15147
rect 14093 15107 14151 15113
rect 14734 15104 14740 15156
rect 14792 15104 14798 15156
rect 14936 15116 15424 15144
rect 11762 15079 11820 15085
rect 11762 15076 11774 15079
rect 10796 15048 11284 15076
rect 11348 15048 11774 15076
rect 7340 14980 9260 15008
rect 9401 15011 9459 15017
rect 7340 14968 7346 14980
rect 9401 14977 9413 15011
rect 9447 14977 9459 15011
rect 9401 14971 9459 14977
rect 9674 14968 9680 15020
rect 9732 15008 9738 15020
rect 10229 15011 10287 15017
rect 10229 15008 10241 15011
rect 9732 14980 10241 15008
rect 9732 14968 9738 14980
rect 10229 14977 10241 14980
rect 10275 14977 10287 15011
rect 10229 14971 10287 14977
rect 10413 15011 10471 15017
rect 10413 14977 10425 15011
rect 10459 15008 10471 15011
rect 10459 14980 10548 15008
rect 10459 14977 10471 14980
rect 10413 14971 10471 14977
rect 10520 14952 10548 14980
rect 10594 14968 10600 15020
rect 10652 14968 10658 15020
rect 10796 15017 10824 15048
rect 10781 15011 10839 15017
rect 10781 14977 10793 15011
rect 10827 14977 10839 15011
rect 10781 14971 10839 14977
rect 10965 15011 11023 15017
rect 10965 14977 10977 15011
rect 11011 14977 11023 15011
rect 10965 14971 11023 14977
rect 3053 14943 3111 14949
rect 3053 14909 3065 14943
rect 3099 14940 3111 14943
rect 3697 14943 3755 14949
rect 3697 14940 3709 14943
rect 3099 14912 3709 14940
rect 3099 14909 3111 14912
rect 3053 14903 3111 14909
rect 3697 14909 3709 14912
rect 3743 14940 3755 14943
rect 4706 14940 4712 14952
rect 3743 14912 4712 14940
rect 3743 14909 3755 14912
rect 3697 14903 3755 14909
rect 4706 14900 4712 14912
rect 4764 14900 4770 14952
rect 8846 14900 8852 14952
rect 8904 14900 8910 14952
rect 9769 14943 9827 14949
rect 9769 14909 9781 14943
rect 9815 14909 9827 14943
rect 9769 14903 9827 14909
rect 9861 14943 9919 14949
rect 9861 14909 9873 14943
rect 9907 14909 9919 14943
rect 9861 14903 9919 14909
rect 4154 14832 4160 14884
rect 4212 14832 4218 14884
rect 4982 14872 4988 14884
rect 4356 14844 4988 14872
rect 3970 14764 3976 14816
rect 4028 14804 4034 14816
rect 4356 14813 4384 14844
rect 4982 14832 4988 14844
rect 5040 14832 5046 14884
rect 8481 14875 8539 14881
rect 8481 14841 8493 14875
rect 8527 14872 8539 14875
rect 8754 14872 8760 14884
rect 8527 14844 8760 14872
rect 8527 14841 8539 14844
rect 8481 14835 8539 14841
rect 8754 14832 8760 14844
rect 8812 14832 8818 14884
rect 8938 14832 8944 14884
rect 8996 14872 9002 14884
rect 9493 14875 9551 14881
rect 9493 14872 9505 14875
rect 8996 14844 9505 14872
rect 8996 14832 9002 14844
rect 9493 14841 9505 14844
rect 9539 14841 9551 14875
rect 9493 14835 9551 14841
rect 4065 14807 4123 14813
rect 4065 14804 4077 14807
rect 4028 14776 4077 14804
rect 4028 14764 4034 14776
rect 4065 14773 4077 14776
rect 4111 14773 4123 14807
rect 4065 14767 4123 14773
rect 4341 14807 4399 14813
rect 4341 14773 4353 14807
rect 4387 14773 4399 14807
rect 4341 14767 4399 14773
rect 4614 14764 4620 14816
rect 4672 14764 4678 14816
rect 5902 14764 5908 14816
rect 5960 14764 5966 14816
rect 6089 14807 6147 14813
rect 6089 14773 6101 14807
rect 6135 14804 6147 14807
rect 6362 14804 6368 14816
rect 6135 14776 6368 14804
rect 6135 14773 6147 14776
rect 6089 14767 6147 14773
rect 6362 14764 6368 14776
rect 6420 14764 6426 14816
rect 6546 14764 6552 14816
rect 6604 14764 6610 14816
rect 8662 14764 8668 14816
rect 8720 14804 8726 14816
rect 9309 14807 9367 14813
rect 9309 14804 9321 14807
rect 8720 14776 9321 14804
rect 8720 14764 8726 14776
rect 9309 14773 9321 14776
rect 9355 14773 9367 14807
rect 9784 14804 9812 14903
rect 9876 14872 9904 14903
rect 9950 14900 9956 14952
rect 10008 14900 10014 14952
rect 10134 14900 10140 14952
rect 10192 14940 10198 14952
rect 10192 14912 10456 14940
rect 10192 14900 10198 14912
rect 10042 14872 10048 14884
rect 9876 14844 10048 14872
rect 10042 14832 10048 14844
rect 10100 14832 10106 14884
rect 10428 14872 10456 14912
rect 10502 14900 10508 14952
rect 10560 14940 10566 14952
rect 10870 14940 10876 14952
rect 10560 14912 10876 14940
rect 10560 14900 10566 14912
rect 10870 14900 10876 14912
rect 10928 14900 10934 14952
rect 10980 14872 11008 14971
rect 11054 14968 11060 15020
rect 11112 14968 11118 15020
rect 11146 14968 11152 15020
rect 11204 14968 11210 15020
rect 11256 15008 11284 15048
rect 11762 15045 11774 15048
rect 11808 15045 11820 15079
rect 11762 15039 11820 15045
rect 13449 15079 13507 15085
rect 13449 15045 13461 15079
rect 13495 15076 13507 15079
rect 13722 15076 13728 15088
rect 13495 15048 13728 15076
rect 13495 15045 13507 15048
rect 13449 15039 13507 15045
rect 13722 15036 13728 15048
rect 13780 15036 13786 15088
rect 13814 15036 13820 15088
rect 13872 15036 13878 15088
rect 13081 15011 13139 15017
rect 13081 15008 13093 15011
rect 11256 14980 13093 15008
rect 13081 14977 13093 14980
rect 13127 14977 13139 15011
rect 13081 14971 13139 14977
rect 13262 14968 13268 15020
rect 13320 14968 13326 15020
rect 13357 15011 13415 15017
rect 13357 14977 13369 15011
rect 13403 14977 13415 15011
rect 13357 14971 13415 14977
rect 13587 15011 13645 15017
rect 13587 14977 13599 15011
rect 13633 15008 13645 15011
rect 13633 14980 13952 15008
rect 13633 14977 13645 14980
rect 13587 14971 13645 14977
rect 11517 14943 11575 14949
rect 11517 14909 11529 14943
rect 11563 14909 11575 14943
rect 11517 14903 11575 14909
rect 10428 14844 11008 14872
rect 10134 14804 10140 14816
rect 9784 14776 10140 14804
rect 9309 14767 9367 14773
rect 10134 14764 10140 14776
rect 10192 14764 10198 14816
rect 11532 14804 11560 14903
rect 13170 14900 13176 14952
rect 13228 14940 13234 14952
rect 13372 14940 13400 14971
rect 13228 14912 13400 14940
rect 13228 14900 13234 14912
rect 13722 14900 13728 14952
rect 13780 14900 13786 14952
rect 13924 14940 13952 14980
rect 13998 14968 14004 15020
rect 14056 14968 14062 15020
rect 14182 14968 14188 15020
rect 14240 14968 14246 15020
rect 14936 15017 14964 15116
rect 15102 15036 15108 15088
rect 15160 15036 15166 15088
rect 15194 15036 15200 15088
rect 15252 15085 15258 15088
rect 15252 15079 15281 15085
rect 15269 15045 15281 15079
rect 15396 15076 15424 15116
rect 15838 15104 15844 15156
rect 15896 15144 15902 15156
rect 16761 15147 16819 15153
rect 15896 15116 16344 15144
rect 15896 15104 15902 15116
rect 16316 15088 16344 15116
rect 16761 15113 16773 15147
rect 16807 15144 16819 15147
rect 16850 15144 16856 15156
rect 16807 15116 16856 15144
rect 16807 15113 16819 15116
rect 16761 15107 16819 15113
rect 16850 15104 16856 15116
rect 16908 15104 16914 15156
rect 17037 15147 17095 15153
rect 17037 15113 17049 15147
rect 17083 15113 17095 15147
rect 17037 15107 17095 15113
rect 16209 15079 16267 15085
rect 16209 15076 16221 15079
rect 15396 15048 16221 15076
rect 15252 15039 15281 15045
rect 16209 15045 16221 15048
rect 16255 15045 16267 15079
rect 16209 15039 16267 15045
rect 15252 15036 15258 15039
rect 16298 15036 16304 15088
rect 16356 15076 16362 15088
rect 17052 15076 17080 15107
rect 17770 15104 17776 15156
rect 17828 15104 17834 15156
rect 19981 15147 20039 15153
rect 19981 15113 19993 15147
rect 20027 15144 20039 15147
rect 20346 15144 20352 15156
rect 20027 15116 20352 15144
rect 20027 15113 20039 15116
rect 19981 15107 20039 15113
rect 20346 15104 20352 15116
rect 20404 15104 20410 15156
rect 20993 15147 21051 15153
rect 20993 15144 21005 15147
rect 20640 15116 21005 15144
rect 16356 15048 17080 15076
rect 17129 15079 17187 15085
rect 16356 15036 16362 15048
rect 14921 15011 14979 15017
rect 14921 14977 14933 15011
rect 14967 14977 14979 15011
rect 14921 14971 14979 14977
rect 15013 15011 15071 15017
rect 15013 14977 15025 15011
rect 15059 14977 15071 15011
rect 15013 14971 15071 14977
rect 15212 14980 15608 15008
rect 14734 14940 14740 14952
rect 13924 14912 14740 14940
rect 14734 14900 14740 14912
rect 14792 14900 14798 14952
rect 15028 14940 15056 14971
rect 15212 14940 15240 14980
rect 15028 14912 15240 14940
rect 15378 14900 15384 14952
rect 15436 14900 15442 14952
rect 15473 14943 15531 14949
rect 15473 14909 15485 14943
rect 15519 14909 15531 14943
rect 15580 14940 15608 14980
rect 15654 14968 15660 15020
rect 15712 14968 15718 15020
rect 15746 14968 15752 15020
rect 15804 15008 15810 15020
rect 16684 15017 16712 15048
rect 17129 15045 17141 15079
rect 17175 15076 17187 15079
rect 17678 15076 17684 15088
rect 17175 15048 17684 15076
rect 17175 15045 17187 15048
rect 17129 15039 17187 15045
rect 17678 15036 17684 15048
rect 17736 15036 17742 15088
rect 18049 15079 18107 15085
rect 18049 15045 18061 15079
rect 18095 15076 18107 15079
rect 20162 15076 20168 15088
rect 18095 15048 20168 15076
rect 18095 15045 18107 15048
rect 18049 15039 18107 15045
rect 20162 15036 20168 15048
rect 20220 15036 20226 15088
rect 15933 15011 15991 15017
rect 15933 15008 15945 15011
rect 15804 14980 15945 15008
rect 15804 14968 15810 14980
rect 15933 14977 15945 14980
rect 15979 14977 15991 15011
rect 16669 15011 16727 15017
rect 15933 14971 15991 14977
rect 16040 14980 16620 15008
rect 16040 14940 16068 14980
rect 15580 14912 16068 14940
rect 16209 14943 16267 14949
rect 15473 14903 15531 14909
rect 16209 14909 16221 14943
rect 16255 14940 16267 14943
rect 16390 14940 16396 14952
rect 16255 14912 16396 14940
rect 16255 14909 16267 14912
rect 16209 14903 16267 14909
rect 12710 14832 12716 14884
rect 12768 14872 12774 14884
rect 13354 14872 13360 14884
rect 12768 14844 13360 14872
rect 12768 14832 12774 14844
rect 13354 14832 13360 14844
rect 13412 14832 13418 14884
rect 13814 14832 13820 14884
rect 13872 14872 13878 14884
rect 15488 14872 15516 14903
rect 16390 14900 16396 14912
rect 16448 14900 16454 14952
rect 16592 14940 16620 14980
rect 16669 14977 16681 15011
rect 16715 14977 16727 15011
rect 16669 14971 16727 14977
rect 16758 14968 16764 15020
rect 16816 15008 16822 15020
rect 16853 15011 16911 15017
rect 16853 15008 16865 15011
rect 16816 14980 16865 15008
rect 16816 14968 16822 14980
rect 16853 14977 16865 14980
rect 16899 14977 16911 15011
rect 16853 14971 16911 14977
rect 17954 14968 17960 15020
rect 18012 14968 18018 15020
rect 18138 14968 18144 15020
rect 18196 14968 18202 15020
rect 18230 14968 18236 15020
rect 18288 15008 18294 15020
rect 18325 15011 18383 15017
rect 18325 15008 18337 15011
rect 18288 14980 18337 15008
rect 18288 14968 18294 14980
rect 18325 14977 18337 14980
rect 18371 15008 18383 15011
rect 18782 15008 18788 15020
rect 18371 14980 18788 15008
rect 18371 14977 18383 14980
rect 18325 14971 18383 14977
rect 18782 14968 18788 14980
rect 18840 14968 18846 15020
rect 18966 14968 18972 15020
rect 19024 15008 19030 15020
rect 19797 15011 19855 15017
rect 19797 15008 19809 15011
rect 19024 14980 19809 15008
rect 19024 14968 19030 14980
rect 19797 14977 19809 14980
rect 19843 14977 19855 15011
rect 19797 14971 19855 14977
rect 20070 14968 20076 15020
rect 20128 14968 20134 15020
rect 20640 15017 20668 15116
rect 20993 15113 21005 15116
rect 21039 15144 21051 15147
rect 22278 15144 22284 15156
rect 21039 15116 22284 15144
rect 21039 15113 21051 15116
rect 20993 15107 21051 15113
rect 22278 15104 22284 15116
rect 22336 15104 22342 15156
rect 22465 15147 22523 15153
rect 22465 15113 22477 15147
rect 22511 15113 22523 15147
rect 22465 15107 22523 15113
rect 23845 15147 23903 15153
rect 23845 15113 23857 15147
rect 23891 15144 23903 15147
rect 24118 15144 24124 15156
rect 23891 15116 24124 15144
rect 23891 15113 23903 15116
rect 23845 15107 23903 15113
rect 20717 15079 20775 15085
rect 20717 15045 20729 15079
rect 20763 15076 20775 15079
rect 22480 15076 22508 15107
rect 24118 15104 24124 15116
rect 24176 15104 24182 15156
rect 24486 15104 24492 15156
rect 24544 15144 24550 15156
rect 24673 15147 24731 15153
rect 24673 15144 24685 15147
rect 24544 15116 24685 15144
rect 24544 15104 24550 15116
rect 24673 15113 24685 15116
rect 24719 15113 24731 15147
rect 24673 15107 24731 15113
rect 24854 15104 24860 15156
rect 24912 15104 24918 15156
rect 25130 15104 25136 15156
rect 25188 15104 25194 15156
rect 20763 15048 21036 15076
rect 20763 15045 20775 15048
rect 20717 15039 20775 15045
rect 21008 15020 21036 15048
rect 21100 15048 22508 15076
rect 24136 15076 24164 15104
rect 24949 15079 25007 15085
rect 24949 15076 24961 15079
rect 24136 15048 24961 15076
rect 20625 15011 20683 15017
rect 20625 14977 20637 15011
rect 20671 14977 20683 15011
rect 20625 14971 20683 14977
rect 20898 14968 20904 15020
rect 20956 14968 20962 15020
rect 20990 14968 20996 15020
rect 21048 14968 21054 15020
rect 21100 14940 21128 15048
rect 24949 15045 24961 15048
rect 24995 15045 25007 15079
rect 24949 15039 25007 15045
rect 21174 14968 21180 15020
rect 21232 14968 21238 15020
rect 21266 14968 21272 15020
rect 21324 14968 21330 15020
rect 21634 14968 21640 15020
rect 21692 14968 21698 15020
rect 21818 14968 21824 15020
rect 21876 14968 21882 15020
rect 21913 15011 21971 15017
rect 21913 14977 21925 15011
rect 21959 14977 21971 15011
rect 21913 14971 21971 14977
rect 16592 14912 21128 14940
rect 15562 14872 15568 14884
rect 13872 14844 15424 14872
rect 15488 14844 15568 14872
rect 13872 14832 13878 14844
rect 12728 14804 12756 14832
rect 15396 14816 15424 14844
rect 15562 14832 15568 14844
rect 15620 14832 15626 14884
rect 17218 14832 17224 14884
rect 17276 14872 17282 14884
rect 18966 14872 18972 14884
rect 17276 14844 18972 14872
rect 17276 14832 17282 14844
rect 18966 14832 18972 14844
rect 19024 14832 19030 14884
rect 19426 14832 19432 14884
rect 19484 14872 19490 14884
rect 19797 14875 19855 14881
rect 19797 14872 19809 14875
rect 19484 14844 19809 14872
rect 19484 14832 19490 14844
rect 19797 14841 19809 14844
rect 19843 14841 19855 14875
rect 19797 14835 19855 14841
rect 20901 14875 20959 14881
rect 20901 14841 20913 14875
rect 20947 14872 20959 14875
rect 21928 14872 21956 14971
rect 22002 14968 22008 15020
rect 22060 15008 22066 15020
rect 22097 15011 22155 15017
rect 22097 15008 22109 15011
rect 22060 14980 22109 15008
rect 22060 14968 22066 14980
rect 22097 14977 22109 14980
rect 22143 14977 22155 15011
rect 22097 14971 22155 14977
rect 22189 15011 22247 15017
rect 22189 14977 22201 15011
rect 22235 14977 22247 15011
rect 22189 14971 22247 14977
rect 22204 14940 22232 14971
rect 22278 14968 22284 15020
rect 22336 14968 22342 15020
rect 23198 14968 23204 15020
rect 23256 15008 23262 15020
rect 23753 15011 23811 15017
rect 23753 15008 23765 15011
rect 23256 14980 23765 15008
rect 23256 14968 23262 14980
rect 23753 14977 23765 14980
rect 23799 14977 23811 15011
rect 23753 14971 23811 14977
rect 23768 14940 23796 14971
rect 23934 14968 23940 15020
rect 23992 14968 23998 15020
rect 24670 14968 24676 15020
rect 24728 15008 24734 15020
rect 25225 15011 25283 15017
rect 24728 14980 24808 15008
rect 24728 14968 24734 14980
rect 24213 14943 24271 14949
rect 24213 14940 24225 14943
rect 22204 14912 22324 14940
rect 23768 14912 24225 14940
rect 22296 14884 22324 14912
rect 24213 14909 24225 14912
rect 24259 14909 24271 14943
rect 24213 14903 24271 14909
rect 20947 14844 21956 14872
rect 20947 14841 20959 14844
rect 20901 14835 20959 14841
rect 22278 14832 22284 14884
rect 22336 14832 22342 14884
rect 24780 14872 24808 14980
rect 25225 14977 25237 15011
rect 25271 14977 25283 15011
rect 25225 14971 25283 14977
rect 24949 14875 25007 14881
rect 24949 14872 24961 14875
rect 24780 14844 24961 14872
rect 24949 14841 24961 14844
rect 24995 14841 25007 14875
rect 24949 14835 25007 14841
rect 11532 14776 12756 14804
rect 12897 14807 12955 14813
rect 12897 14773 12909 14807
rect 12943 14804 12955 14807
rect 12986 14804 12992 14816
rect 12943 14776 12992 14804
rect 12943 14773 12955 14776
rect 12897 14767 12955 14773
rect 12986 14764 12992 14776
rect 13044 14764 13050 14816
rect 14366 14764 14372 14816
rect 14424 14764 14430 14816
rect 15378 14764 15384 14816
rect 15436 14764 15442 14816
rect 15838 14764 15844 14816
rect 15896 14764 15902 14816
rect 16022 14764 16028 14816
rect 16080 14764 16086 14816
rect 16666 14764 16672 14816
rect 16724 14804 16730 14816
rect 18414 14804 18420 14816
rect 16724 14776 18420 14804
rect 16724 14764 16730 14776
rect 18414 14764 18420 14776
rect 18472 14804 18478 14816
rect 18874 14804 18880 14816
rect 18472 14776 18880 14804
rect 18472 14764 18478 14776
rect 18874 14764 18880 14776
rect 18932 14764 18938 14816
rect 20622 14764 20628 14816
rect 20680 14804 20686 14816
rect 21177 14807 21235 14813
rect 21177 14804 21189 14807
rect 20680 14776 21189 14804
rect 20680 14764 20686 14776
rect 21177 14773 21189 14776
rect 21223 14773 21235 14807
rect 21177 14767 21235 14773
rect 24302 14764 24308 14816
rect 24360 14764 24366 14816
rect 24578 14764 24584 14816
rect 24636 14804 24642 14816
rect 25240 14804 25268 14971
rect 24636 14776 25268 14804
rect 24636 14764 24642 14776
rect 1104 14714 27876 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 27876 14714
rect 1104 14640 27876 14662
rect 1946 14560 1952 14612
rect 2004 14560 2010 14612
rect 4982 14560 4988 14612
rect 5040 14600 5046 14612
rect 5350 14600 5356 14612
rect 5040 14572 5356 14600
rect 5040 14560 5046 14572
rect 5350 14560 5356 14572
rect 5408 14600 5414 14612
rect 10134 14600 10140 14612
rect 5408 14572 10140 14600
rect 5408 14560 5414 14572
rect 2774 14532 2780 14544
rect 1596 14504 2780 14532
rect 1596 14405 1624 14504
rect 2774 14492 2780 14504
rect 2832 14532 2838 14544
rect 3694 14532 3700 14544
rect 2832 14504 3700 14532
rect 2832 14492 2838 14504
rect 3694 14492 3700 14504
rect 3752 14492 3758 14544
rect 3970 14492 3976 14544
rect 4028 14532 4034 14544
rect 7190 14532 7196 14544
rect 4028 14504 4476 14532
rect 4028 14492 4034 14504
rect 1673 14467 1731 14473
rect 1673 14433 1685 14467
rect 1719 14433 1731 14467
rect 1673 14427 1731 14433
rect 1581 14399 1639 14405
rect 1581 14365 1593 14399
rect 1627 14365 1639 14399
rect 1688 14396 1716 14427
rect 3234 14424 3240 14476
rect 3292 14464 3298 14476
rect 4448 14473 4476 14504
rect 6748 14504 7196 14532
rect 6748 14473 6776 14504
rect 7190 14492 7196 14504
rect 7248 14492 7254 14544
rect 4433 14467 4491 14473
rect 3292 14436 4016 14464
rect 3292 14424 3298 14436
rect 1854 14396 1860 14408
rect 1688 14368 1860 14396
rect 1581 14359 1639 14365
rect 1854 14356 1860 14368
rect 1912 14396 1918 14408
rect 2041 14399 2099 14405
rect 2041 14396 2053 14399
rect 1912 14368 2053 14396
rect 1912 14356 1918 14368
rect 2041 14365 2053 14368
rect 2087 14365 2099 14399
rect 2041 14359 2099 14365
rect 2130 14356 2136 14408
rect 2188 14396 2194 14408
rect 2225 14399 2283 14405
rect 2225 14396 2237 14399
rect 2188 14368 2237 14396
rect 2188 14356 2194 14368
rect 2225 14365 2237 14368
rect 2271 14365 2283 14399
rect 2225 14359 2283 14365
rect 3602 14356 3608 14408
rect 3660 14356 3666 14408
rect 3988 14405 4016 14436
rect 4433 14433 4445 14467
rect 4479 14433 4491 14467
rect 4433 14427 4491 14433
rect 6733 14467 6791 14473
rect 6733 14433 6745 14467
rect 6779 14433 6791 14467
rect 6733 14427 6791 14433
rect 7009 14467 7067 14473
rect 7009 14433 7021 14467
rect 7055 14464 7067 14467
rect 7374 14464 7380 14476
rect 7055 14436 7380 14464
rect 7055 14433 7067 14436
rect 7009 14427 7067 14433
rect 7374 14424 7380 14436
rect 7432 14424 7438 14476
rect 7742 14424 7748 14476
rect 7800 14464 7806 14476
rect 8496 14473 8524 14572
rect 10134 14560 10140 14572
rect 10192 14600 10198 14612
rect 10229 14603 10287 14609
rect 10229 14600 10241 14603
rect 10192 14572 10241 14600
rect 10192 14560 10198 14572
rect 10229 14569 10241 14572
rect 10275 14569 10287 14603
rect 10229 14563 10287 14569
rect 10962 14560 10968 14612
rect 11020 14600 11026 14612
rect 12986 14600 12992 14612
rect 11020 14572 12992 14600
rect 11020 14560 11026 14572
rect 12986 14560 12992 14572
rect 13044 14560 13050 14612
rect 13170 14560 13176 14612
rect 13228 14560 13234 14612
rect 13998 14600 14004 14612
rect 13648 14572 14004 14600
rect 8846 14492 8852 14544
rect 8904 14532 8910 14544
rect 8904 14504 10732 14532
rect 8904 14492 8910 14504
rect 8389 14467 8447 14473
rect 8389 14464 8401 14467
rect 7800 14436 8401 14464
rect 7800 14424 7806 14436
rect 8389 14433 8401 14436
rect 8435 14433 8447 14467
rect 8389 14427 8447 14433
rect 8481 14467 8539 14473
rect 8481 14433 8493 14467
rect 8527 14433 8539 14467
rect 8481 14427 8539 14433
rect 8662 14424 8668 14476
rect 8720 14424 8726 14476
rect 9030 14424 9036 14476
rect 9088 14464 9094 14476
rect 10704 14464 10732 14504
rect 10778 14492 10784 14544
rect 10836 14492 10842 14544
rect 13648 14532 13676 14572
rect 13998 14560 14004 14572
rect 14056 14560 14062 14612
rect 14182 14560 14188 14612
rect 14240 14600 14246 14612
rect 14829 14603 14887 14609
rect 14829 14600 14841 14603
rect 14240 14572 14841 14600
rect 14240 14560 14246 14572
rect 14829 14569 14841 14572
rect 14875 14600 14887 14603
rect 16022 14600 16028 14612
rect 14875 14572 16028 14600
rect 14875 14569 14887 14572
rect 14829 14563 14887 14569
rect 16022 14560 16028 14572
rect 16080 14560 16086 14612
rect 18138 14560 18144 14612
rect 18196 14600 18202 14612
rect 18509 14603 18567 14609
rect 18509 14600 18521 14603
rect 18196 14572 18521 14600
rect 18196 14560 18202 14572
rect 18509 14569 18521 14572
rect 18555 14569 18567 14603
rect 18509 14563 18567 14569
rect 21174 14560 21180 14612
rect 21232 14600 21238 14612
rect 21637 14603 21695 14609
rect 21637 14600 21649 14603
rect 21232 14572 21649 14600
rect 21232 14560 21238 14572
rect 21637 14569 21649 14572
rect 21683 14600 21695 14603
rect 22373 14603 22431 14609
rect 22373 14600 22385 14603
rect 21683 14572 22385 14600
rect 21683 14569 21695 14572
rect 21637 14563 21695 14569
rect 22373 14569 22385 14572
rect 22419 14569 22431 14603
rect 24118 14600 24124 14612
rect 22373 14563 22431 14569
rect 22664 14572 24124 14600
rect 12636 14504 13676 14532
rect 12636 14464 12664 14504
rect 13722 14492 13728 14544
rect 13780 14532 13786 14544
rect 17865 14535 17923 14541
rect 17865 14532 17877 14535
rect 13780 14504 17877 14532
rect 13780 14492 13786 14504
rect 17865 14501 17877 14504
rect 17911 14501 17923 14535
rect 17865 14495 17923 14501
rect 18248 14504 20116 14532
rect 12894 14464 12900 14476
rect 9088 14436 10640 14464
rect 10704 14436 12664 14464
rect 12728 14436 12900 14464
rect 9088 14424 9094 14436
rect 3973 14399 4031 14405
rect 3973 14365 3985 14399
rect 4019 14365 4031 14399
rect 3973 14359 4031 14365
rect 4062 14356 4068 14408
rect 4120 14356 4126 14408
rect 4341 14399 4399 14405
rect 4341 14365 4353 14399
rect 4387 14396 4399 14399
rect 4982 14396 4988 14408
rect 4387 14368 4988 14396
rect 4387 14365 4399 14368
rect 4341 14359 4399 14365
rect 4982 14356 4988 14368
rect 5040 14356 5046 14408
rect 6641 14399 6699 14405
rect 6641 14365 6653 14399
rect 6687 14396 6699 14399
rect 7282 14396 7288 14408
rect 6687 14368 7288 14396
rect 6687 14365 6699 14368
rect 6641 14359 6699 14365
rect 7282 14356 7288 14368
rect 7340 14356 7346 14408
rect 8570 14356 8576 14408
rect 8628 14356 8634 14408
rect 9493 14399 9551 14405
rect 9493 14365 9505 14399
rect 9539 14365 9551 14399
rect 9493 14359 9551 14365
rect 1394 14288 1400 14340
rect 1452 14328 1458 14340
rect 2866 14328 2872 14340
rect 1452 14300 2872 14328
rect 1452 14288 1458 14300
rect 2866 14288 2872 14300
rect 2924 14288 2930 14340
rect 9508 14328 9536 14359
rect 9674 14356 9680 14408
rect 9732 14396 9738 14408
rect 10612 14405 10640 14436
rect 10505 14399 10563 14405
rect 10505 14396 10517 14399
rect 9732 14368 10517 14396
rect 9732 14356 9738 14368
rect 9766 14328 9772 14340
rect 9508 14300 9772 14328
rect 9766 14288 9772 14300
rect 9824 14288 9830 14340
rect 10042 14288 10048 14340
rect 10100 14288 10106 14340
rect 10244 14337 10272 14368
rect 10505 14365 10517 14368
rect 10551 14365 10563 14399
rect 10505 14359 10563 14365
rect 10597 14399 10655 14405
rect 10597 14365 10609 14399
rect 10643 14365 10655 14399
rect 10597 14359 10655 14365
rect 10781 14399 10839 14405
rect 10781 14365 10793 14399
rect 10827 14396 10839 14399
rect 11238 14396 11244 14408
rect 10827 14368 11244 14396
rect 10827 14365 10839 14368
rect 10781 14359 10839 14365
rect 10244 14331 10303 14337
rect 10244 14300 10257 14331
rect 10245 14297 10257 14300
rect 10291 14297 10303 14331
rect 10796 14328 10824 14359
rect 11238 14356 11244 14368
rect 11296 14356 11302 14408
rect 12728 14405 12756 14436
rect 12894 14424 12900 14436
rect 12952 14464 12958 14476
rect 14366 14464 14372 14476
rect 12952 14436 14372 14464
rect 12952 14424 12958 14436
rect 14366 14424 14372 14436
rect 14424 14424 14430 14476
rect 14734 14424 14740 14476
rect 14792 14464 14798 14476
rect 18248 14464 18276 14504
rect 20088 14464 20116 14504
rect 20162 14492 20168 14544
rect 20220 14532 20226 14544
rect 22664 14532 22692 14572
rect 24118 14560 24124 14572
rect 24176 14560 24182 14612
rect 24486 14560 24492 14612
rect 24544 14560 24550 14612
rect 20220 14504 22692 14532
rect 20220 14492 20226 14504
rect 22738 14492 22744 14544
rect 22796 14532 22802 14544
rect 23106 14532 23112 14544
rect 22796 14504 23112 14532
rect 22796 14492 22802 14504
rect 23106 14492 23112 14504
rect 23164 14532 23170 14544
rect 23293 14535 23351 14541
rect 23293 14532 23305 14535
rect 23164 14504 23305 14532
rect 23164 14492 23170 14504
rect 23293 14501 23305 14504
rect 23339 14501 23351 14535
rect 23293 14495 23351 14501
rect 20438 14464 20444 14476
rect 14792 14436 18276 14464
rect 18340 14436 18644 14464
rect 20088 14436 20444 14464
rect 14792 14424 14798 14436
rect 12713 14399 12771 14405
rect 12713 14365 12725 14399
rect 12759 14365 12771 14399
rect 12713 14359 12771 14365
rect 12802 14356 12808 14408
rect 12860 14356 12866 14408
rect 12986 14356 12992 14408
rect 13044 14356 13050 14408
rect 13265 14399 13323 14405
rect 13265 14365 13277 14399
rect 13311 14365 13323 14399
rect 13265 14359 13323 14365
rect 10245 14291 10303 14297
rect 10336 14300 10824 14328
rect 1762 14220 1768 14272
rect 1820 14260 1826 14272
rect 2133 14263 2191 14269
rect 2133 14260 2145 14263
rect 1820 14232 2145 14260
rect 1820 14220 1826 14232
rect 2133 14229 2145 14232
rect 2179 14229 2191 14263
rect 2133 14223 2191 14229
rect 2222 14220 2228 14272
rect 2280 14260 2286 14272
rect 2961 14263 3019 14269
rect 2961 14260 2973 14263
rect 2280 14232 2973 14260
rect 2280 14220 2286 14232
rect 2961 14229 2973 14232
rect 3007 14229 3019 14263
rect 2961 14223 3019 14229
rect 3789 14263 3847 14269
rect 3789 14229 3801 14263
rect 3835 14260 3847 14263
rect 3878 14260 3884 14272
rect 3835 14232 3884 14260
rect 3835 14229 3847 14232
rect 3789 14223 3847 14229
rect 3878 14220 3884 14232
rect 3936 14220 3942 14272
rect 4798 14220 4804 14272
rect 4856 14260 4862 14272
rect 5442 14260 5448 14272
rect 4856 14232 5448 14260
rect 4856 14220 4862 14232
rect 5442 14220 5448 14232
rect 5500 14260 5506 14272
rect 5626 14260 5632 14272
rect 5500 14232 5632 14260
rect 5500 14220 5506 14232
rect 5626 14220 5632 14232
rect 5684 14220 5690 14272
rect 8202 14220 8208 14272
rect 8260 14220 8266 14272
rect 9490 14220 9496 14272
rect 9548 14220 9554 14272
rect 10060 14260 10088 14288
rect 10336 14260 10364 14300
rect 12342 14288 12348 14340
rect 12400 14328 12406 14340
rect 13280 14328 13308 14359
rect 15010 14356 15016 14408
rect 15068 14356 15074 14408
rect 15197 14399 15255 14405
rect 15197 14365 15209 14399
rect 15243 14396 15255 14399
rect 15838 14396 15844 14408
rect 15243 14368 15844 14396
rect 15243 14365 15255 14368
rect 15197 14359 15255 14365
rect 15212 14328 15240 14359
rect 15838 14356 15844 14368
rect 15896 14356 15902 14408
rect 16209 14399 16267 14405
rect 16209 14365 16221 14399
rect 16255 14365 16267 14399
rect 16209 14359 16267 14365
rect 16301 14399 16359 14405
rect 16301 14365 16313 14399
rect 16347 14396 16359 14399
rect 16666 14396 16672 14408
rect 16347 14368 16672 14396
rect 16347 14365 16359 14368
rect 16301 14359 16359 14365
rect 12400 14300 13308 14328
rect 13832 14300 15240 14328
rect 16224 14328 16252 14359
rect 16666 14356 16672 14368
rect 16724 14356 16730 14408
rect 18340 14405 18368 14436
rect 18616 14408 18644 14436
rect 20438 14424 20444 14436
rect 20496 14424 20502 14476
rect 20622 14424 20628 14476
rect 20680 14464 20686 14476
rect 23477 14467 23535 14473
rect 20680 14436 21864 14464
rect 20680 14424 20686 14436
rect 18049 14399 18107 14405
rect 18049 14365 18061 14399
rect 18095 14365 18107 14399
rect 18049 14359 18107 14365
rect 18325 14399 18383 14405
rect 18325 14365 18337 14399
rect 18371 14365 18383 14399
rect 18325 14359 18383 14365
rect 17586 14328 17592 14340
rect 16224 14300 17592 14328
rect 12400 14288 12406 14300
rect 10060 14232 10364 14260
rect 10410 14220 10416 14272
rect 10468 14220 10474 14272
rect 10686 14220 10692 14272
rect 10744 14260 10750 14272
rect 13832 14260 13860 14300
rect 17586 14288 17592 14300
rect 17644 14288 17650 14340
rect 18064 14328 18092 14359
rect 18414 14356 18420 14408
rect 18472 14356 18478 14408
rect 18598 14356 18604 14408
rect 18656 14356 18662 14408
rect 20898 14356 20904 14408
rect 20956 14396 20962 14408
rect 21726 14396 21732 14408
rect 20956 14368 21732 14396
rect 20956 14356 20962 14368
rect 21726 14356 21732 14368
rect 21784 14356 21790 14408
rect 21836 14405 21864 14436
rect 23477 14433 23489 14467
rect 23523 14464 23535 14467
rect 23934 14464 23940 14476
rect 23523 14436 23940 14464
rect 23523 14433 23535 14436
rect 23477 14427 23535 14433
rect 23934 14424 23940 14436
rect 23992 14464 23998 14476
rect 23992 14436 24440 14464
rect 23992 14424 23998 14436
rect 21821 14399 21879 14405
rect 21821 14365 21833 14399
rect 21867 14365 21879 14399
rect 21821 14359 21879 14365
rect 22278 14356 22284 14408
rect 22336 14356 22342 14408
rect 22465 14399 22523 14405
rect 22465 14365 22477 14399
rect 22511 14396 22523 14399
rect 22554 14396 22560 14408
rect 22511 14368 22560 14396
rect 22511 14365 22523 14368
rect 22465 14359 22523 14365
rect 22554 14356 22560 14368
rect 22612 14356 22618 14408
rect 24412 14405 24440 14436
rect 24397 14399 24455 14405
rect 24397 14365 24409 14399
rect 24443 14365 24455 14399
rect 24397 14359 24455 14365
rect 24581 14399 24639 14405
rect 24581 14365 24593 14399
rect 24627 14365 24639 14399
rect 24581 14359 24639 14365
rect 20346 14328 20352 14340
rect 18064 14300 20352 14328
rect 20346 14288 20352 14300
rect 20404 14288 20410 14340
rect 21744 14328 21772 14356
rect 22002 14328 22008 14340
rect 21744 14300 22008 14328
rect 22002 14288 22008 14300
rect 22060 14288 22066 14340
rect 22830 14288 22836 14340
rect 22888 14328 22894 14340
rect 23017 14331 23075 14337
rect 23017 14328 23029 14331
rect 22888 14300 23029 14328
rect 22888 14288 22894 14300
rect 23017 14297 23029 14300
rect 23063 14297 23075 14331
rect 23017 14291 23075 14297
rect 23198 14288 23204 14340
rect 23256 14328 23262 14340
rect 24596 14328 24624 14359
rect 26602 14356 26608 14408
rect 26660 14356 26666 14408
rect 26694 14356 26700 14408
rect 26752 14356 26758 14408
rect 23256 14300 24624 14328
rect 23256 14288 23262 14300
rect 10744 14232 13860 14260
rect 13909 14263 13967 14269
rect 10744 14220 10750 14232
rect 13909 14229 13921 14263
rect 13955 14260 13967 14263
rect 14274 14260 14280 14272
rect 13955 14232 14280 14260
rect 13955 14229 13967 14232
rect 13909 14223 13967 14229
rect 14274 14220 14280 14232
rect 14332 14220 14338 14272
rect 16022 14220 16028 14272
rect 16080 14220 16086 14272
rect 16669 14263 16727 14269
rect 16669 14229 16681 14263
rect 16715 14260 16727 14263
rect 18138 14260 18144 14272
rect 16715 14232 18144 14260
rect 16715 14229 16727 14232
rect 16669 14223 16727 14229
rect 18138 14220 18144 14232
rect 18196 14220 18202 14272
rect 18230 14220 18236 14272
rect 18288 14260 18294 14272
rect 18874 14260 18880 14272
rect 18288 14232 18880 14260
rect 18288 14220 18294 14232
rect 18874 14220 18880 14232
rect 18932 14260 18938 14272
rect 20806 14260 20812 14272
rect 18932 14232 20812 14260
rect 18932 14220 18938 14232
rect 20806 14220 20812 14232
rect 20864 14220 20870 14272
rect 21174 14220 21180 14272
rect 21232 14260 21238 14272
rect 21453 14263 21511 14269
rect 21453 14260 21465 14263
rect 21232 14232 21465 14260
rect 21232 14220 21238 14232
rect 21453 14229 21465 14232
rect 21499 14229 21511 14263
rect 21453 14223 21511 14229
rect 24118 14220 24124 14272
rect 24176 14260 24182 14272
rect 26053 14263 26111 14269
rect 26053 14260 26065 14263
rect 24176 14232 26065 14260
rect 24176 14220 24182 14232
rect 26053 14229 26065 14232
rect 26099 14229 26111 14263
rect 26053 14223 26111 14229
rect 1104 14170 27876 14192
rect 1104 14118 4874 14170
rect 4926 14118 4938 14170
rect 4990 14118 5002 14170
rect 5054 14118 5066 14170
rect 5118 14118 5130 14170
rect 5182 14118 27876 14170
rect 1104 14096 27876 14118
rect 1574 14059 1632 14065
rect 1574 14025 1586 14059
rect 1620 14056 1632 14059
rect 2130 14056 2136 14068
rect 1620 14028 2136 14056
rect 1620 14025 1632 14028
rect 1574 14019 1632 14025
rect 2130 14016 2136 14028
rect 2188 14016 2194 14068
rect 2317 14059 2375 14065
rect 2317 14025 2329 14059
rect 2363 14025 2375 14059
rect 2317 14019 2375 14025
rect 3973 14059 4031 14065
rect 3973 14025 3985 14059
rect 4019 14056 4031 14059
rect 4019 14028 4660 14056
rect 4019 14025 4031 14028
rect 3973 14019 4031 14025
rect 2041 13991 2099 13997
rect 2041 13957 2053 13991
rect 2087 13988 2099 13991
rect 2222 13988 2228 14000
rect 2087 13960 2228 13988
rect 2087 13957 2099 13960
rect 2041 13951 2099 13957
rect 2222 13948 2228 13960
rect 2280 13948 2286 14000
rect 2332 13988 2360 14019
rect 2654 13991 2712 13997
rect 2654 13988 2666 13991
rect 2332 13960 2666 13988
rect 2654 13957 2666 13960
rect 2700 13957 2712 13991
rect 2654 13951 2712 13957
rect 4062 13948 4068 14000
rect 4120 13988 4126 14000
rect 4120 13960 4384 13988
rect 4120 13948 4126 13960
rect 1394 13880 1400 13932
rect 1452 13880 1458 13932
rect 1486 13880 1492 13932
rect 1544 13880 1550 13932
rect 1670 13880 1676 13932
rect 1728 13880 1734 13932
rect 1762 13880 1768 13932
rect 1820 13880 1826 13932
rect 1949 13923 2007 13929
rect 1949 13889 1961 13923
rect 1995 13889 2007 13923
rect 1949 13883 2007 13889
rect 2133 13923 2191 13929
rect 2133 13889 2145 13923
rect 2179 13920 2191 13923
rect 2314 13920 2320 13932
rect 2179 13892 2320 13920
rect 2179 13889 2191 13892
rect 2133 13883 2191 13889
rect 1964 13852 1992 13883
rect 2314 13880 2320 13892
rect 2372 13880 2378 13932
rect 4356 13929 4384 13960
rect 4248 13923 4306 13929
rect 4248 13889 4260 13923
rect 4294 13889 4306 13923
rect 4248 13883 4306 13889
rect 4341 13923 4399 13929
rect 4341 13889 4353 13923
rect 4387 13920 4399 13923
rect 4433 13923 4491 13929
rect 4433 13920 4445 13923
rect 4387 13892 4445 13920
rect 4387 13889 4399 13892
rect 4341 13883 4399 13889
rect 4433 13889 4445 13892
rect 4479 13889 4491 13923
rect 4632 13920 4660 14028
rect 4706 14016 4712 14068
rect 4764 14056 4770 14068
rect 4985 14059 5043 14065
rect 4985 14056 4997 14059
rect 4764 14028 4997 14056
rect 4764 14016 4770 14028
rect 4985 14025 4997 14028
rect 5031 14025 5043 14059
rect 5902 14056 5908 14068
rect 4985 14019 5043 14025
rect 5184 14028 5908 14056
rect 4798 13948 4804 14000
rect 4856 13948 4862 14000
rect 5184 13920 5212 14028
rect 5902 14016 5908 14028
rect 5960 14016 5966 14068
rect 6362 14016 6368 14068
rect 6420 14016 6426 14068
rect 7650 14016 7656 14068
rect 7708 14056 7714 14068
rect 7745 14059 7803 14065
rect 7745 14056 7757 14059
rect 7708 14028 7757 14056
rect 7708 14016 7714 14028
rect 7745 14025 7757 14028
rect 7791 14025 7803 14059
rect 8570 14056 8576 14068
rect 7745 14019 7803 14025
rect 8404 14028 8576 14056
rect 8404 13997 8432 14028
rect 8570 14016 8576 14028
rect 8628 14056 8634 14068
rect 11885 14059 11943 14065
rect 11885 14056 11897 14059
rect 8628 14028 11897 14056
rect 8628 14016 8634 14028
rect 11885 14025 11897 14028
rect 11931 14056 11943 14059
rect 16143 14059 16201 14065
rect 11931 14028 14596 14056
rect 11931 14025 11943 14028
rect 11885 14019 11943 14025
rect 7009 13991 7067 13997
rect 7009 13988 7021 13991
rect 4632 13892 5212 13920
rect 5828 13960 7021 13988
rect 5828 13906 5856 13960
rect 7009 13957 7021 13960
rect 7055 13957 7067 13991
rect 8173 13991 8231 13997
rect 8173 13988 8185 13991
rect 7009 13951 7067 13957
rect 7668 13960 8185 13988
rect 7668 13932 7696 13960
rect 8173 13957 8185 13960
rect 8219 13957 8231 13991
rect 8389 13991 8447 13997
rect 8389 13988 8401 13991
rect 8173 13951 8231 13957
rect 8312 13960 8401 13988
rect 4433 13883 4491 13889
rect 2038 13852 2044 13864
rect 1964 13824 2044 13852
rect 2038 13812 2044 13824
rect 2096 13812 2102 13864
rect 2406 13812 2412 13864
rect 2464 13812 2470 13864
rect 4264 13852 4292 13883
rect 7650 13880 7656 13932
rect 7708 13880 7714 13932
rect 7929 13923 7987 13929
rect 7929 13889 7941 13923
rect 7975 13920 7987 13923
rect 8312 13920 8340 13960
rect 8389 13957 8401 13960
rect 8435 13957 8447 13991
rect 8389 13951 8447 13957
rect 9766 13948 9772 14000
rect 9824 13988 9830 14000
rect 10686 13988 10692 14000
rect 9824 13960 10692 13988
rect 9824 13948 9830 13960
rect 10060 13929 10088 13960
rect 10686 13948 10692 13960
rect 10744 13948 10750 14000
rect 13296 13991 13354 13997
rect 13296 13957 13308 13991
rect 13342 13988 13354 13991
rect 13633 13991 13691 13997
rect 13633 13988 13645 13991
rect 13342 13960 13645 13988
rect 13342 13957 13354 13960
rect 13296 13951 13354 13957
rect 13633 13957 13645 13960
rect 13679 13957 13691 13991
rect 13633 13951 13691 13957
rect 13722 13948 13728 14000
rect 13780 13988 13786 14000
rect 14001 13991 14059 13997
rect 14001 13988 14013 13991
rect 13780 13960 14013 13988
rect 13780 13948 13786 13960
rect 14001 13957 14013 13960
rect 14047 13957 14059 13991
rect 14001 13951 14059 13957
rect 14090 13948 14096 14000
rect 14148 13997 14154 14000
rect 14148 13991 14177 13997
rect 14165 13957 14177 13991
rect 14568 13988 14596 14028
rect 16143 14025 16155 14059
rect 16189 14056 16201 14059
rect 16758 14056 16764 14068
rect 16189 14028 16764 14056
rect 16189 14025 16201 14028
rect 16143 14019 16201 14025
rect 16758 14016 16764 14028
rect 16816 14016 16822 14068
rect 17954 14056 17960 14068
rect 17512 14028 17960 14056
rect 15933 13991 15991 13997
rect 14568 13960 14688 13988
rect 14148 13951 14177 13957
rect 14148 13948 14154 13951
rect 7975 13892 8340 13920
rect 10045 13923 10103 13929
rect 7975 13889 7987 13892
rect 7929 13883 7987 13889
rect 10045 13889 10057 13923
rect 10091 13889 10103 13923
rect 10045 13883 10103 13889
rect 10321 13923 10379 13929
rect 10321 13889 10333 13923
rect 10367 13889 10379 13923
rect 10321 13883 10379 13889
rect 4614 13852 4620 13864
rect 4264 13824 4620 13852
rect 4614 13812 4620 13824
rect 4672 13812 4678 13864
rect 5353 13855 5411 13861
rect 5353 13821 5365 13855
rect 5399 13852 5411 13855
rect 5626 13852 5632 13864
rect 5399 13824 5632 13852
rect 5399 13821 5411 13824
rect 5353 13815 5411 13821
rect 5626 13812 5632 13824
rect 5684 13812 5690 13864
rect 6086 13812 6092 13864
rect 6144 13812 6150 13864
rect 6687 13855 6745 13861
rect 6687 13852 6699 13855
rect 6196 13824 6699 13852
rect 5534 13744 5540 13796
rect 5592 13784 5598 13796
rect 6196 13784 6224 13824
rect 6687 13821 6699 13824
rect 6733 13821 6745 13855
rect 6687 13815 6745 13821
rect 6825 13855 6883 13861
rect 6825 13821 6837 13855
rect 6871 13852 6883 13855
rect 6914 13852 6920 13864
rect 6871 13824 6920 13852
rect 6871 13821 6883 13824
rect 6825 13815 6883 13821
rect 6914 13812 6920 13824
rect 6972 13812 6978 13864
rect 9769 13855 9827 13861
rect 9769 13821 9781 13855
rect 9815 13852 9827 13855
rect 9858 13852 9864 13864
rect 9815 13824 9864 13852
rect 9815 13821 9827 13824
rect 9769 13815 9827 13821
rect 9858 13812 9864 13824
rect 9916 13852 9922 13864
rect 10336 13852 10364 13883
rect 10502 13880 10508 13932
rect 10560 13880 10566 13932
rect 11977 13923 12035 13929
rect 11977 13889 11989 13923
rect 12023 13920 12035 13923
rect 12342 13920 12348 13932
rect 12023 13892 12348 13920
rect 12023 13889 12035 13892
rect 11977 13883 12035 13889
rect 10594 13852 10600 13864
rect 9916 13824 10272 13852
rect 10336 13824 10600 13852
rect 9916 13812 9922 13824
rect 5592 13756 6224 13784
rect 5592 13744 5598 13756
rect 7190 13744 7196 13796
rect 7248 13784 7254 13796
rect 7834 13784 7840 13796
rect 7248 13756 7840 13784
rect 7248 13744 7254 13756
rect 7834 13744 7840 13756
rect 7892 13784 7898 13796
rect 8754 13784 8760 13796
rect 7892 13756 8760 13784
rect 7892 13744 7898 13756
rect 8754 13744 8760 13756
rect 8812 13744 8818 13796
rect 10134 13784 10140 13796
rect 8864 13756 10140 13784
rect 1670 13676 1676 13728
rect 1728 13716 1734 13728
rect 3602 13716 3608 13728
rect 1728 13688 3608 13716
rect 1728 13676 1734 13688
rect 3602 13676 3608 13688
rect 3660 13716 3666 13728
rect 3789 13719 3847 13725
rect 3789 13716 3801 13719
rect 3660 13688 3801 13716
rect 3660 13676 3666 13688
rect 3789 13685 3801 13688
rect 3835 13716 3847 13719
rect 3970 13716 3976 13728
rect 3835 13688 3976 13716
rect 3835 13685 3847 13688
rect 3789 13679 3847 13685
rect 3970 13676 3976 13688
rect 4028 13676 4034 13728
rect 4614 13676 4620 13728
rect 4672 13716 4678 13728
rect 4801 13719 4859 13725
rect 4801 13716 4813 13719
rect 4672 13688 4813 13716
rect 4672 13676 4678 13688
rect 4801 13685 4813 13688
rect 4847 13685 4859 13719
rect 4801 13679 4859 13685
rect 7926 13676 7932 13728
rect 7984 13676 7990 13728
rect 8018 13676 8024 13728
rect 8076 13676 8082 13728
rect 8205 13719 8263 13725
rect 8205 13685 8217 13719
rect 8251 13716 8263 13719
rect 8864 13716 8892 13756
rect 10134 13744 10140 13756
rect 10192 13744 10198 13796
rect 10244 13784 10272 13824
rect 10594 13812 10600 13824
rect 10652 13812 10658 13864
rect 11054 13852 11060 13864
rect 10704 13824 11060 13852
rect 10704 13784 10732 13824
rect 11054 13812 11060 13824
rect 11112 13812 11118 13864
rect 12176 13793 12204 13892
rect 12342 13880 12348 13892
rect 12400 13880 12406 13932
rect 13446 13880 13452 13932
rect 13504 13920 13510 13932
rect 13541 13923 13599 13929
rect 13541 13920 13553 13923
rect 13504 13892 13553 13920
rect 13504 13880 13510 13892
rect 13541 13889 13553 13892
rect 13587 13889 13599 13923
rect 13541 13883 13599 13889
rect 13814 13880 13820 13932
rect 13872 13880 13878 13932
rect 13906 13880 13912 13932
rect 13964 13880 13970 13932
rect 14274 13880 14280 13932
rect 14332 13880 14338 13932
rect 14550 13880 14556 13932
rect 14608 13880 14614 13932
rect 14660 13929 14688 13960
rect 15933 13957 15945 13991
rect 15979 13988 15991 13991
rect 16298 13988 16304 14000
rect 15979 13960 16304 13988
rect 15979 13957 15991 13960
rect 15933 13951 15991 13957
rect 16298 13948 16304 13960
rect 16356 13948 16362 14000
rect 14645 13923 14703 13929
rect 14645 13889 14657 13923
rect 14691 13889 14703 13923
rect 14645 13883 14703 13889
rect 17218 13880 17224 13932
rect 17276 13880 17282 13932
rect 17512 13929 17540 14028
rect 17954 14016 17960 14028
rect 18012 14016 18018 14068
rect 18598 14016 18604 14068
rect 18656 14056 18662 14068
rect 19613 14059 19671 14065
rect 19613 14056 19625 14059
rect 18656 14028 19625 14056
rect 18656 14016 18662 14028
rect 19613 14025 19625 14028
rect 19659 14025 19671 14059
rect 20714 14056 20720 14068
rect 19613 14019 19671 14025
rect 20272 14028 20720 14056
rect 19334 13988 19340 14000
rect 17972 13960 19340 13988
rect 17497 13923 17555 13929
rect 17497 13889 17509 13923
rect 17543 13889 17555 13923
rect 17497 13883 17555 13889
rect 17586 13880 17592 13932
rect 17644 13880 17650 13932
rect 17681 13923 17739 13929
rect 17681 13889 17693 13923
rect 17727 13920 17739 13923
rect 17770 13920 17776 13932
rect 17727 13892 17776 13920
rect 17727 13889 17739 13892
rect 17681 13883 17739 13889
rect 17770 13880 17776 13892
rect 17828 13880 17834 13932
rect 17972 13929 18000 13960
rect 17865 13923 17923 13929
rect 17865 13889 17877 13923
rect 17911 13920 17923 13923
rect 17957 13923 18015 13929
rect 17957 13920 17969 13923
rect 17911 13892 17969 13920
rect 17911 13889 17923 13892
rect 17865 13883 17923 13889
rect 17957 13889 17969 13892
rect 18003 13889 18015 13923
rect 17957 13883 18015 13889
rect 18049 13923 18107 13929
rect 18049 13889 18061 13923
rect 18095 13920 18107 13923
rect 18138 13920 18144 13932
rect 18095 13892 18144 13920
rect 18095 13889 18107 13892
rect 18049 13883 18107 13889
rect 18138 13880 18144 13892
rect 18196 13880 18202 13932
rect 19076 13929 19104 13960
rect 19334 13948 19340 13960
rect 19392 13948 19398 14000
rect 19705 13991 19763 13997
rect 18233 13923 18291 13929
rect 18233 13889 18245 13923
rect 18279 13889 18291 13923
rect 18233 13883 18291 13889
rect 19061 13923 19119 13929
rect 19061 13889 19073 13923
rect 19107 13889 19119 13923
rect 19061 13883 19119 13889
rect 17604 13852 17632 13880
rect 18248 13852 18276 13883
rect 19150 13880 19156 13932
rect 19208 13880 19214 13932
rect 19426 13914 19432 13966
rect 19484 13914 19490 13966
rect 19705 13957 19717 13991
rect 19751 13988 19763 13991
rect 19886 13988 19892 14000
rect 19751 13960 19892 13988
rect 19751 13957 19763 13960
rect 19705 13951 19763 13957
rect 19886 13948 19892 13960
rect 19944 13988 19950 14000
rect 20272 13988 20300 14028
rect 20714 14016 20720 14028
rect 20772 14016 20778 14068
rect 20990 14016 20996 14068
rect 21048 14056 21054 14068
rect 21361 14059 21419 14065
rect 21361 14056 21373 14059
rect 21048 14028 21373 14056
rect 21048 14016 21054 14028
rect 21361 14025 21373 14028
rect 21407 14056 21419 14059
rect 21542 14056 21548 14068
rect 21407 14028 21548 14056
rect 21407 14025 21419 14028
rect 21361 14019 21419 14025
rect 21542 14016 21548 14028
rect 21600 14016 21606 14068
rect 22554 14016 22560 14068
rect 22612 14016 22618 14068
rect 26237 14059 26295 14065
rect 26237 14056 26249 14059
rect 22664 14028 26249 14056
rect 22664 13988 22692 14028
rect 26237 14025 26249 14028
rect 26283 14025 26295 14059
rect 26237 14019 26295 14025
rect 26602 14016 26608 14068
rect 26660 14056 26666 14068
rect 26697 14059 26755 14065
rect 26697 14056 26709 14059
rect 26660 14028 26709 14056
rect 26660 14016 26666 14028
rect 26697 14025 26709 14028
rect 26743 14025 26755 14059
rect 26697 14019 26755 14025
rect 19944 13960 20300 13988
rect 21100 13960 22692 13988
rect 19944 13948 19950 13960
rect 19521 13926 19579 13929
rect 19610 13926 19616 13932
rect 19521 13923 19616 13926
rect 19521 13889 19533 13923
rect 19567 13898 19616 13923
rect 19567 13889 19579 13898
rect 19521 13883 19579 13889
rect 19610 13880 19616 13898
rect 19668 13880 19674 13932
rect 20073 13923 20131 13929
rect 19781 13913 19839 13919
rect 19781 13910 19793 13913
rect 19720 13882 19793 13910
rect 19245 13855 19303 13861
rect 17604 13824 19196 13852
rect 10244 13756 10732 13784
rect 12161 13787 12219 13793
rect 12161 13753 12173 13787
rect 12207 13753 12219 13787
rect 16945 13787 17003 13793
rect 16945 13784 16957 13787
rect 12161 13747 12219 13753
rect 14134 13756 16957 13784
rect 8251 13688 8892 13716
rect 8251 13685 8263 13688
rect 8205 13679 8263 13685
rect 9122 13676 9128 13728
rect 9180 13716 9186 13728
rect 9493 13719 9551 13725
rect 9493 13716 9505 13719
rect 9180 13688 9505 13716
rect 9180 13676 9186 13688
rect 9493 13685 9505 13688
rect 9539 13685 9551 13719
rect 9493 13679 9551 13685
rect 9953 13719 10011 13725
rect 9953 13685 9965 13719
rect 9999 13716 10011 13719
rect 10318 13716 10324 13728
rect 9999 13688 10324 13716
rect 9999 13685 10011 13688
rect 9953 13679 10011 13685
rect 10318 13676 10324 13688
rect 10376 13676 10382 13728
rect 13906 13676 13912 13728
rect 13964 13716 13970 13728
rect 14134 13716 14162 13756
rect 16945 13753 16957 13756
rect 16991 13753 17003 13787
rect 19168 13784 19196 13824
rect 19245 13821 19257 13855
rect 19291 13852 19303 13855
rect 19426 13852 19432 13864
rect 19291 13824 19432 13852
rect 19291 13821 19303 13824
rect 19245 13815 19303 13821
rect 19426 13812 19432 13824
rect 19484 13812 19490 13864
rect 19334 13784 19340 13796
rect 19168 13756 19340 13784
rect 16945 13747 17003 13753
rect 19334 13744 19340 13756
rect 19392 13744 19398 13796
rect 19518 13744 19524 13796
rect 19576 13744 19582 13796
rect 19720 13784 19748 13882
rect 19781 13879 19793 13882
rect 19827 13879 19839 13913
rect 20073 13889 20085 13923
rect 20119 13920 20131 13923
rect 20162 13920 20168 13932
rect 20119 13892 20168 13920
rect 20119 13889 20131 13892
rect 20073 13883 20131 13889
rect 20162 13880 20168 13892
rect 20220 13880 20226 13932
rect 20346 13880 20352 13932
rect 20404 13929 20410 13932
rect 20404 13920 20415 13929
rect 21100 13920 21128 13960
rect 22922 13948 22928 14000
rect 22980 13988 22986 14000
rect 23201 13991 23259 13997
rect 23201 13988 23213 13991
rect 22980 13960 23213 13988
rect 22980 13948 22986 13960
rect 23201 13957 23213 13960
rect 23247 13988 23259 13991
rect 25133 13991 25191 13997
rect 25133 13988 25145 13991
rect 23247 13960 25145 13988
rect 23247 13957 23259 13960
rect 23201 13951 23259 13957
rect 25133 13957 25145 13960
rect 25179 13957 25191 13991
rect 26620 13988 26648 14016
rect 25133 13951 25191 13957
rect 26068 13960 26648 13988
rect 20404 13892 21128 13920
rect 20404 13883 20415 13892
rect 20404 13880 20410 13883
rect 21174 13880 21180 13932
rect 21232 13880 21238 13932
rect 21450 13880 21456 13932
rect 21508 13880 21514 13932
rect 22741 13923 22799 13929
rect 22741 13889 22753 13923
rect 22787 13889 22799 13923
rect 22741 13883 22799 13889
rect 19781 13873 19839 13879
rect 22756 13852 22784 13883
rect 23014 13880 23020 13932
rect 23072 13880 23078 13932
rect 23109 13923 23167 13929
rect 23109 13889 23121 13923
rect 23155 13889 23167 13923
rect 23109 13883 23167 13889
rect 23124 13852 23152 13883
rect 23382 13880 23388 13932
rect 23440 13880 23446 13932
rect 25038 13880 25044 13932
rect 25096 13880 25102 13932
rect 25222 13880 25228 13932
rect 25280 13880 25286 13932
rect 26068 13929 26096 13960
rect 26053 13923 26111 13929
rect 26053 13889 26065 13923
rect 26099 13889 26111 13923
rect 26053 13883 26111 13889
rect 26418 13880 26424 13932
rect 26476 13920 26482 13932
rect 26513 13923 26571 13929
rect 26513 13920 26525 13923
rect 26476 13892 26525 13920
rect 26476 13880 26482 13892
rect 26513 13889 26525 13892
rect 26559 13889 26571 13923
rect 26513 13883 26571 13889
rect 23290 13852 23296 13864
rect 22756 13824 23296 13852
rect 23290 13812 23296 13824
rect 23348 13812 23354 13864
rect 19794 13784 19800 13796
rect 19720 13756 19800 13784
rect 19794 13744 19800 13756
rect 19852 13784 19858 13796
rect 19981 13787 20039 13793
rect 19981 13784 19993 13787
rect 19852 13756 19993 13784
rect 19852 13744 19858 13756
rect 19981 13753 19993 13756
rect 20027 13753 20039 13787
rect 20257 13787 20315 13793
rect 20257 13784 20269 13787
rect 19981 13747 20039 13753
rect 20088 13756 20269 13784
rect 13964 13688 14162 13716
rect 13964 13676 13970 13688
rect 14366 13676 14372 13728
rect 14424 13676 14430 13728
rect 15838 13676 15844 13728
rect 15896 13716 15902 13728
rect 16117 13719 16175 13725
rect 16117 13716 16129 13719
rect 15896 13688 16129 13716
rect 15896 13676 15902 13688
rect 16117 13685 16129 13688
rect 16163 13685 16175 13719
rect 16117 13679 16175 13685
rect 16298 13676 16304 13728
rect 16356 13676 16362 13728
rect 17405 13719 17463 13725
rect 17405 13685 17417 13719
rect 17451 13716 17463 13719
rect 17865 13719 17923 13725
rect 17865 13716 17877 13719
rect 17451 13688 17877 13716
rect 17451 13685 17463 13688
rect 17405 13679 17463 13685
rect 17865 13685 17877 13688
rect 17911 13685 17923 13719
rect 17865 13679 17923 13685
rect 19426 13676 19432 13728
rect 19484 13676 19490 13728
rect 19536 13716 19564 13744
rect 20088 13716 20116 13756
rect 20257 13753 20269 13756
rect 20303 13753 20315 13787
rect 20257 13747 20315 13753
rect 22278 13744 22284 13796
rect 22336 13784 22342 13796
rect 23109 13787 23167 13793
rect 23109 13784 23121 13787
rect 22336 13756 23121 13784
rect 22336 13744 22342 13756
rect 23109 13753 23121 13756
rect 23155 13753 23167 13787
rect 23400 13784 23428 13880
rect 25056 13852 25084 13880
rect 25406 13852 25412 13864
rect 25056 13824 25412 13852
rect 25406 13812 25412 13824
rect 25464 13812 25470 13864
rect 25590 13812 25596 13864
rect 25648 13812 25654 13864
rect 25961 13855 26019 13861
rect 25961 13821 25973 13855
rect 26007 13852 26019 13855
rect 26234 13852 26240 13864
rect 26007 13824 26240 13852
rect 26007 13821 26019 13824
rect 25961 13815 26019 13821
rect 26234 13812 26240 13824
rect 26292 13812 26298 13864
rect 26326 13812 26332 13864
rect 26384 13812 26390 13864
rect 25774 13784 25780 13796
rect 23400 13756 25780 13784
rect 23109 13747 23167 13753
rect 25774 13744 25780 13756
rect 25832 13784 25838 13796
rect 26436 13784 26464 13880
rect 25832 13756 26464 13784
rect 25832 13744 25838 13756
rect 19536 13688 20116 13716
rect 20162 13676 20168 13728
rect 20220 13716 20226 13728
rect 20993 13719 21051 13725
rect 20993 13716 21005 13719
rect 20220 13688 21005 13716
rect 20220 13676 20226 13688
rect 20993 13685 21005 13688
rect 21039 13685 21051 13719
rect 20993 13679 21051 13685
rect 21266 13676 21272 13728
rect 21324 13716 21330 13728
rect 26418 13716 26424 13728
rect 21324 13688 26424 13716
rect 21324 13676 21330 13688
rect 26418 13676 26424 13688
rect 26476 13676 26482 13728
rect 1104 13626 27876 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 27876 13626
rect 1104 13552 27876 13574
rect 1670 13472 1676 13524
rect 1728 13512 1734 13524
rect 2041 13515 2099 13521
rect 2041 13512 2053 13515
rect 1728 13484 2053 13512
rect 1728 13472 1734 13484
rect 2041 13481 2053 13484
rect 2087 13481 2099 13515
rect 2041 13475 2099 13481
rect 4157 13515 4215 13521
rect 4157 13481 4169 13515
rect 4203 13512 4215 13515
rect 5258 13512 5264 13524
rect 4203 13484 5264 13512
rect 4203 13481 4215 13484
rect 4157 13475 4215 13481
rect 5258 13472 5264 13484
rect 5316 13472 5322 13524
rect 7926 13472 7932 13524
rect 7984 13512 7990 13524
rect 8113 13515 8171 13521
rect 8113 13512 8125 13515
rect 7984 13484 8125 13512
rect 7984 13472 7990 13484
rect 8113 13481 8125 13484
rect 8159 13481 8171 13515
rect 8113 13475 8171 13481
rect 8205 13515 8263 13521
rect 8205 13481 8217 13515
rect 8251 13512 8263 13515
rect 8754 13512 8760 13524
rect 8251 13484 8760 13512
rect 8251 13481 8263 13484
rect 8205 13475 8263 13481
rect 8754 13472 8760 13484
rect 8812 13472 8818 13524
rect 11054 13472 11060 13524
rect 11112 13512 11118 13524
rect 11112 13484 11376 13512
rect 11112 13472 11118 13484
rect 1854 13404 1860 13456
rect 1912 13404 1918 13456
rect 5534 13404 5540 13456
rect 5592 13404 5598 13456
rect 7190 13404 7196 13456
rect 7248 13404 7254 13456
rect 5552 13376 5580 13404
rect 7944 13376 7972 13472
rect 8018 13404 8024 13456
rect 8076 13444 8082 13456
rect 8297 13447 8355 13453
rect 8297 13444 8309 13447
rect 8076 13416 8309 13444
rect 8076 13404 8082 13416
rect 8297 13413 8309 13416
rect 8343 13413 8355 13447
rect 8297 13407 8355 13413
rect 5459 13348 5580 13376
rect 7576 13348 7972 13376
rect 1486 13268 1492 13320
rect 1544 13308 1550 13320
rect 5459 13317 5487 13348
rect 3973 13311 4031 13317
rect 3973 13308 3985 13311
rect 1544 13280 2268 13308
rect 1544 13268 1550 13280
rect 1394 13200 1400 13252
rect 1452 13240 1458 13252
rect 2240 13249 2268 13280
rect 2792 13280 3985 13308
rect 2009 13243 2067 13249
rect 2009 13240 2021 13243
rect 1452 13212 2021 13240
rect 1452 13200 1458 13212
rect 2009 13209 2021 13212
rect 2055 13209 2067 13243
rect 2009 13203 2067 13209
rect 2225 13243 2283 13249
rect 2225 13209 2237 13243
rect 2271 13240 2283 13243
rect 2682 13240 2688 13252
rect 2271 13212 2688 13240
rect 2271 13209 2283 13212
rect 2225 13203 2283 13209
rect 2682 13200 2688 13212
rect 2740 13240 2746 13252
rect 2792 13240 2820 13280
rect 3973 13277 3985 13280
rect 4019 13277 4031 13311
rect 3973 13271 4031 13277
rect 5444 13311 5502 13317
rect 5444 13277 5456 13311
rect 5490 13277 5502 13311
rect 5444 13271 5502 13277
rect 5537 13311 5595 13317
rect 5537 13277 5549 13311
rect 5583 13308 5595 13311
rect 5626 13308 5632 13320
rect 5583 13280 5632 13308
rect 5583 13277 5595 13280
rect 5537 13271 5595 13277
rect 5626 13268 5632 13280
rect 5684 13268 5690 13320
rect 7576 13317 7604 13348
rect 7285 13311 7343 13317
rect 7285 13277 7297 13311
rect 7331 13308 7343 13311
rect 7561 13311 7619 13317
rect 7561 13308 7573 13311
rect 7331 13280 7573 13308
rect 7331 13277 7343 13280
rect 7285 13271 7343 13277
rect 7561 13277 7573 13280
rect 7607 13277 7619 13311
rect 7561 13271 7619 13277
rect 7745 13311 7803 13317
rect 7745 13277 7757 13311
rect 7791 13308 7803 13311
rect 8036 13308 8064 13404
rect 8404 13348 8984 13376
rect 8404 13317 8432 13348
rect 8956 13320 8984 13348
rect 10594 13336 10600 13388
rect 10652 13376 10658 13388
rect 11348 13385 11376 13484
rect 13814 13472 13820 13524
rect 13872 13512 13878 13524
rect 14185 13515 14243 13521
rect 14185 13512 14197 13515
rect 13872 13484 14197 13512
rect 13872 13472 13878 13484
rect 14185 13481 14197 13484
rect 14231 13481 14243 13515
rect 14185 13475 14243 13481
rect 14274 13472 14280 13524
rect 14332 13472 14338 13524
rect 16390 13512 16396 13524
rect 14936 13484 16396 13512
rect 10873 13379 10931 13385
rect 10873 13376 10885 13379
rect 10652 13348 10885 13376
rect 10652 13336 10658 13348
rect 10873 13345 10885 13348
rect 10919 13345 10931 13379
rect 10873 13339 10931 13345
rect 11333 13379 11391 13385
rect 11333 13345 11345 13379
rect 11379 13345 11391 13379
rect 11333 13339 11391 13345
rect 14093 13379 14151 13385
rect 14093 13345 14105 13379
rect 14139 13376 14151 13379
rect 14936 13376 14964 13484
rect 16390 13472 16396 13484
rect 16448 13472 16454 13524
rect 19610 13472 19616 13524
rect 19668 13512 19674 13524
rect 19797 13515 19855 13521
rect 19797 13512 19809 13515
rect 19668 13484 19809 13512
rect 19668 13472 19674 13484
rect 19797 13481 19809 13484
rect 19843 13512 19855 13515
rect 20993 13515 21051 13521
rect 20993 13512 21005 13515
rect 19843 13484 21005 13512
rect 19843 13481 19855 13484
rect 19797 13475 19855 13481
rect 20993 13481 21005 13484
rect 21039 13481 21051 13515
rect 20993 13475 21051 13481
rect 21085 13515 21143 13521
rect 21085 13481 21097 13515
rect 21131 13512 21143 13515
rect 21174 13512 21180 13524
rect 21131 13484 21180 13512
rect 21131 13481 21143 13484
rect 21085 13475 21143 13481
rect 21174 13472 21180 13484
rect 21232 13472 21238 13524
rect 22922 13472 22928 13524
rect 22980 13472 22986 13524
rect 24118 13472 24124 13524
rect 24176 13512 24182 13524
rect 24581 13515 24639 13521
rect 24581 13512 24593 13515
rect 24176 13484 24593 13512
rect 24176 13472 24182 13484
rect 24581 13481 24593 13484
rect 24627 13481 24639 13515
rect 24581 13475 24639 13481
rect 25590 13472 25596 13524
rect 25648 13512 25654 13524
rect 25685 13515 25743 13521
rect 25685 13512 25697 13515
rect 25648 13484 25697 13512
rect 25648 13472 25654 13484
rect 25685 13481 25697 13484
rect 25731 13481 25743 13515
rect 25685 13475 25743 13481
rect 15378 13404 15384 13456
rect 15436 13444 15442 13456
rect 20073 13447 20131 13453
rect 15436 13416 16160 13444
rect 15436 13404 15442 13416
rect 14139 13348 14964 13376
rect 14139 13345 14151 13348
rect 14093 13339 14151 13345
rect 7791 13280 8064 13308
rect 8389 13311 8447 13317
rect 7791 13277 7803 13280
rect 7745 13271 7803 13277
rect 8389 13277 8401 13311
rect 8435 13277 8447 13311
rect 8389 13271 8447 13277
rect 8573 13311 8631 13317
rect 8573 13277 8585 13311
rect 8619 13277 8631 13311
rect 8573 13271 8631 13277
rect 2740 13212 2820 13240
rect 3789 13243 3847 13249
rect 2740 13200 2746 13212
rect 3789 13209 3801 13243
rect 3835 13240 3847 13243
rect 7009 13243 7067 13249
rect 3835 13212 4016 13240
rect 3835 13209 3847 13212
rect 3789 13203 3847 13209
rect 3988 13184 4016 13212
rect 7009 13209 7021 13243
rect 7055 13240 7067 13243
rect 7760 13240 7788 13271
rect 7055 13212 7788 13240
rect 8588 13240 8616 13271
rect 8938 13268 8944 13320
rect 8996 13268 9002 13320
rect 9122 13268 9128 13320
rect 9180 13268 9186 13320
rect 9766 13268 9772 13320
rect 9824 13308 9830 13320
rect 10134 13308 10140 13320
rect 9824 13280 10140 13308
rect 9824 13268 9830 13280
rect 10134 13268 10140 13280
rect 10192 13268 10198 13320
rect 10318 13268 10324 13320
rect 10376 13268 10382 13320
rect 10502 13268 10508 13320
rect 10560 13308 10566 13320
rect 11149 13311 11207 13317
rect 11149 13308 11161 13311
rect 10560 13280 11161 13308
rect 10560 13268 10566 13280
rect 11149 13277 11161 13280
rect 11195 13308 11207 13311
rect 11425 13311 11483 13317
rect 11425 13308 11437 13311
rect 11195 13280 11437 13308
rect 11195 13277 11207 13280
rect 11149 13271 11207 13277
rect 11425 13277 11437 13280
rect 11471 13277 11483 13311
rect 11425 13271 11483 13277
rect 14366 13268 14372 13320
rect 14424 13268 14430 13320
rect 14550 13268 14556 13320
rect 14608 13308 14614 13320
rect 14936 13317 14964 13348
rect 15197 13379 15255 13385
rect 15197 13345 15209 13379
rect 15243 13376 15255 13379
rect 16022 13376 16028 13388
rect 15243 13348 16028 13376
rect 15243 13345 15255 13348
rect 15197 13339 15255 13345
rect 16022 13336 16028 13348
rect 16080 13336 16086 13388
rect 16132 13385 16160 13416
rect 20073 13413 20085 13447
rect 20119 13444 20131 13447
rect 20622 13444 20628 13456
rect 20119 13416 20628 13444
rect 20119 13413 20131 13416
rect 20073 13407 20131 13413
rect 20622 13404 20628 13416
rect 20680 13404 20686 13456
rect 21266 13444 21272 13456
rect 20916 13416 21272 13444
rect 16117 13379 16175 13385
rect 16117 13345 16129 13379
rect 16163 13345 16175 13379
rect 16117 13339 16175 13345
rect 19245 13379 19303 13385
rect 19245 13345 19257 13379
rect 19291 13376 19303 13379
rect 19334 13376 19340 13388
rect 19291 13348 19340 13376
rect 19291 13345 19303 13348
rect 19245 13339 19303 13345
rect 19334 13336 19340 13348
rect 19392 13336 19398 13388
rect 19426 13336 19432 13388
rect 19484 13376 19490 13388
rect 20254 13376 20260 13388
rect 19484 13348 20260 13376
rect 19484 13336 19490 13348
rect 20254 13336 20260 13348
rect 20312 13336 20318 13388
rect 20346 13336 20352 13388
rect 20404 13376 20410 13388
rect 20717 13379 20775 13385
rect 20717 13376 20729 13379
rect 20404 13348 20729 13376
rect 20404 13336 20410 13348
rect 20717 13345 20729 13348
rect 20763 13345 20775 13379
rect 20717 13339 20775 13345
rect 14737 13311 14795 13317
rect 14737 13308 14749 13311
rect 14608 13280 14749 13308
rect 14608 13268 14614 13280
rect 14737 13277 14749 13280
rect 14783 13277 14795 13311
rect 14737 13271 14795 13277
rect 14921 13311 14979 13317
rect 14921 13277 14933 13311
rect 14967 13277 14979 13311
rect 14921 13271 14979 13277
rect 9140 13240 9168 13268
rect 8588 13212 9168 13240
rect 7055 13209 7067 13212
rect 7009 13203 7067 13209
rect 3970 13132 3976 13184
rect 4028 13132 4034 13184
rect 5169 13175 5227 13181
rect 5169 13141 5181 13175
rect 5215 13172 5227 13175
rect 5258 13172 5264 13184
rect 5215 13144 5264 13172
rect 5215 13141 5227 13144
rect 5169 13135 5227 13141
rect 5258 13132 5264 13144
rect 5316 13132 5322 13184
rect 7282 13132 7288 13184
rect 7340 13132 7346 13184
rect 7650 13132 7656 13184
rect 7708 13132 7714 13184
rect 7837 13175 7895 13181
rect 7837 13141 7849 13175
rect 7883 13172 7895 13175
rect 8110 13172 8116 13184
rect 7883 13144 8116 13172
rect 7883 13141 7895 13144
rect 7837 13135 7895 13141
rect 8110 13132 8116 13144
rect 8168 13132 8174 13184
rect 9030 13132 9036 13184
rect 9088 13132 9094 13184
rect 10134 13132 10140 13184
rect 10192 13132 10198 13184
rect 10686 13132 10692 13184
rect 10744 13172 10750 13184
rect 10873 13175 10931 13181
rect 10873 13172 10885 13175
rect 10744 13144 10885 13172
rect 10744 13132 10750 13144
rect 10873 13141 10885 13144
rect 10919 13141 10931 13175
rect 10873 13135 10931 13141
rect 11790 13132 11796 13184
rect 11848 13132 11854 13184
rect 14550 13132 14556 13184
rect 14608 13132 14614 13184
rect 14752 13172 14780 13271
rect 15286 13268 15292 13320
rect 15344 13268 15350 13320
rect 15473 13311 15531 13317
rect 15473 13277 15485 13311
rect 15519 13277 15531 13311
rect 15473 13271 15531 13277
rect 14826 13200 14832 13252
rect 14884 13200 14890 13252
rect 15102 13249 15108 13252
rect 15059 13243 15108 13249
rect 15059 13209 15071 13243
rect 15105 13209 15108 13243
rect 15059 13203 15108 13209
rect 15102 13200 15108 13203
rect 15160 13200 15166 13252
rect 15381 13243 15439 13249
rect 15381 13240 15393 13243
rect 15212 13212 15393 13240
rect 15212 13172 15240 13212
rect 15381 13209 15393 13212
rect 15427 13209 15439 13243
rect 15488 13240 15516 13271
rect 16298 13268 16304 13320
rect 16356 13268 16362 13320
rect 19150 13268 19156 13320
rect 19208 13308 19214 13320
rect 19613 13311 19671 13317
rect 19613 13308 19625 13311
rect 19208 13280 19625 13308
rect 19208 13268 19214 13280
rect 19613 13277 19625 13280
rect 19659 13308 19671 13311
rect 19702 13308 19708 13320
rect 19659 13280 19708 13308
rect 19659 13277 19671 13280
rect 19613 13271 19671 13277
rect 19702 13268 19708 13280
rect 19760 13268 19766 13320
rect 20441 13311 20499 13317
rect 20441 13277 20453 13311
rect 20487 13277 20499 13311
rect 20441 13271 20499 13277
rect 20533 13311 20591 13317
rect 20533 13277 20545 13311
rect 20579 13308 20591 13311
rect 20916 13308 20944 13416
rect 21266 13404 21272 13416
rect 21324 13404 21330 13456
rect 24397 13447 24455 13453
rect 24397 13444 24409 13447
rect 22066 13416 24409 13444
rect 21177 13379 21235 13385
rect 21177 13345 21189 13379
rect 21223 13376 21235 13379
rect 21223 13348 21772 13376
rect 21223 13345 21235 13348
rect 21177 13339 21235 13345
rect 20579 13280 20944 13308
rect 20579 13277 20591 13280
rect 20533 13271 20591 13277
rect 15746 13240 15752 13252
rect 15488 13212 15752 13240
rect 15381 13203 15439 13209
rect 15746 13200 15752 13212
rect 15804 13240 15810 13252
rect 15804 13212 16528 13240
rect 15804 13200 15810 13212
rect 16500 13181 16528 13212
rect 19334 13200 19340 13252
rect 19392 13240 19398 13252
rect 20162 13240 20168 13252
rect 19392 13212 20168 13240
rect 19392 13200 19398 13212
rect 20162 13200 20168 13212
rect 20220 13200 20226 13252
rect 14752 13144 15240 13172
rect 16485 13175 16543 13181
rect 16485 13141 16497 13175
rect 16531 13172 16543 13175
rect 16942 13172 16948 13184
rect 16531 13144 16948 13172
rect 16531 13141 16543 13144
rect 16485 13135 16543 13141
rect 16942 13132 16948 13144
rect 17000 13132 17006 13184
rect 19429 13175 19487 13181
rect 19429 13141 19441 13175
rect 19475 13172 19487 13175
rect 19518 13172 19524 13184
rect 19475 13144 19524 13172
rect 19475 13141 19487 13144
rect 19429 13135 19487 13141
rect 19518 13132 19524 13144
rect 19576 13132 19582 13184
rect 20456 13172 20484 13271
rect 20990 13268 20996 13320
rect 21048 13308 21054 13320
rect 21269 13311 21327 13317
rect 21269 13308 21281 13311
rect 21048 13280 21281 13308
rect 21048 13268 21054 13280
rect 21269 13277 21281 13280
rect 21315 13277 21327 13311
rect 21269 13271 21327 13277
rect 21450 13268 21456 13320
rect 21508 13268 21514 13320
rect 21744 13317 21772 13348
rect 21729 13311 21787 13317
rect 21729 13277 21741 13311
rect 21775 13308 21787 13311
rect 22066 13308 22094 13416
rect 24397 13413 24409 13416
rect 24443 13413 24455 13447
rect 25314 13444 25320 13456
rect 24397 13407 24455 13413
rect 24596 13416 25320 13444
rect 24596 13317 24624 13416
rect 25314 13404 25320 13416
rect 25372 13444 25378 13456
rect 26142 13444 26148 13456
rect 25372 13416 26148 13444
rect 25372 13404 25378 13416
rect 26142 13404 26148 13416
rect 26200 13404 26206 13456
rect 25774 13336 25780 13388
rect 25832 13376 25838 13388
rect 25869 13379 25927 13385
rect 25869 13376 25881 13379
rect 25832 13348 25881 13376
rect 25832 13336 25838 13348
rect 25869 13345 25881 13348
rect 25915 13345 25927 13379
rect 25869 13339 25927 13345
rect 25961 13379 26019 13385
rect 25961 13345 25973 13379
rect 26007 13376 26019 13379
rect 26326 13376 26332 13388
rect 26007 13348 26332 13376
rect 26007 13345 26019 13348
rect 25961 13339 26019 13345
rect 26326 13336 26332 13348
rect 26384 13336 26390 13388
rect 21775 13280 22094 13308
rect 24581 13311 24639 13317
rect 21775 13277 21787 13280
rect 21729 13271 21787 13277
rect 24581 13277 24593 13311
rect 24627 13277 24639 13311
rect 24581 13271 24639 13277
rect 24673 13311 24731 13317
rect 24673 13277 24685 13311
rect 24719 13277 24731 13311
rect 24673 13271 24731 13277
rect 26053 13311 26111 13317
rect 26053 13277 26065 13311
rect 26099 13277 26111 13311
rect 26053 13271 26111 13277
rect 20622 13200 20628 13252
rect 20680 13240 20686 13252
rect 21545 13243 21603 13249
rect 21545 13240 21557 13243
rect 20680 13212 21557 13240
rect 20680 13200 20686 13212
rect 21545 13209 21557 13212
rect 21591 13209 21603 13243
rect 23109 13243 23167 13249
rect 21545 13203 21603 13209
rect 22756 13212 23060 13240
rect 20530 13172 20536 13184
rect 20456 13144 20536 13172
rect 20530 13132 20536 13144
rect 20588 13172 20594 13184
rect 22756 13181 22784 13212
rect 22922 13181 22928 13184
rect 21913 13175 21971 13181
rect 21913 13172 21925 13175
rect 20588 13144 21925 13172
rect 20588 13132 20594 13144
rect 21913 13141 21925 13144
rect 21959 13141 21971 13175
rect 21913 13135 21971 13141
rect 22741 13175 22799 13181
rect 22741 13141 22753 13175
rect 22787 13141 22799 13175
rect 22741 13135 22799 13141
rect 22909 13175 22928 13181
rect 22909 13141 22921 13175
rect 22909 13135 22928 13141
rect 22922 13132 22928 13135
rect 22980 13132 22986 13184
rect 23032 13172 23060 13212
rect 23109 13209 23121 13243
rect 23155 13240 23167 13243
rect 23290 13240 23296 13252
rect 23155 13212 23296 13240
rect 23155 13209 23167 13212
rect 23109 13203 23167 13209
rect 23290 13200 23296 13212
rect 23348 13200 23354 13252
rect 23842 13200 23848 13252
rect 23900 13240 23906 13252
rect 24688 13240 24716 13271
rect 24762 13240 24768 13252
rect 23900 13212 24768 13240
rect 23900 13200 23906 13212
rect 24762 13200 24768 13212
rect 24820 13200 24826 13252
rect 24946 13200 24952 13252
rect 25004 13240 25010 13252
rect 25041 13243 25099 13249
rect 25041 13240 25053 13243
rect 25004 13212 25053 13240
rect 25004 13200 25010 13212
rect 25041 13209 25053 13212
rect 25087 13209 25099 13243
rect 26068 13240 26096 13271
rect 26142 13268 26148 13320
rect 26200 13268 26206 13320
rect 26694 13240 26700 13252
rect 26068 13212 26700 13240
rect 25041 13203 25099 13209
rect 26694 13200 26700 13212
rect 26752 13200 26758 13252
rect 23382 13172 23388 13184
rect 23032 13144 23388 13172
rect 23382 13132 23388 13144
rect 23440 13132 23446 13184
rect 1104 13082 27876 13104
rect 1104 13030 4874 13082
rect 4926 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 27876 13082
rect 1104 13008 27876 13030
rect 10318 12928 10324 12980
rect 10376 12968 10382 12980
rect 10376 12940 10824 12968
rect 10376 12928 10382 12940
rect 10796 12912 10824 12940
rect 14826 12928 14832 12980
rect 14884 12928 14890 12980
rect 15746 12968 15752 12980
rect 15304 12940 15752 12968
rect 10060 12872 10732 12900
rect 2682 12792 2688 12844
rect 2740 12832 2746 12844
rect 3697 12835 3755 12841
rect 3697 12832 3709 12835
rect 2740 12804 3709 12832
rect 2740 12792 2746 12804
rect 3697 12801 3709 12804
rect 3743 12801 3755 12835
rect 3697 12795 3755 12801
rect 3786 12792 3792 12844
rect 3844 12792 3850 12844
rect 3970 12792 3976 12844
rect 4028 12792 4034 12844
rect 5534 12792 5540 12844
rect 5592 12832 5598 12844
rect 7009 12835 7067 12841
rect 7009 12832 7021 12835
rect 5592 12804 7021 12832
rect 5592 12792 5598 12804
rect 7009 12801 7021 12804
rect 7055 12801 7067 12835
rect 7009 12795 7067 12801
rect 8018 12792 8024 12844
rect 8076 12832 8082 12844
rect 8113 12835 8171 12841
rect 8113 12832 8125 12835
rect 8076 12804 8125 12832
rect 8076 12792 8082 12804
rect 8113 12801 8125 12804
rect 8159 12801 8171 12835
rect 8113 12795 8171 12801
rect 8386 12792 8392 12844
rect 8444 12832 8450 12844
rect 10060 12841 10088 12872
rect 10704 12844 10732 12872
rect 10778 12860 10784 12912
rect 10836 12900 10842 12912
rect 10965 12903 11023 12909
rect 10965 12900 10977 12903
rect 10836 12872 10977 12900
rect 10836 12860 10842 12872
rect 10965 12869 10977 12872
rect 11011 12869 11023 12903
rect 10965 12863 11023 12869
rect 13449 12903 13507 12909
rect 13449 12869 13461 12903
rect 13495 12900 13507 12903
rect 14093 12903 14151 12909
rect 14093 12900 14105 12903
rect 13495 12872 14105 12900
rect 13495 12869 13507 12872
rect 13449 12863 13507 12869
rect 14093 12869 14105 12872
rect 14139 12869 14151 12903
rect 14093 12863 14151 12869
rect 15197 12903 15255 12909
rect 15197 12869 15209 12903
rect 15243 12900 15255 12903
rect 15304 12900 15332 12940
rect 15746 12928 15752 12940
rect 15804 12928 15810 12980
rect 16669 12971 16727 12977
rect 16669 12968 16681 12971
rect 15856 12940 16681 12968
rect 15243 12872 15332 12900
rect 15243 12869 15255 12872
rect 15197 12863 15255 12869
rect 15378 12860 15384 12912
rect 15436 12900 15442 12912
rect 15565 12903 15623 12909
rect 15565 12900 15577 12903
rect 15436 12872 15577 12900
rect 15436 12860 15442 12872
rect 15565 12869 15577 12872
rect 15611 12869 15623 12903
rect 15565 12863 15623 12869
rect 9861 12835 9919 12841
rect 9861 12832 9873 12835
rect 8444 12804 9873 12832
rect 8444 12792 8450 12804
rect 9861 12801 9873 12804
rect 9907 12801 9919 12835
rect 9861 12795 9919 12801
rect 10045 12835 10103 12841
rect 10045 12801 10057 12835
rect 10091 12801 10103 12835
rect 10045 12795 10103 12801
rect 10134 12792 10140 12844
rect 10192 12792 10198 12844
rect 10318 12792 10324 12844
rect 10376 12792 10382 12844
rect 10410 12792 10416 12844
rect 10468 12832 10474 12844
rect 10468 12804 10640 12832
rect 10468 12792 10474 12804
rect 3881 12767 3939 12773
rect 3881 12733 3893 12767
rect 3927 12764 3939 12767
rect 4062 12764 4068 12776
rect 3927 12736 4068 12764
rect 3927 12733 3939 12736
rect 3881 12727 3939 12733
rect 4062 12724 4068 12736
rect 4120 12724 4126 12776
rect 6362 12724 6368 12776
rect 6420 12724 6426 12776
rect 6914 12724 6920 12776
rect 6972 12724 6978 12776
rect 8297 12767 8355 12773
rect 8297 12733 8309 12767
rect 8343 12764 8355 12767
rect 10152 12764 10180 12792
rect 10505 12767 10563 12773
rect 10505 12764 10517 12767
rect 8343 12736 8432 12764
rect 10152 12736 10517 12764
rect 8343 12733 8355 12736
rect 8297 12727 8355 12733
rect 8404 12708 8432 12736
rect 10505 12733 10517 12736
rect 10551 12733 10563 12767
rect 10612 12764 10640 12804
rect 10686 12792 10692 12844
rect 10744 12792 10750 12844
rect 11149 12835 11207 12841
rect 11149 12801 11161 12835
rect 11195 12801 11207 12835
rect 11149 12795 11207 12801
rect 13357 12835 13415 12841
rect 13357 12801 13369 12835
rect 13403 12801 13415 12835
rect 13357 12795 13415 12801
rect 11164 12764 11192 12795
rect 10612 12736 11192 12764
rect 10505 12727 10563 12733
rect 3786 12656 3792 12708
rect 3844 12696 3850 12708
rect 5350 12696 5356 12708
rect 3844 12668 5356 12696
rect 3844 12656 3850 12668
rect 5350 12656 5356 12668
rect 5408 12656 5414 12708
rect 8386 12656 8392 12708
rect 8444 12656 8450 12708
rect 13372 12696 13400 12795
rect 13538 12792 13544 12844
rect 13596 12792 13602 12844
rect 13725 12835 13783 12841
rect 13725 12801 13737 12835
rect 13771 12832 13783 12835
rect 14550 12832 14556 12844
rect 13771 12804 14556 12832
rect 13771 12801 13783 12804
rect 13725 12795 13783 12801
rect 14550 12792 14556 12804
rect 14608 12792 14614 12844
rect 15013 12835 15071 12841
rect 15013 12832 15025 12835
rect 14660 12804 15025 12832
rect 14660 12776 14688 12804
rect 15013 12801 15025 12804
rect 15059 12832 15071 12835
rect 15286 12832 15292 12844
rect 15059 12804 15292 12832
rect 15059 12801 15071 12804
rect 15013 12795 15071 12801
rect 15286 12792 15292 12804
rect 15344 12792 15350 12844
rect 15473 12835 15531 12841
rect 15473 12801 15485 12835
rect 15519 12801 15531 12835
rect 15473 12795 15531 12801
rect 13998 12724 14004 12776
rect 14056 12764 14062 12776
rect 14642 12764 14648 12776
rect 14056 12736 14648 12764
rect 14056 12724 14062 12736
rect 14642 12724 14648 12736
rect 14700 12724 14706 12776
rect 15488 12764 15516 12795
rect 15028 12736 15516 12764
rect 15580 12764 15608 12863
rect 15654 12860 15660 12912
rect 15712 12860 15718 12912
rect 15856 12841 15884 12940
rect 16669 12937 16681 12940
rect 16715 12937 16727 12971
rect 16669 12931 16727 12937
rect 18325 12971 18383 12977
rect 18325 12937 18337 12971
rect 18371 12968 18383 12971
rect 19150 12968 19156 12980
rect 18371 12940 19156 12968
rect 18371 12937 18383 12940
rect 18325 12931 18383 12937
rect 19150 12928 19156 12940
rect 19208 12928 19214 12980
rect 20346 12928 20352 12980
rect 20404 12968 20410 12980
rect 20441 12971 20499 12977
rect 20441 12968 20453 12971
rect 20404 12940 20453 12968
rect 20404 12928 20410 12940
rect 20441 12937 20453 12940
rect 20487 12937 20499 12971
rect 20441 12931 20499 12937
rect 20714 12928 20720 12980
rect 20772 12968 20778 12980
rect 20772 12940 24164 12968
rect 20772 12928 20778 12940
rect 16485 12903 16543 12909
rect 16485 12869 16497 12903
rect 16531 12869 16543 12903
rect 16485 12863 16543 12869
rect 18785 12903 18843 12909
rect 18785 12869 18797 12903
rect 18831 12900 18843 12903
rect 19334 12900 19340 12912
rect 18831 12872 19340 12900
rect 18831 12869 18843 12872
rect 18785 12863 18843 12869
rect 15841 12835 15899 12841
rect 15841 12801 15853 12835
rect 15887 12801 15899 12835
rect 15841 12795 15899 12801
rect 16209 12835 16267 12841
rect 16209 12801 16221 12835
rect 16255 12801 16267 12835
rect 16209 12795 16267 12801
rect 16114 12764 16120 12776
rect 15580 12736 16120 12764
rect 14090 12696 14096 12708
rect 13372 12668 14096 12696
rect 14090 12656 14096 12668
rect 14148 12696 14154 12708
rect 15028 12696 15056 12736
rect 16114 12724 16120 12736
rect 16172 12764 16178 12776
rect 16224 12764 16252 12795
rect 16298 12792 16304 12844
rect 16356 12792 16362 12844
rect 16500 12832 16528 12863
rect 16853 12835 16911 12841
rect 16853 12832 16865 12835
rect 16500 12804 16865 12832
rect 16853 12801 16865 12804
rect 16899 12801 16911 12835
rect 16853 12795 16911 12801
rect 16942 12792 16948 12844
rect 17000 12792 17006 12844
rect 17221 12835 17279 12841
rect 17221 12801 17233 12835
rect 17267 12832 17279 12835
rect 18417 12835 18475 12841
rect 18417 12832 18429 12835
rect 17267 12804 18429 12832
rect 17267 12801 17279 12804
rect 17221 12795 17279 12801
rect 18417 12801 18429 12804
rect 18463 12801 18475 12835
rect 18417 12795 18475 12801
rect 18601 12835 18659 12841
rect 18601 12801 18613 12835
rect 18647 12801 18659 12835
rect 18601 12795 18659 12801
rect 16172 12736 16252 12764
rect 16172 12724 16178 12736
rect 16390 12724 16396 12776
rect 16448 12764 16454 12776
rect 16485 12767 16543 12773
rect 16485 12764 16497 12767
rect 16448 12736 16497 12764
rect 16448 12724 16454 12736
rect 16485 12733 16497 12736
rect 16531 12733 16543 12767
rect 16485 12727 16543 12733
rect 17310 12724 17316 12776
rect 17368 12724 17374 12776
rect 17862 12724 17868 12776
rect 17920 12724 17926 12776
rect 17957 12767 18015 12773
rect 17957 12733 17969 12767
rect 18003 12764 18015 12767
rect 18616 12764 18644 12795
rect 18874 12792 18880 12844
rect 18932 12792 18938 12844
rect 19168 12841 19196 12872
rect 19334 12860 19340 12872
rect 19392 12860 19398 12912
rect 19702 12860 19708 12912
rect 19760 12900 19766 12912
rect 23842 12900 23848 12912
rect 19760 12872 23848 12900
rect 19760 12860 19766 12872
rect 23842 12860 23848 12872
rect 23900 12860 23906 12912
rect 24136 12909 24164 12940
rect 24854 12928 24860 12980
rect 24912 12968 24918 12980
rect 26145 12971 26203 12977
rect 24912 12940 26004 12968
rect 24912 12928 24918 12940
rect 23937 12903 23995 12909
rect 23937 12869 23949 12903
rect 23983 12900 23995 12903
rect 24029 12903 24087 12909
rect 24029 12900 24041 12903
rect 23983 12872 24041 12900
rect 23983 12869 23995 12872
rect 23937 12863 23995 12869
rect 24029 12869 24041 12872
rect 24075 12869 24087 12903
rect 24029 12863 24087 12869
rect 24121 12903 24179 12909
rect 24121 12869 24133 12903
rect 24167 12869 24179 12903
rect 24121 12863 24179 12869
rect 24670 12860 24676 12912
rect 24728 12900 24734 12912
rect 25976 12909 26004 12940
rect 26145 12937 26157 12971
rect 26191 12968 26203 12971
rect 26326 12968 26332 12980
rect 26191 12940 26332 12968
rect 26191 12937 26203 12940
rect 26145 12931 26203 12937
rect 26326 12928 26332 12940
rect 26384 12928 26390 12980
rect 25961 12903 26019 12909
rect 24728 12872 25084 12900
rect 24728 12860 24734 12872
rect 19153 12835 19211 12841
rect 19153 12801 19165 12835
rect 19199 12801 19211 12835
rect 19153 12795 19211 12801
rect 20254 12792 20260 12844
rect 20312 12832 20318 12844
rect 20349 12835 20407 12841
rect 20349 12832 20361 12835
rect 20312 12804 20361 12832
rect 20312 12792 20318 12804
rect 20349 12801 20361 12804
rect 20395 12801 20407 12835
rect 20349 12795 20407 12801
rect 20717 12835 20775 12841
rect 20717 12801 20729 12835
rect 20763 12832 20775 12835
rect 21818 12832 21824 12844
rect 20763 12804 21824 12832
rect 20763 12801 20775 12804
rect 20717 12795 20775 12801
rect 21818 12792 21824 12804
rect 21876 12792 21882 12844
rect 25056 12841 25084 12872
rect 25961 12869 25973 12903
rect 26007 12869 26019 12903
rect 25961 12863 26019 12869
rect 26234 12860 26240 12912
rect 26292 12900 26298 12912
rect 26602 12900 26608 12912
rect 26292 12872 26608 12900
rect 26292 12860 26298 12872
rect 26602 12860 26608 12872
rect 26660 12860 26666 12912
rect 23661 12835 23719 12841
rect 23661 12801 23673 12835
rect 23707 12801 23719 12835
rect 23661 12795 23719 12801
rect 23753 12835 23811 12841
rect 23753 12801 23765 12835
rect 23799 12832 23811 12835
rect 24397 12835 24455 12841
rect 24397 12832 24409 12835
rect 23799 12804 24409 12832
rect 23799 12801 23811 12804
rect 23753 12795 23811 12801
rect 24397 12801 24409 12804
rect 24443 12832 24455 12835
rect 25041 12835 25099 12841
rect 24443 12804 24992 12832
rect 24443 12801 24455 12804
rect 24397 12795 24455 12801
rect 19337 12767 19395 12773
rect 19337 12764 19349 12767
rect 18003 12733 18016 12764
rect 18616 12736 19349 12764
rect 17957 12727 18016 12733
rect 19337 12733 19349 12736
rect 19383 12733 19395 12767
rect 19337 12727 19395 12733
rect 14148 12668 15056 12696
rect 14148 12656 14154 12668
rect 15102 12656 15108 12708
rect 15160 12696 15166 12708
rect 17681 12699 17739 12705
rect 17681 12696 17693 12699
rect 15160 12668 17693 12696
rect 15160 12656 15166 12668
rect 17681 12665 17693 12668
rect 17727 12665 17739 12699
rect 17681 12659 17739 12665
rect 17770 12656 17776 12708
rect 17828 12696 17834 12708
rect 17988 12696 18016 12727
rect 18969 12699 19027 12705
rect 18969 12696 18981 12699
rect 17828 12668 18981 12696
rect 17828 12656 17834 12668
rect 18969 12665 18981 12668
rect 19015 12665 19027 12699
rect 19352 12696 19380 12727
rect 20530 12724 20536 12776
rect 20588 12724 20594 12776
rect 20622 12696 20628 12708
rect 19352 12668 20628 12696
rect 18969 12659 19027 12665
rect 20622 12656 20628 12668
rect 20680 12656 20686 12708
rect 3513 12631 3571 12637
rect 3513 12597 3525 12631
rect 3559 12628 3571 12631
rect 4614 12628 4620 12640
rect 3559 12600 4620 12628
rect 3559 12597 3571 12600
rect 3513 12591 3571 12597
rect 4614 12588 4620 12600
rect 4672 12588 4678 12640
rect 7926 12588 7932 12640
rect 7984 12588 7990 12640
rect 8110 12588 8116 12640
rect 8168 12588 8174 12640
rect 10870 12588 10876 12640
rect 10928 12588 10934 12640
rect 11238 12588 11244 12640
rect 11296 12588 11302 12640
rect 13170 12588 13176 12640
rect 13228 12588 13234 12640
rect 15286 12588 15292 12640
rect 15344 12588 15350 12640
rect 20438 12588 20444 12640
rect 20496 12628 20502 12640
rect 20717 12631 20775 12637
rect 20717 12628 20729 12631
rect 20496 12600 20729 12628
rect 20496 12588 20502 12600
rect 20717 12597 20729 12600
rect 20763 12597 20775 12631
rect 23676 12628 23704 12795
rect 23937 12767 23995 12773
rect 23937 12733 23949 12767
rect 23983 12733 23995 12767
rect 23937 12727 23995 12733
rect 24581 12767 24639 12773
rect 24581 12733 24593 12767
rect 24627 12764 24639 12767
rect 24854 12764 24860 12776
rect 24627 12736 24860 12764
rect 24627 12733 24639 12736
rect 24581 12727 24639 12733
rect 23952 12696 23980 12727
rect 24854 12724 24860 12736
rect 24912 12724 24918 12776
rect 24964 12773 24992 12804
rect 25041 12801 25053 12835
rect 25087 12801 25099 12835
rect 25041 12795 25099 12801
rect 25592 12835 25650 12841
rect 25592 12801 25604 12835
rect 25638 12801 25650 12835
rect 25592 12795 25650 12801
rect 24949 12767 25007 12773
rect 24949 12733 24961 12767
rect 24995 12764 25007 12767
rect 25317 12767 25375 12773
rect 25317 12764 25329 12767
rect 24995 12736 25329 12764
rect 24995 12733 25007 12736
rect 24949 12727 25007 12733
rect 25317 12733 25329 12736
rect 25363 12733 25375 12767
rect 25607 12764 25635 12795
rect 25682 12792 25688 12844
rect 25740 12832 25746 12844
rect 25777 12835 25835 12841
rect 25777 12832 25789 12835
rect 25740 12804 25789 12832
rect 25740 12792 25746 12804
rect 25777 12801 25789 12804
rect 25823 12801 25835 12835
rect 25777 12795 25835 12801
rect 26142 12792 26148 12844
rect 26200 12832 26206 12844
rect 26421 12835 26479 12841
rect 26421 12832 26433 12835
rect 26200 12804 26433 12832
rect 26200 12792 26206 12804
rect 26421 12801 26433 12804
rect 26467 12832 26479 12835
rect 26694 12832 26700 12844
rect 26467 12804 26700 12832
rect 26467 12801 26479 12804
rect 26421 12795 26479 12801
rect 26694 12792 26700 12804
rect 26752 12792 26758 12844
rect 25607 12736 25820 12764
rect 25317 12727 25375 12733
rect 25792 12708 25820 12736
rect 26050 12724 26056 12776
rect 26108 12764 26114 12776
rect 26237 12767 26295 12773
rect 26237 12764 26249 12767
rect 26108 12736 26249 12764
rect 26108 12724 26114 12736
rect 26237 12733 26249 12736
rect 26283 12733 26295 12767
rect 26237 12727 26295 12733
rect 23952 12668 24992 12696
rect 24964 12640 24992 12668
rect 25774 12656 25780 12708
rect 25832 12656 25838 12708
rect 24394 12628 24400 12640
rect 23676 12600 24400 12628
rect 20717 12591 20775 12597
rect 24394 12588 24400 12600
rect 24452 12628 24458 12640
rect 24670 12628 24676 12640
rect 24452 12600 24676 12628
rect 24452 12588 24458 12600
rect 24670 12588 24676 12600
rect 24728 12588 24734 12640
rect 24762 12588 24768 12640
rect 24820 12588 24826 12640
rect 24946 12588 24952 12640
rect 25004 12588 25010 12640
rect 1104 12538 27876 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 27876 12538
rect 1104 12464 27876 12486
rect 4246 12384 4252 12436
rect 4304 12384 4310 12436
rect 4356 12396 5856 12424
rect 3694 12316 3700 12368
rect 3752 12356 3758 12368
rect 4356 12356 4384 12396
rect 3752 12328 4384 12356
rect 3752 12316 3758 12328
rect 5350 12316 5356 12368
rect 5408 12356 5414 12368
rect 5408 12328 5764 12356
rect 5408 12316 5414 12328
rect 3053 12291 3111 12297
rect 3053 12288 3065 12291
rect 1964 12260 3065 12288
rect 1964 12229 1992 12260
rect 3053 12257 3065 12260
rect 3099 12257 3111 12291
rect 3053 12251 3111 12257
rect 4062 12248 4068 12300
rect 4120 12248 4126 12300
rect 4706 12288 4712 12300
rect 4356 12260 4712 12288
rect 1949 12223 2007 12229
rect 1949 12189 1961 12223
rect 1995 12189 2007 12223
rect 1949 12183 2007 12189
rect 2130 12180 2136 12232
rect 2188 12180 2194 12232
rect 2314 12229 2320 12232
rect 2271 12223 2320 12229
rect 2271 12189 2283 12223
rect 2317 12189 2320 12223
rect 2271 12183 2320 12189
rect 2314 12180 2320 12183
rect 2372 12180 2378 12232
rect 2409 12223 2467 12229
rect 2409 12189 2421 12223
rect 2455 12220 2467 12223
rect 2498 12220 2504 12232
rect 2455 12192 2504 12220
rect 2455 12189 2467 12192
rect 2409 12183 2467 12189
rect 2498 12180 2504 12192
rect 2556 12220 2562 12232
rect 2685 12223 2743 12229
rect 2685 12220 2697 12223
rect 2556 12192 2697 12220
rect 2556 12180 2562 12192
rect 2685 12189 2697 12192
rect 2731 12189 2743 12223
rect 2685 12183 2743 12189
rect 2041 12155 2099 12161
rect 2041 12121 2053 12155
rect 2087 12121 2099 12155
rect 2041 12115 2099 12121
rect 1670 12044 1676 12096
rect 1728 12084 1734 12096
rect 1765 12087 1823 12093
rect 1765 12084 1777 12087
rect 1728 12056 1777 12084
rect 1728 12044 1734 12056
rect 1765 12053 1777 12056
rect 1811 12053 1823 12087
rect 2056 12084 2084 12115
rect 2501 12087 2559 12093
rect 2501 12084 2513 12087
rect 2056 12056 2513 12084
rect 1765 12047 1823 12053
rect 2501 12053 2513 12056
rect 2547 12053 2559 12087
rect 2700 12084 2728 12183
rect 2866 12180 2872 12232
rect 2924 12220 2930 12232
rect 2961 12223 3019 12229
rect 2961 12220 2973 12223
rect 2924 12192 2973 12220
rect 2924 12180 2930 12192
rect 2961 12189 2973 12192
rect 3007 12189 3019 12223
rect 2961 12183 3019 12189
rect 3145 12223 3203 12229
rect 3145 12189 3157 12223
rect 3191 12189 3203 12223
rect 3145 12183 3203 12189
rect 3160 12152 3188 12183
rect 3786 12180 3792 12232
rect 3844 12180 3850 12232
rect 3973 12223 4031 12229
rect 3973 12189 3985 12223
rect 4019 12220 4031 12223
rect 4080 12220 4108 12248
rect 4019 12192 4108 12220
rect 4019 12189 4031 12192
rect 3973 12183 4031 12189
rect 2976 12124 3188 12152
rect 4065 12155 4123 12161
rect 2976 12084 3004 12124
rect 4065 12121 4077 12155
rect 4111 12152 4123 12155
rect 4154 12152 4160 12164
rect 4111 12124 4160 12152
rect 4111 12121 4123 12124
rect 4065 12115 4123 12121
rect 4154 12112 4160 12124
rect 4212 12112 4218 12164
rect 4270 12155 4328 12161
rect 4270 12121 4282 12155
rect 4316 12152 4328 12155
rect 4356 12152 4384 12260
rect 4706 12248 4712 12260
rect 4764 12248 4770 12300
rect 5736 12297 5764 12328
rect 5261 12291 5319 12297
rect 5261 12257 5273 12291
rect 5307 12257 5319 12291
rect 5261 12251 5319 12257
rect 5721 12291 5779 12297
rect 5721 12257 5733 12291
rect 5767 12257 5779 12291
rect 5721 12251 5779 12257
rect 4525 12223 4583 12229
rect 4525 12220 4537 12223
rect 4316 12124 4384 12152
rect 4448 12192 4537 12220
rect 4316 12121 4328 12124
rect 4270 12115 4328 12121
rect 2700 12056 3004 12084
rect 2501 12047 2559 12053
rect 3234 12044 3240 12096
rect 3292 12084 3298 12096
rect 4448 12093 4476 12192
rect 4525 12189 4537 12192
rect 4571 12189 4583 12223
rect 4525 12183 4583 12189
rect 4614 12180 4620 12232
rect 4672 12220 4678 12232
rect 5276 12220 5304 12251
rect 4672 12192 5304 12220
rect 4672 12180 4678 12192
rect 5350 12180 5356 12232
rect 5408 12180 5414 12232
rect 5828 12229 5856 12396
rect 6730 12384 6736 12436
rect 6788 12424 6794 12436
rect 7285 12427 7343 12433
rect 7285 12424 7297 12427
rect 6788 12396 7297 12424
rect 6788 12384 6794 12396
rect 7285 12393 7297 12396
rect 7331 12424 7343 12427
rect 7331 12396 7696 12424
rect 7331 12393 7343 12396
rect 7285 12387 7343 12393
rect 6656 12260 7052 12288
rect 6656 12229 6684 12260
rect 7024 12232 7052 12260
rect 7282 12248 7288 12300
rect 7340 12288 7346 12300
rect 7668 12297 7696 12396
rect 8018 12384 8024 12436
rect 8076 12424 8082 12436
rect 8205 12427 8263 12433
rect 8205 12424 8217 12427
rect 8076 12396 8217 12424
rect 8076 12384 8082 12396
rect 8205 12393 8217 12396
rect 8251 12393 8263 12427
rect 8205 12387 8263 12393
rect 8386 12384 8392 12436
rect 8444 12424 8450 12436
rect 8570 12424 8576 12436
rect 8444 12396 8576 12424
rect 8444 12384 8450 12396
rect 8570 12384 8576 12396
rect 8628 12384 8634 12436
rect 9401 12427 9459 12433
rect 8680 12396 9352 12424
rect 7653 12291 7711 12297
rect 7340 12260 7604 12288
rect 7340 12248 7346 12260
rect 7576 12232 7604 12260
rect 7653 12257 7665 12291
rect 7699 12257 7711 12291
rect 7653 12251 7711 12257
rect 7745 12291 7803 12297
rect 7745 12257 7757 12291
rect 7791 12288 7803 12291
rect 8036 12288 8064 12384
rect 7791 12260 8064 12288
rect 8128 12328 8616 12356
rect 7791 12257 7803 12260
rect 7745 12251 7803 12257
rect 5813 12223 5871 12229
rect 5813 12189 5825 12223
rect 5859 12189 5871 12223
rect 5813 12183 5871 12189
rect 6641 12223 6699 12229
rect 6641 12189 6653 12223
rect 6687 12189 6699 12223
rect 6641 12183 6699 12189
rect 6825 12223 6883 12229
rect 6825 12189 6837 12223
rect 6871 12189 6883 12223
rect 6825 12183 6883 12189
rect 6840 12152 6868 12183
rect 7006 12180 7012 12232
rect 7064 12180 7070 12232
rect 7101 12223 7159 12229
rect 7101 12189 7113 12223
rect 7147 12189 7159 12223
rect 7101 12183 7159 12189
rect 7116 12152 7144 12183
rect 7374 12180 7380 12232
rect 7432 12180 7438 12232
rect 7558 12180 7564 12232
rect 7616 12180 7622 12232
rect 7929 12223 7987 12229
rect 7929 12189 7941 12223
rect 7975 12220 7987 12223
rect 8128 12220 8156 12328
rect 8202 12248 8208 12300
rect 8260 12288 8266 12300
rect 8260 12260 8524 12288
rect 8260 12248 8266 12260
rect 7975 12192 8156 12220
rect 7975 12189 7987 12192
rect 7929 12183 7987 12189
rect 8386 12180 8392 12232
rect 8444 12180 8450 12232
rect 8496 12229 8524 12260
rect 8481 12223 8539 12229
rect 8481 12189 8493 12223
rect 8527 12189 8539 12223
rect 8481 12183 8539 12189
rect 8404 12152 8432 12180
rect 6840 12124 8432 12152
rect 8588 12152 8616 12328
rect 8680 12232 8708 12396
rect 9122 12356 9128 12368
rect 8772 12328 9128 12356
rect 8662 12180 8668 12232
rect 8720 12180 8726 12232
rect 8772 12229 8800 12328
rect 9122 12316 9128 12328
rect 9180 12356 9186 12368
rect 9217 12359 9275 12365
rect 9217 12356 9229 12359
rect 9180 12328 9229 12356
rect 9180 12316 9186 12328
rect 9217 12325 9229 12328
rect 9263 12325 9275 12359
rect 9324 12356 9352 12396
rect 9401 12393 9413 12427
rect 9447 12424 9459 12427
rect 9766 12424 9772 12436
rect 9447 12396 9772 12424
rect 9447 12393 9459 12396
rect 9401 12387 9459 12393
rect 9766 12384 9772 12396
rect 9824 12384 9830 12436
rect 16114 12384 16120 12436
rect 16172 12424 16178 12436
rect 16853 12427 16911 12433
rect 16853 12424 16865 12427
rect 16172 12396 16865 12424
rect 16172 12384 16178 12396
rect 16853 12393 16865 12396
rect 16899 12393 16911 12427
rect 16853 12387 16911 12393
rect 17310 12384 17316 12436
rect 17368 12424 17374 12436
rect 17589 12427 17647 12433
rect 17589 12424 17601 12427
rect 17368 12396 17601 12424
rect 17368 12384 17374 12396
rect 17589 12393 17601 12396
rect 17635 12393 17647 12427
rect 17589 12387 17647 12393
rect 19610 12384 19616 12436
rect 19668 12384 19674 12436
rect 20349 12427 20407 12433
rect 20349 12393 20361 12427
rect 20395 12424 20407 12427
rect 20622 12424 20628 12436
rect 20395 12396 20628 12424
rect 20395 12393 20407 12396
rect 20349 12387 20407 12393
rect 20622 12384 20628 12396
rect 20680 12384 20686 12436
rect 21637 12427 21695 12433
rect 21637 12393 21649 12427
rect 21683 12424 21695 12427
rect 21726 12424 21732 12436
rect 21683 12396 21732 12424
rect 21683 12393 21695 12396
rect 21637 12387 21695 12393
rect 21726 12384 21732 12396
rect 21784 12384 21790 12436
rect 25685 12427 25743 12433
rect 25685 12393 25697 12427
rect 25731 12424 25743 12427
rect 25774 12424 25780 12436
rect 25731 12396 25780 12424
rect 25731 12393 25743 12396
rect 25685 12387 25743 12393
rect 25774 12384 25780 12396
rect 25832 12384 25838 12436
rect 9953 12359 10011 12365
rect 9953 12356 9965 12359
rect 9324 12328 9965 12356
rect 9217 12319 9275 12325
rect 9953 12325 9965 12328
rect 9999 12325 10011 12359
rect 22833 12359 22891 12365
rect 22833 12356 22845 12359
rect 9953 12319 10011 12325
rect 20548 12328 22845 12356
rect 12176 12260 12664 12288
rect 12176 12232 12204 12260
rect 8757 12223 8815 12229
rect 8757 12189 8769 12223
rect 8803 12189 8815 12223
rect 8757 12183 8815 12189
rect 9490 12180 9496 12232
rect 9548 12220 9554 12232
rect 9677 12223 9735 12229
rect 9677 12220 9689 12223
rect 9548 12192 9689 12220
rect 9548 12180 9554 12192
rect 9677 12189 9689 12192
rect 9723 12189 9735 12223
rect 9677 12183 9735 12189
rect 9766 12180 9772 12232
rect 9824 12180 9830 12232
rect 9953 12223 10011 12229
rect 9953 12189 9965 12223
rect 9999 12220 10011 12223
rect 10226 12220 10232 12232
rect 9999 12192 10232 12220
rect 9999 12189 10011 12192
rect 9953 12183 10011 12189
rect 9030 12152 9036 12164
rect 8588 12124 9036 12152
rect 9030 12112 9036 12124
rect 9088 12112 9094 12164
rect 9385 12155 9443 12161
rect 9385 12121 9397 12155
rect 9431 12152 9443 12155
rect 9508 12152 9536 12180
rect 9431 12124 9536 12152
rect 9585 12155 9643 12161
rect 9431 12121 9443 12124
rect 9385 12115 9443 12121
rect 9585 12121 9597 12155
rect 9631 12152 9643 12155
rect 9968 12152 9996 12183
rect 10226 12180 10232 12192
rect 10284 12180 10290 12232
rect 10778 12180 10784 12232
rect 10836 12220 10842 12232
rect 11606 12220 11612 12232
rect 10836 12192 11612 12220
rect 10836 12180 10842 12192
rect 11606 12180 11612 12192
rect 11664 12180 11670 12232
rect 11790 12180 11796 12232
rect 11848 12220 11854 12232
rect 11977 12223 12035 12229
rect 11977 12220 11989 12223
rect 11848 12192 11989 12220
rect 11848 12180 11854 12192
rect 11977 12189 11989 12192
rect 12023 12189 12035 12223
rect 11977 12183 12035 12189
rect 9631 12124 9996 12152
rect 11992 12152 12020 12183
rect 12158 12180 12164 12232
rect 12216 12180 12222 12232
rect 12636 12229 12664 12260
rect 15470 12248 15476 12300
rect 15528 12248 15534 12300
rect 20548 12297 20576 12328
rect 22833 12325 22845 12328
rect 22879 12325 22891 12359
rect 27154 12356 27160 12368
rect 22833 12319 22891 12325
rect 25056 12328 27160 12356
rect 20073 12291 20131 12297
rect 20073 12257 20085 12291
rect 20119 12288 20131 12291
rect 20533 12291 20591 12297
rect 20533 12288 20545 12291
rect 20119 12260 20545 12288
rect 20119 12257 20131 12260
rect 20073 12251 20131 12257
rect 20533 12257 20545 12260
rect 20579 12257 20591 12291
rect 20533 12251 20591 12257
rect 22005 12291 22063 12297
rect 22005 12257 22017 12291
rect 22051 12288 22063 12291
rect 22465 12291 22523 12297
rect 22465 12288 22477 12291
rect 22051 12260 22477 12288
rect 22051 12257 22063 12260
rect 22005 12251 22063 12257
rect 22465 12257 22477 12260
rect 22511 12257 22523 12291
rect 22465 12251 22523 12257
rect 22741 12291 22799 12297
rect 22741 12257 22753 12291
rect 22787 12288 22799 12291
rect 22787 12260 23244 12288
rect 22787 12257 22799 12260
rect 22741 12251 22799 12257
rect 12437 12223 12495 12229
rect 12437 12189 12449 12223
rect 12483 12189 12495 12223
rect 12437 12183 12495 12189
rect 12621 12223 12679 12229
rect 12621 12189 12633 12223
rect 12667 12189 12679 12223
rect 12621 12183 12679 12189
rect 12452 12152 12480 12183
rect 15286 12180 15292 12232
rect 15344 12220 15350 12232
rect 15729 12223 15787 12229
rect 15729 12220 15741 12223
rect 15344 12192 15741 12220
rect 15344 12180 15350 12192
rect 15729 12189 15741 12192
rect 15775 12189 15787 12223
rect 15729 12183 15787 12189
rect 17218 12180 17224 12232
rect 17276 12220 17282 12232
rect 17589 12223 17647 12229
rect 17589 12220 17601 12223
rect 17276 12192 17601 12220
rect 17276 12180 17282 12192
rect 17589 12189 17601 12192
rect 17635 12189 17647 12223
rect 17589 12183 17647 12189
rect 17770 12180 17776 12232
rect 17828 12180 17834 12232
rect 17865 12223 17923 12229
rect 17865 12189 17877 12223
rect 17911 12220 17923 12223
rect 18230 12220 18236 12232
rect 17911 12192 18236 12220
rect 17911 12189 17923 12192
rect 17865 12183 17923 12189
rect 18230 12180 18236 12192
rect 18288 12180 18294 12232
rect 19981 12223 20039 12229
rect 19981 12189 19993 12223
rect 20027 12220 20039 12223
rect 20625 12223 20683 12229
rect 20625 12220 20637 12223
rect 20027 12192 20637 12220
rect 20027 12189 20039 12192
rect 19981 12183 20039 12189
rect 20625 12189 20637 12192
rect 20671 12189 20683 12223
rect 20625 12183 20683 12189
rect 21913 12223 21971 12229
rect 21913 12189 21925 12223
rect 21959 12220 21971 12223
rect 22373 12223 22431 12229
rect 21959 12192 22094 12220
rect 21959 12189 21971 12192
rect 21913 12183 21971 12189
rect 11992 12124 12480 12152
rect 9631 12121 9643 12124
rect 9585 12115 9643 12121
rect 3881 12087 3939 12093
rect 3881 12084 3893 12087
rect 3292 12056 3893 12084
rect 3292 12044 3298 12056
rect 3881 12053 3893 12056
rect 3927 12053 3939 12087
rect 3881 12047 3939 12053
rect 4433 12087 4491 12093
rect 4433 12053 4445 12087
rect 4479 12053 4491 12087
rect 4433 12047 4491 12053
rect 4798 12044 4804 12096
rect 4856 12044 4862 12096
rect 6733 12087 6791 12093
rect 6733 12053 6745 12087
rect 6779 12084 6791 12087
rect 6822 12084 6828 12096
rect 6779 12056 6828 12084
rect 6779 12053 6791 12056
rect 6733 12047 6791 12053
rect 6822 12044 6828 12056
rect 6880 12044 6886 12096
rect 7006 12044 7012 12096
rect 7064 12084 7070 12096
rect 8018 12084 8024 12096
rect 7064 12056 8024 12084
rect 7064 12044 7070 12056
rect 8018 12044 8024 12056
rect 8076 12044 8082 12096
rect 8110 12044 8116 12096
rect 8168 12044 8174 12096
rect 11330 12044 11336 12096
rect 11388 12084 11394 12096
rect 11701 12087 11759 12093
rect 11701 12084 11713 12087
rect 11388 12056 11713 12084
rect 11388 12044 11394 12056
rect 11701 12053 11713 12056
rect 11747 12053 11759 12087
rect 11701 12047 11759 12053
rect 12345 12087 12403 12093
rect 12345 12053 12357 12087
rect 12391 12084 12403 12087
rect 12434 12084 12440 12096
rect 12391 12056 12440 12084
rect 12391 12053 12403 12056
rect 12345 12047 12403 12053
rect 12434 12044 12440 12056
rect 12492 12044 12498 12096
rect 12529 12087 12587 12093
rect 12529 12053 12541 12087
rect 12575 12084 12587 12087
rect 12618 12084 12624 12096
rect 12575 12056 12624 12084
rect 12575 12053 12587 12056
rect 12529 12047 12587 12053
rect 12618 12044 12624 12056
rect 12676 12044 12682 12096
rect 20640 12084 20668 12183
rect 22066 12152 22094 12192
rect 22373 12189 22385 12223
rect 22419 12189 22431 12223
rect 22480 12220 22508 12251
rect 23216 12232 23244 12260
rect 24486 12248 24492 12300
rect 24544 12288 24550 12300
rect 25056 12297 25084 12328
rect 27154 12316 27160 12328
rect 27212 12316 27218 12368
rect 25041 12291 25099 12297
rect 25041 12288 25053 12291
rect 24544 12260 25053 12288
rect 24544 12248 24550 12260
rect 25041 12257 25053 12260
rect 25087 12257 25099 12291
rect 25041 12251 25099 12257
rect 25225 12291 25283 12297
rect 25225 12257 25237 12291
rect 25271 12288 25283 12291
rect 25682 12288 25688 12300
rect 25271 12260 25688 12288
rect 25271 12257 25283 12260
rect 25225 12251 25283 12257
rect 25682 12248 25688 12260
rect 25740 12248 25746 12300
rect 23014 12220 23020 12232
rect 22480 12192 23020 12220
rect 22373 12183 22431 12189
rect 22388 12152 22416 12183
rect 23014 12180 23020 12192
rect 23072 12180 23078 12232
rect 23198 12180 23204 12232
rect 23256 12180 23262 12232
rect 23382 12180 23388 12232
rect 23440 12180 23446 12232
rect 25498 12220 25504 12232
rect 25240 12192 25504 12220
rect 25240 12164 25268 12192
rect 25498 12180 25504 12192
rect 25556 12180 25562 12232
rect 25869 12223 25927 12229
rect 25869 12189 25881 12223
rect 25915 12220 25927 12223
rect 25958 12220 25964 12232
rect 25915 12192 25964 12220
rect 25915 12189 25927 12192
rect 25869 12183 25927 12189
rect 25958 12180 25964 12192
rect 26016 12180 26022 12232
rect 23109 12155 23167 12161
rect 23109 12152 23121 12155
rect 22066 12124 23121 12152
rect 23109 12121 23121 12124
rect 23155 12152 23167 12155
rect 24026 12152 24032 12164
rect 23155 12124 24032 12152
rect 23155 12121 23167 12124
rect 23109 12115 23167 12121
rect 24026 12112 24032 12124
rect 24084 12112 24090 12164
rect 25222 12112 25228 12164
rect 25280 12112 25286 12164
rect 22922 12084 22928 12096
rect 20640 12056 22928 12084
rect 22922 12044 22928 12056
rect 22980 12084 22986 12096
rect 23934 12084 23940 12096
rect 22980 12056 23940 12084
rect 22980 12044 22986 12056
rect 23934 12044 23940 12056
rect 23992 12044 23998 12096
rect 25406 12044 25412 12096
rect 25464 12084 25470 12096
rect 25682 12084 25688 12096
rect 25464 12056 25688 12084
rect 25464 12044 25470 12056
rect 25682 12044 25688 12056
rect 25740 12044 25746 12096
rect 1104 11994 27876 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 27876 11994
rect 1104 11920 27876 11942
rect 2498 11840 2504 11892
rect 2556 11880 2562 11892
rect 2777 11883 2835 11889
rect 2777 11880 2789 11883
rect 2556 11852 2789 11880
rect 2556 11840 2562 11852
rect 2777 11849 2789 11852
rect 2823 11849 2835 11883
rect 2777 11843 2835 11849
rect 10689 11883 10747 11889
rect 10689 11849 10701 11883
rect 10735 11880 10747 11883
rect 12158 11880 12164 11892
rect 10735 11852 12164 11880
rect 10735 11849 10747 11852
rect 10689 11843 10747 11849
rect 2406 11812 2412 11824
rect 1412 11784 2412 11812
rect 1412 11753 1440 11784
rect 2406 11772 2412 11784
rect 2464 11772 2470 11824
rect 1670 11753 1676 11756
rect 1397 11747 1455 11753
rect 1397 11713 1409 11747
rect 1443 11713 1455 11747
rect 1664 11744 1676 11753
rect 1631 11716 1676 11744
rect 1397 11707 1455 11713
rect 1664 11707 1676 11716
rect 1670 11704 1676 11707
rect 1728 11704 1734 11756
rect 2792 11744 2820 11843
rect 12158 11840 12164 11852
rect 12216 11840 12222 11892
rect 14642 11840 14648 11892
rect 14700 11840 14706 11892
rect 18969 11883 19027 11889
rect 18969 11849 18981 11883
rect 19015 11880 19027 11883
rect 19978 11880 19984 11892
rect 19015 11852 19984 11880
rect 19015 11849 19027 11852
rect 18969 11843 19027 11849
rect 19978 11840 19984 11852
rect 20036 11840 20042 11892
rect 23198 11840 23204 11892
rect 23256 11880 23262 11892
rect 24137 11883 24195 11889
rect 24137 11880 24149 11883
rect 23256 11852 24149 11880
rect 23256 11840 23262 11852
rect 24137 11849 24149 11852
rect 24183 11849 24195 11883
rect 24137 11843 24195 11849
rect 24305 11883 24363 11889
rect 24305 11849 24317 11883
rect 24351 11880 24363 11883
rect 24486 11880 24492 11892
rect 24351 11852 24492 11880
rect 24351 11849 24363 11852
rect 24305 11843 24363 11849
rect 24486 11840 24492 11852
rect 24544 11840 24550 11892
rect 24765 11883 24823 11889
rect 24765 11849 24777 11883
rect 24811 11880 24823 11883
rect 24854 11880 24860 11892
rect 24811 11852 24860 11880
rect 24811 11849 24823 11852
rect 24765 11843 24823 11849
rect 24854 11840 24860 11852
rect 24912 11880 24918 11892
rect 24912 11852 25452 11880
rect 24912 11840 24918 11852
rect 25424 11824 25452 11852
rect 3789 11815 3847 11821
rect 3789 11781 3801 11815
rect 3835 11812 3847 11815
rect 5350 11812 5356 11824
rect 3835 11784 5356 11812
rect 3835 11781 3847 11784
rect 3789 11775 3847 11781
rect 3145 11747 3203 11753
rect 3145 11744 3157 11747
rect 2792 11716 3157 11744
rect 3145 11713 3157 11716
rect 3191 11713 3203 11747
rect 3697 11747 3755 11753
rect 3697 11744 3709 11747
rect 3145 11707 3203 11713
rect 3528 11716 3709 11744
rect 3234 11636 3240 11688
rect 3292 11636 3298 11688
rect 3528 11620 3556 11716
rect 3697 11713 3709 11716
rect 3743 11713 3755 11747
rect 3697 11707 3755 11713
rect 3878 11704 3884 11756
rect 3936 11704 3942 11756
rect 4154 11704 4160 11756
rect 4212 11744 4218 11756
rect 5077 11747 5135 11753
rect 5077 11744 5089 11747
rect 4212 11716 5089 11744
rect 4212 11704 4218 11716
rect 5077 11713 5089 11716
rect 5123 11744 5135 11747
rect 5166 11744 5172 11756
rect 5123 11716 5172 11744
rect 5123 11713 5135 11716
rect 5077 11707 5135 11713
rect 5166 11704 5172 11716
rect 5224 11704 5230 11756
rect 5276 11753 5304 11784
rect 5350 11772 5356 11784
rect 5408 11772 5414 11824
rect 8110 11812 8116 11824
rect 5552 11784 8116 11812
rect 5552 11756 5580 11784
rect 8110 11772 8116 11784
rect 8168 11772 8174 11824
rect 8220 11784 10364 11812
rect 5261 11747 5319 11753
rect 5261 11713 5273 11747
rect 5307 11713 5319 11747
rect 5261 11707 5319 11713
rect 5534 11704 5540 11756
rect 5592 11704 5598 11756
rect 5718 11704 5724 11756
rect 5776 11744 5782 11756
rect 6549 11747 6607 11753
rect 5776 11716 6500 11744
rect 5776 11704 5782 11716
rect 4709 11679 4767 11685
rect 4709 11645 4721 11679
rect 4755 11676 4767 11679
rect 4798 11676 4804 11688
rect 4755 11648 4804 11676
rect 4755 11645 4767 11648
rect 4709 11639 4767 11645
rect 4798 11636 4804 11648
rect 4856 11636 4862 11688
rect 3510 11568 3516 11620
rect 3568 11568 3574 11620
rect 6089 11543 6147 11549
rect 6089 11509 6101 11543
rect 6135 11540 6147 11543
rect 6178 11540 6184 11552
rect 6135 11512 6184 11540
rect 6135 11509 6147 11512
rect 6089 11503 6147 11509
rect 6178 11500 6184 11512
rect 6236 11500 6242 11552
rect 6472 11540 6500 11716
rect 6549 11713 6561 11747
rect 6595 11744 6607 11747
rect 6638 11744 6644 11756
rect 6595 11716 6644 11744
rect 6595 11713 6607 11716
rect 6549 11707 6607 11713
rect 6638 11704 6644 11716
rect 6696 11704 6702 11756
rect 6914 11704 6920 11756
rect 6972 11704 6978 11756
rect 7193 11747 7251 11753
rect 7193 11713 7205 11747
rect 7239 11713 7251 11747
rect 7193 11707 7251 11713
rect 7837 11747 7895 11753
rect 7837 11713 7849 11747
rect 7883 11744 7895 11747
rect 8220 11744 8248 11784
rect 10336 11756 10364 11784
rect 12176 11784 12664 11812
rect 7883 11716 8248 11744
rect 7883 11713 7895 11716
rect 7837 11707 7895 11713
rect 6822 11636 6828 11688
rect 6880 11676 6886 11688
rect 7101 11679 7159 11685
rect 7101 11676 7113 11679
rect 6880 11648 7113 11676
rect 6880 11636 6886 11648
rect 7101 11645 7113 11648
rect 7147 11645 7159 11679
rect 7101 11639 7159 11645
rect 6546 11568 6552 11620
rect 6604 11608 6610 11620
rect 7208 11608 7236 11707
rect 8662 11704 8668 11756
rect 8720 11744 8726 11756
rect 8941 11747 8999 11753
rect 8941 11744 8953 11747
rect 8720 11716 8953 11744
rect 8720 11704 8726 11716
rect 8941 11713 8953 11716
rect 8987 11713 8999 11747
rect 8941 11707 8999 11713
rect 9122 11704 9128 11756
rect 9180 11704 9186 11756
rect 9398 11704 9404 11756
rect 9456 11744 9462 11756
rect 10229 11747 10287 11753
rect 10229 11744 10241 11747
rect 9456 11716 10241 11744
rect 9456 11704 9462 11716
rect 10229 11713 10241 11716
rect 10275 11713 10287 11747
rect 10229 11707 10287 11713
rect 7466 11636 7472 11688
rect 7524 11676 7530 11688
rect 7561 11679 7619 11685
rect 7561 11676 7573 11679
rect 7524 11648 7573 11676
rect 7524 11636 7530 11648
rect 7561 11645 7573 11648
rect 7607 11645 7619 11679
rect 10244 11676 10272 11707
rect 10318 11704 10324 11756
rect 10376 11704 10382 11756
rect 10505 11747 10563 11753
rect 10505 11713 10517 11747
rect 10551 11744 10563 11747
rect 10778 11744 10784 11756
rect 10551 11716 10784 11744
rect 10551 11713 10563 11716
rect 10505 11707 10563 11713
rect 10778 11704 10784 11716
rect 10836 11704 10842 11756
rect 11609 11747 11667 11753
rect 11609 11713 11621 11747
rect 11655 11744 11667 11747
rect 11698 11744 11704 11756
rect 11655 11716 11704 11744
rect 11655 11713 11667 11716
rect 11609 11707 11667 11713
rect 11698 11704 11704 11716
rect 11756 11704 11762 11756
rect 11790 11704 11796 11756
rect 11848 11704 11854 11756
rect 12176 11753 12204 11784
rect 12636 11756 12664 11784
rect 13170 11772 13176 11824
rect 13228 11812 13234 11824
rect 13510 11815 13568 11821
rect 13510 11812 13522 11815
rect 13228 11784 13522 11812
rect 13228 11772 13234 11784
rect 13510 11781 13522 11784
rect 13556 11781 13568 11815
rect 13510 11775 13568 11781
rect 18046 11772 18052 11824
rect 18104 11812 18110 11824
rect 18785 11815 18843 11821
rect 18785 11812 18797 11815
rect 18104 11784 18797 11812
rect 18104 11772 18110 11784
rect 18785 11781 18797 11784
rect 18831 11812 18843 11815
rect 19242 11812 19248 11824
rect 18831 11784 19248 11812
rect 18831 11781 18843 11784
rect 18785 11775 18843 11781
rect 19242 11772 19248 11784
rect 19300 11772 19306 11824
rect 23014 11772 23020 11824
rect 23072 11812 23078 11824
rect 23753 11815 23811 11821
rect 23753 11812 23765 11815
rect 23072 11784 23765 11812
rect 23072 11772 23078 11784
rect 23753 11781 23765 11784
rect 23799 11781 23811 11815
rect 23753 11775 23811 11781
rect 23934 11772 23940 11824
rect 23992 11772 23998 11824
rect 25406 11772 25412 11824
rect 25464 11772 25470 11824
rect 12161 11747 12219 11753
rect 12161 11713 12173 11747
rect 12207 11713 12219 11747
rect 12434 11744 12440 11756
rect 12161 11707 12219 11713
rect 12268 11716 12440 11744
rect 10962 11676 10968 11688
rect 10244 11648 10968 11676
rect 7561 11639 7619 11645
rect 10962 11636 10968 11648
rect 11020 11636 11026 11688
rect 11514 11636 11520 11688
rect 11572 11676 11578 11688
rect 11885 11679 11943 11685
rect 11885 11676 11897 11679
rect 11572 11648 11897 11676
rect 11572 11636 11578 11648
rect 11885 11645 11897 11648
rect 11931 11645 11943 11679
rect 11885 11639 11943 11645
rect 11977 11679 12035 11685
rect 11977 11645 11989 11679
rect 12023 11676 12035 11679
rect 12268 11676 12296 11716
rect 12434 11704 12440 11716
rect 12492 11704 12498 11756
rect 12618 11704 12624 11756
rect 12676 11704 12682 11756
rect 13265 11747 13323 11753
rect 13265 11713 13277 11747
rect 13311 11744 13323 11747
rect 13354 11744 13360 11756
rect 13311 11716 13360 11744
rect 13311 11713 13323 11716
rect 13265 11707 13323 11713
rect 13354 11704 13360 11716
rect 13412 11704 13418 11756
rect 18598 11704 18604 11756
rect 18656 11704 18662 11756
rect 20530 11704 20536 11756
rect 20588 11744 20594 11756
rect 20809 11747 20867 11753
rect 20809 11744 20821 11747
rect 20588 11716 20821 11744
rect 20588 11704 20594 11716
rect 20809 11713 20821 11716
rect 20855 11713 20867 11747
rect 20809 11707 20867 11713
rect 23474 11704 23480 11756
rect 23532 11704 23538 11756
rect 24394 11704 24400 11756
rect 24452 11704 24458 11756
rect 24581 11747 24639 11753
rect 24581 11713 24593 11747
rect 24627 11744 24639 11747
rect 24946 11744 24952 11756
rect 24627 11716 24952 11744
rect 24627 11713 24639 11716
rect 24581 11707 24639 11713
rect 24946 11704 24952 11716
rect 25004 11704 25010 11756
rect 25498 11704 25504 11756
rect 25556 11744 25562 11756
rect 26145 11747 26203 11753
rect 26145 11744 26157 11747
rect 25556 11716 26157 11744
rect 25556 11704 25562 11716
rect 26145 11713 26157 11716
rect 26191 11713 26203 11747
rect 26145 11707 26203 11713
rect 26237 11747 26295 11753
rect 26237 11713 26249 11747
rect 26283 11744 26295 11747
rect 26973 11747 27031 11753
rect 26973 11744 26985 11747
rect 26283 11716 26985 11744
rect 26283 11713 26295 11716
rect 26237 11707 26295 11713
rect 26973 11713 26985 11716
rect 27019 11713 27031 11747
rect 26973 11707 27031 11713
rect 27154 11704 27160 11756
rect 27212 11704 27218 11756
rect 27246 11704 27252 11756
rect 27304 11704 27310 11756
rect 12023 11648 12296 11676
rect 12023 11645 12035 11648
rect 11977 11639 12035 11645
rect 6604 11580 7236 11608
rect 11900 11608 11928 11639
rect 20898 11636 20904 11688
rect 20956 11636 20962 11688
rect 21177 11679 21235 11685
rect 21177 11645 21189 11679
rect 21223 11676 21235 11679
rect 22738 11676 22744 11688
rect 21223 11648 22744 11676
rect 21223 11645 21235 11648
rect 21177 11639 21235 11645
rect 22738 11636 22744 11648
rect 22796 11636 22802 11688
rect 23293 11679 23351 11685
rect 23293 11645 23305 11679
rect 23339 11676 23351 11679
rect 23566 11676 23572 11688
rect 23339 11648 23572 11676
rect 23339 11645 23351 11648
rect 23293 11639 23351 11645
rect 23566 11636 23572 11648
rect 23624 11636 23630 11688
rect 23842 11636 23848 11688
rect 23900 11636 23906 11688
rect 26050 11636 26056 11688
rect 26108 11636 26114 11688
rect 26329 11679 26387 11685
rect 26329 11645 26341 11679
rect 26375 11645 26387 11679
rect 26329 11639 26387 11645
rect 12526 11608 12532 11620
rect 11900 11580 12532 11608
rect 6604 11568 6610 11580
rect 12526 11568 12532 11580
rect 12584 11568 12590 11620
rect 25682 11568 25688 11620
rect 25740 11568 25746 11620
rect 25869 11611 25927 11617
rect 25869 11577 25881 11611
rect 25915 11608 25927 11611
rect 26344 11608 26372 11639
rect 25915 11580 26372 11608
rect 25915 11577 25927 11580
rect 25869 11571 25927 11577
rect 7926 11540 7932 11552
rect 6472 11512 7932 11540
rect 7926 11500 7932 11512
rect 7984 11500 7990 11552
rect 8202 11500 8208 11552
rect 8260 11540 8266 11552
rect 9125 11543 9183 11549
rect 9125 11540 9137 11543
rect 8260 11512 9137 11540
rect 8260 11500 8266 11512
rect 9125 11509 9137 11512
rect 9171 11509 9183 11543
rect 9125 11503 9183 11509
rect 11606 11500 11612 11552
rect 11664 11540 11670 11552
rect 12345 11543 12403 11549
rect 12345 11540 12357 11543
rect 11664 11512 12357 11540
rect 11664 11500 11670 11512
rect 12345 11509 12357 11512
rect 12391 11509 12403 11543
rect 12345 11503 12403 11509
rect 12437 11543 12495 11549
rect 12437 11509 12449 11543
rect 12483 11540 12495 11543
rect 12618 11540 12624 11552
rect 12483 11512 12624 11540
rect 12483 11509 12495 11512
rect 12437 11503 12495 11509
rect 12618 11500 12624 11512
rect 12676 11500 12682 11552
rect 23382 11500 23388 11552
rect 23440 11540 23446 11552
rect 24121 11543 24179 11549
rect 24121 11540 24133 11543
rect 23440 11512 24133 11540
rect 23440 11500 23446 11512
rect 24121 11509 24133 11512
rect 24167 11509 24179 11543
rect 24121 11503 24179 11509
rect 26510 11500 26516 11552
rect 26568 11500 26574 11552
rect 1104 11450 27876 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 27876 11450
rect 1104 11376 27876 11398
rect 4798 11296 4804 11348
rect 4856 11296 4862 11348
rect 8294 11296 8300 11348
rect 8352 11296 8358 11348
rect 8386 11296 8392 11348
rect 8444 11336 8450 11348
rect 8570 11336 8576 11348
rect 8444 11308 8576 11336
rect 8444 11296 8450 11308
rect 8570 11296 8576 11308
rect 8628 11336 8634 11348
rect 9125 11339 9183 11345
rect 9125 11336 9137 11339
rect 8628 11308 9137 11336
rect 8628 11296 8634 11308
rect 9125 11305 9137 11308
rect 9171 11336 9183 11339
rect 10873 11339 10931 11345
rect 9171 11308 10272 11336
rect 9171 11305 9183 11308
rect 9125 11299 9183 11305
rect 8202 11268 8208 11280
rect 7760 11240 8208 11268
rect 7377 11203 7435 11209
rect 7377 11169 7389 11203
rect 7423 11200 7435 11203
rect 7558 11200 7564 11212
rect 7423 11172 7564 11200
rect 7423 11169 7435 11172
rect 7377 11163 7435 11169
rect 7558 11160 7564 11172
rect 7616 11160 7622 11212
rect 7760 11209 7788 11240
rect 8202 11228 8208 11240
rect 8260 11228 8266 11280
rect 7745 11203 7803 11209
rect 7745 11169 7757 11203
rect 7791 11169 7803 11203
rect 7745 11163 7803 11169
rect 8113 11203 8171 11209
rect 8113 11169 8125 11203
rect 8159 11200 8171 11203
rect 8312 11200 8340 11296
rect 8159 11172 8248 11200
rect 8312 11172 8984 11200
rect 8159 11169 8171 11172
rect 8113 11163 8171 11169
rect 4338 11092 4344 11144
rect 4396 11132 4402 11144
rect 4614 11132 4620 11144
rect 4396 11104 4620 11132
rect 4396 11092 4402 11104
rect 4614 11092 4620 11104
rect 4672 11132 4678 11144
rect 4709 11135 4767 11141
rect 4709 11132 4721 11135
rect 4672 11104 4721 11132
rect 4672 11092 4678 11104
rect 4709 11101 4721 11104
rect 4755 11101 4767 11135
rect 4709 11095 4767 11101
rect 4798 11092 4804 11144
rect 4856 11132 4862 11144
rect 4893 11135 4951 11141
rect 4893 11132 4905 11135
rect 4856 11104 4905 11132
rect 4856 11092 4862 11104
rect 4893 11101 4905 11104
rect 4939 11101 4951 11135
rect 4893 11095 4951 11101
rect 5077 11135 5135 11141
rect 5077 11101 5089 11135
rect 5123 11132 5135 11135
rect 5166 11132 5172 11144
rect 5123 11104 5172 11132
rect 5123 11101 5135 11104
rect 5077 11095 5135 11101
rect 5166 11092 5172 11104
rect 5224 11092 5230 11144
rect 5534 11092 5540 11144
rect 5592 11092 5598 11144
rect 5718 11092 5724 11144
rect 5776 11092 5782 11144
rect 7837 11135 7895 11141
rect 7837 11101 7849 11135
rect 7883 11132 7895 11135
rect 7883 11104 8156 11132
rect 7883 11101 7895 11104
rect 7837 11095 7895 11101
rect 5261 11067 5319 11073
rect 5261 11033 5273 11067
rect 5307 11064 5319 11067
rect 5629 11067 5687 11073
rect 5629 11064 5641 11067
rect 5307 11036 5641 11064
rect 5307 11033 5319 11036
rect 5261 11027 5319 11033
rect 5629 11033 5641 11036
rect 5675 11033 5687 11067
rect 5629 11027 5687 11033
rect 6546 11024 6552 11076
rect 6604 11064 6610 11076
rect 8021 11067 8079 11073
rect 8021 11064 8033 11067
rect 6604 11036 8033 11064
rect 6604 11024 6610 11036
rect 8021 11033 8033 11036
rect 8067 11033 8079 11067
rect 8021 11027 8079 11033
rect 4706 10956 4712 11008
rect 4764 10996 4770 11008
rect 4890 10996 4896 11008
rect 4764 10968 4896 10996
rect 4764 10956 4770 10968
rect 4890 10956 4896 10968
rect 4948 10956 4954 11008
rect 5350 10956 5356 11008
rect 5408 10996 5414 11008
rect 8128 11005 8156 11104
rect 8220 11064 8248 11172
rect 8386 11092 8392 11144
rect 8444 11092 8450 11144
rect 8956 11141 8984 11172
rect 9030 11160 9036 11212
rect 9088 11160 9094 11212
rect 8941 11135 8999 11141
rect 8941 11101 8953 11135
rect 8987 11101 8999 11135
rect 8941 11095 8999 11101
rect 9398 11092 9404 11144
rect 9456 11132 9462 11144
rect 10244 11141 10272 11308
rect 10873 11305 10885 11339
rect 10919 11336 10931 11339
rect 11698 11336 11704 11348
rect 10919 11308 11704 11336
rect 10919 11305 10931 11308
rect 10873 11299 10931 11305
rect 11698 11296 11704 11308
rect 11756 11296 11762 11348
rect 19242 11296 19248 11348
rect 19300 11296 19306 11348
rect 22097 11339 22155 11345
rect 22097 11305 22109 11339
rect 22143 11336 22155 11339
rect 23106 11336 23112 11348
rect 22143 11308 23112 11336
rect 22143 11305 22155 11308
rect 22097 11299 22155 11305
rect 23106 11296 23112 11308
rect 23164 11296 23170 11348
rect 24302 11296 24308 11348
rect 24360 11336 24366 11348
rect 24581 11339 24639 11345
rect 24581 11336 24593 11339
rect 24360 11308 24593 11336
rect 24360 11296 24366 11308
rect 24581 11305 24593 11308
rect 24627 11305 24639 11339
rect 24581 11299 24639 11305
rect 26050 11296 26056 11348
rect 26108 11336 26114 11348
rect 26145 11339 26203 11345
rect 26145 11336 26157 11339
rect 26108 11308 26157 11336
rect 26108 11296 26114 11308
rect 26145 11305 26157 11308
rect 26191 11305 26203 11339
rect 26145 11299 26203 11305
rect 11333 11271 11391 11277
rect 11333 11268 11345 11271
rect 10704 11240 11345 11268
rect 10704 11209 10732 11240
rect 11333 11237 11345 11240
rect 11379 11237 11391 11271
rect 11333 11231 11391 11237
rect 14829 11271 14887 11277
rect 14829 11237 14841 11271
rect 14875 11268 14887 11271
rect 15470 11268 15476 11280
rect 14875 11240 15476 11268
rect 14875 11237 14887 11240
rect 14829 11231 14887 11237
rect 15470 11228 15476 11240
rect 15528 11228 15534 11280
rect 27154 11268 27160 11280
rect 26068 11240 27160 11268
rect 10689 11203 10747 11209
rect 10689 11169 10701 11203
rect 10735 11169 10747 11203
rect 10689 11163 10747 11169
rect 12618 11160 12624 11212
rect 12676 11200 12682 11212
rect 12676 11172 12848 11200
rect 12676 11160 12682 11172
rect 9953 11135 10011 11141
rect 9953 11132 9965 11135
rect 9456 11104 9965 11132
rect 9456 11092 9462 11104
rect 9953 11101 9965 11104
rect 9999 11101 10011 11135
rect 9953 11095 10011 11101
rect 10045 11135 10103 11141
rect 10045 11101 10057 11135
rect 10091 11132 10103 11135
rect 10229 11135 10287 11141
rect 10091 11104 10180 11132
rect 10091 11101 10103 11104
rect 10045 11095 10103 11101
rect 9030 11064 9036 11076
rect 8220 11036 9036 11064
rect 9030 11024 9036 11036
rect 9088 11024 9094 11076
rect 9766 11024 9772 11076
rect 9824 11024 9830 11076
rect 5445 10999 5503 11005
rect 5445 10996 5457 10999
rect 5408 10968 5457 10996
rect 5408 10956 5414 10968
rect 5445 10965 5457 10968
rect 5491 10965 5503 10999
rect 5445 10959 5503 10965
rect 8113 10999 8171 11005
rect 8113 10965 8125 10999
rect 8159 10996 8171 10999
rect 8294 10996 8300 11008
rect 8159 10968 8300 10996
rect 8159 10965 8171 10968
rect 8113 10959 8171 10965
rect 8294 10956 8300 10968
rect 8352 10956 8358 11008
rect 9122 10956 9128 11008
rect 9180 10996 9186 11008
rect 9309 10999 9367 11005
rect 9309 10996 9321 10999
rect 9180 10968 9321 10996
rect 9180 10956 9186 10968
rect 9309 10965 9321 10968
rect 9355 10965 9367 10999
rect 10152 10996 10180 11104
rect 10229 11101 10241 11135
rect 10275 11101 10287 11135
rect 10229 11095 10287 11101
rect 10321 11135 10379 11141
rect 10321 11101 10333 11135
rect 10367 11132 10379 11135
rect 10597 11135 10655 11141
rect 10597 11132 10609 11135
rect 10367 11104 10609 11132
rect 10367 11101 10379 11104
rect 10321 11095 10379 11101
rect 10597 11101 10609 11104
rect 10643 11132 10655 11135
rect 10870 11132 10876 11144
rect 10643 11104 10876 11132
rect 10643 11101 10655 11104
rect 10597 11095 10655 11101
rect 10244 11064 10272 11095
rect 10870 11092 10876 11104
rect 10928 11092 10934 11144
rect 10962 11092 10968 11144
rect 11020 11132 11026 11144
rect 11057 11135 11115 11141
rect 11057 11132 11069 11135
rect 11020 11104 11069 11132
rect 11020 11092 11026 11104
rect 11057 11101 11069 11104
rect 11103 11101 11115 11135
rect 11057 11095 11115 11101
rect 11330 11092 11336 11144
rect 11388 11092 11394 11144
rect 12526 11092 12532 11144
rect 12584 11092 12590 11144
rect 12713 11135 12771 11141
rect 12713 11101 12725 11135
rect 12759 11101 12771 11135
rect 12820 11132 12848 11172
rect 12986 11160 12992 11212
rect 13044 11160 13050 11212
rect 14553 11203 14611 11209
rect 14553 11169 14565 11203
rect 14599 11200 14611 11203
rect 14918 11200 14924 11212
rect 14599 11172 14924 11200
rect 14599 11169 14611 11172
rect 14553 11163 14611 11169
rect 14918 11160 14924 11172
rect 14976 11160 14982 11212
rect 16025 11203 16083 11209
rect 16025 11169 16037 11203
rect 16071 11200 16083 11203
rect 16114 11200 16120 11212
rect 16071 11172 16120 11200
rect 16071 11169 16083 11172
rect 16025 11163 16083 11169
rect 16114 11160 16120 11172
rect 16172 11200 16178 11212
rect 16172 11172 18276 11200
rect 16172 11160 16178 11172
rect 15108 11144 15160 11150
rect 13081 11135 13139 11141
rect 13081 11132 13093 11135
rect 12820 11104 13093 11132
rect 12713 11095 12771 11101
rect 13081 11101 13093 11104
rect 13127 11101 13139 11135
rect 13081 11095 13139 11101
rect 11348 11064 11376 11092
rect 10244 11036 11376 11064
rect 11790 11024 11796 11076
rect 11848 11064 11854 11076
rect 12728 11064 12756 11095
rect 14182 11092 14188 11144
rect 14240 11132 14246 11144
rect 14461 11135 14519 11141
rect 14461 11132 14473 11135
rect 14240 11104 14473 11132
rect 14240 11092 14246 11104
rect 14461 11101 14473 11104
rect 14507 11132 14519 11135
rect 14826 11132 14832 11144
rect 14507 11104 14832 11132
rect 14507 11101 14519 11104
rect 14461 11095 14519 11101
rect 14826 11092 14832 11104
rect 14884 11132 14890 11144
rect 15013 11135 15071 11141
rect 15013 11132 15025 11135
rect 14884 11104 15025 11132
rect 14884 11092 14890 11104
rect 15013 11101 15025 11104
rect 15059 11101 15071 11135
rect 15013 11095 15071 11101
rect 17126 11092 17132 11144
rect 17184 11132 17190 11144
rect 17221 11135 17279 11141
rect 17221 11132 17233 11135
rect 17184 11104 17233 11132
rect 17184 11092 17190 11104
rect 17221 11101 17233 11104
rect 17267 11101 17279 11135
rect 17221 11095 17279 11101
rect 17405 11135 17463 11141
rect 17405 11101 17417 11135
rect 17451 11132 17463 11135
rect 17494 11132 17500 11144
rect 17451 11104 17500 11132
rect 17451 11101 17463 11104
rect 17405 11095 17463 11101
rect 17494 11092 17500 11104
rect 17552 11092 17558 11144
rect 17770 11141 17776 11144
rect 17752 11135 17776 11141
rect 17752 11132 17764 11135
rect 17600 11104 17764 11132
rect 15108 11086 15160 11092
rect 11848 11036 12756 11064
rect 11848 11024 11854 11036
rect 16206 11024 16212 11076
rect 16264 11064 16270 11076
rect 17600 11064 17628 11104
rect 17752 11101 17764 11104
rect 17752 11095 17776 11101
rect 17770 11092 17776 11095
rect 17828 11092 17834 11144
rect 18046 11132 18052 11144
rect 17972 11104 18052 11132
rect 16264 11036 17628 11064
rect 16264 11024 16270 11036
rect 10318 10996 10324 11008
rect 10152 10968 10324 10996
rect 9309 10959 9367 10965
rect 10318 10956 10324 10968
rect 10376 10996 10382 11008
rect 11149 10999 11207 11005
rect 11149 10996 11161 10999
rect 10376 10968 11161 10996
rect 10376 10956 10382 10968
rect 11149 10965 11161 10968
rect 11195 10965 11207 10999
rect 11149 10959 11207 10965
rect 12621 10999 12679 11005
rect 12621 10965 12633 10999
rect 12667 10996 12679 10999
rect 12710 10996 12716 11008
rect 12667 10968 12716 10996
rect 12667 10965 12679 10968
rect 12621 10959 12679 10965
rect 12710 10956 12716 10968
rect 12768 10956 12774 11008
rect 13906 10956 13912 11008
rect 13964 10956 13970 11008
rect 17681 10999 17739 11005
rect 17681 10965 17693 10999
rect 17727 10996 17739 10999
rect 17972 10996 18000 11104
rect 18046 11092 18052 11104
rect 18104 11092 18110 11144
rect 18248 11141 18276 11172
rect 23474 11160 23480 11212
rect 23532 11200 23538 11212
rect 23750 11200 23756 11212
rect 23532 11172 23756 11200
rect 23532 11160 23538 11172
rect 23750 11160 23756 11172
rect 23808 11200 23814 11212
rect 26068 11209 26096 11240
rect 27154 11228 27160 11240
rect 27212 11228 27218 11280
rect 26053 11203 26111 11209
rect 23808 11172 24716 11200
rect 23808 11160 23814 11172
rect 18233 11135 18291 11141
rect 18233 11101 18245 11135
rect 18279 11101 18291 11135
rect 18233 11095 18291 11101
rect 18598 11092 18604 11144
rect 18656 11132 18662 11144
rect 19245 11135 19303 11141
rect 19245 11132 19257 11135
rect 18656 11104 19257 11132
rect 18656 11092 18662 11104
rect 19245 11101 19257 11104
rect 19291 11101 19303 11135
rect 19245 11095 19303 11101
rect 19429 11135 19487 11141
rect 19429 11101 19441 11135
rect 19475 11132 19487 11135
rect 19886 11132 19892 11144
rect 19475 11104 19892 11132
rect 19475 11101 19487 11104
rect 19429 11095 19487 11101
rect 19886 11092 19892 11104
rect 19944 11092 19950 11144
rect 22370 11092 22376 11144
rect 22428 11092 22434 11144
rect 24489 11135 24547 11141
rect 24489 11101 24501 11135
rect 24535 11132 24547 11135
rect 24578 11132 24584 11144
rect 24535 11104 24584 11132
rect 24535 11101 24547 11104
rect 24489 11095 24547 11101
rect 24578 11092 24584 11104
rect 24636 11092 24642 11144
rect 24688 11141 24716 11172
rect 26053 11169 26065 11203
rect 26099 11169 26111 11203
rect 26053 11163 26111 11169
rect 26237 11203 26295 11209
rect 26237 11169 26249 11203
rect 26283 11200 26295 11203
rect 26602 11200 26608 11212
rect 26283 11172 26608 11200
rect 26283 11169 26295 11172
rect 26237 11163 26295 11169
rect 26602 11160 26608 11172
rect 26660 11200 26666 11212
rect 27246 11200 27252 11212
rect 26660 11172 27252 11200
rect 26660 11160 26666 11172
rect 27246 11160 27252 11172
rect 27304 11160 27310 11212
rect 24673 11135 24731 11141
rect 24673 11101 24685 11135
rect 24719 11101 24731 11135
rect 24673 11095 24731 11101
rect 25406 11092 25412 11144
rect 25464 11132 25470 11144
rect 25961 11135 26019 11141
rect 25961 11132 25973 11135
rect 25464 11104 25973 11132
rect 25464 11092 25470 11104
rect 25961 11101 25973 11104
rect 26007 11101 26019 11135
rect 25961 11095 26019 11101
rect 19061 11067 19119 11073
rect 19061 11033 19073 11067
rect 19107 11064 19119 11067
rect 19334 11064 19340 11076
rect 19107 11036 19340 11064
rect 19107 11033 19119 11036
rect 19061 11027 19119 11033
rect 19334 11024 19340 11036
rect 19392 11024 19398 11076
rect 21174 11024 21180 11076
rect 21232 11064 21238 11076
rect 22097 11067 22155 11073
rect 22097 11064 22109 11067
rect 21232 11036 22109 11064
rect 21232 11024 21238 11036
rect 22097 11033 22109 11036
rect 22143 11033 22155 11067
rect 22097 11027 22155 11033
rect 17727 10968 18000 10996
rect 19613 10999 19671 11005
rect 17727 10965 17739 10968
rect 17681 10959 17739 10965
rect 19613 10965 19625 10999
rect 19659 10996 19671 10999
rect 19794 10996 19800 11008
rect 19659 10968 19800 10996
rect 19659 10965 19671 10968
rect 19613 10959 19671 10965
rect 19794 10956 19800 10968
rect 19852 10956 19858 11008
rect 22278 10956 22284 11008
rect 22336 10956 22342 11008
rect 1104 10906 27876 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 27876 10906
rect 1104 10832 27876 10854
rect 3510 10752 3516 10804
rect 3568 10792 3574 10804
rect 12897 10795 12955 10801
rect 12897 10792 12909 10795
rect 3568 10764 4660 10792
rect 3568 10752 3574 10764
rect 3878 10684 3884 10736
rect 3936 10724 3942 10736
rect 3936 10696 4568 10724
rect 3936 10684 3942 10696
rect 4540 10665 4568 10696
rect 4632 10665 4660 10764
rect 12452 10764 12909 10792
rect 9030 10684 9036 10736
rect 9088 10724 9094 10736
rect 9401 10727 9459 10733
rect 9401 10724 9413 10727
rect 9088 10696 9413 10724
rect 9088 10684 9094 10696
rect 9401 10693 9413 10696
rect 9447 10693 9459 10727
rect 9401 10687 9459 10693
rect 12452 10668 12480 10764
rect 12897 10761 12909 10764
rect 12943 10761 12955 10795
rect 12897 10755 12955 10761
rect 18141 10795 18199 10801
rect 18141 10761 18153 10795
rect 18187 10792 18199 10795
rect 18598 10792 18604 10804
rect 18187 10764 18604 10792
rect 18187 10761 18199 10764
rect 18141 10755 18199 10761
rect 18598 10752 18604 10764
rect 18656 10752 18662 10804
rect 20346 10752 20352 10804
rect 20404 10792 20410 10804
rect 20641 10795 20699 10801
rect 20641 10792 20653 10795
rect 20404 10764 20653 10792
rect 20404 10752 20410 10764
rect 20641 10761 20653 10764
rect 20687 10761 20699 10795
rect 20641 10755 20699 10761
rect 20809 10795 20867 10801
rect 20809 10761 20821 10795
rect 20855 10792 20867 10795
rect 20898 10792 20904 10804
rect 20855 10764 20904 10792
rect 20855 10761 20867 10764
rect 20809 10755 20867 10761
rect 20898 10752 20904 10764
rect 20956 10792 20962 10804
rect 22189 10795 22247 10801
rect 20956 10764 21036 10792
rect 20956 10752 20962 10764
rect 13081 10727 13139 10733
rect 13081 10724 13093 10727
rect 12728 10696 13093 10724
rect 12728 10668 12756 10696
rect 13081 10693 13093 10696
rect 13127 10693 13139 10727
rect 13081 10687 13139 10693
rect 17221 10727 17279 10733
rect 17221 10693 17233 10727
rect 17267 10724 17279 10727
rect 17267 10696 17632 10724
rect 17267 10693 17279 10696
rect 17221 10687 17279 10693
rect 4525 10659 4583 10665
rect 3818 10628 4292 10656
rect 3329 10591 3387 10597
rect 3329 10557 3341 10591
rect 3375 10557 3387 10591
rect 3329 10551 3387 10557
rect 3344 10520 3372 10551
rect 4154 10548 4160 10600
rect 4212 10548 4218 10600
rect 4264 10597 4292 10628
rect 4525 10625 4537 10659
rect 4571 10625 4583 10659
rect 4525 10619 4583 10625
rect 4617 10659 4675 10665
rect 4617 10625 4629 10659
rect 4663 10625 4675 10659
rect 4617 10619 4675 10625
rect 4798 10616 4804 10668
rect 4856 10656 4862 10668
rect 4893 10659 4951 10665
rect 4893 10656 4905 10659
rect 4856 10628 4905 10656
rect 4856 10616 4862 10628
rect 4893 10625 4905 10628
rect 4939 10625 4951 10659
rect 4893 10619 4951 10625
rect 5077 10659 5135 10665
rect 5077 10625 5089 10659
rect 5123 10656 5135 10659
rect 5258 10656 5264 10668
rect 5123 10628 5264 10656
rect 5123 10625 5135 10628
rect 5077 10619 5135 10625
rect 5258 10616 5264 10628
rect 5316 10616 5322 10668
rect 6638 10616 6644 10668
rect 6696 10616 6702 10668
rect 7466 10616 7472 10668
rect 7524 10656 7530 10668
rect 7653 10659 7711 10665
rect 7653 10656 7665 10659
rect 7524 10628 7665 10656
rect 7524 10616 7530 10628
rect 7653 10625 7665 10628
rect 7699 10625 7711 10659
rect 7653 10619 7711 10625
rect 9122 10616 9128 10668
rect 9180 10616 9186 10668
rect 9306 10616 9312 10668
rect 9364 10616 9370 10668
rect 9490 10616 9496 10668
rect 9548 10616 9554 10668
rect 12342 10616 12348 10668
rect 12400 10616 12406 10668
rect 12434 10616 12440 10668
rect 12492 10616 12498 10668
rect 12618 10616 12624 10668
rect 12676 10616 12682 10668
rect 12710 10616 12716 10668
rect 12768 10616 12774 10668
rect 12805 10659 12863 10665
rect 12805 10625 12817 10659
rect 12851 10625 12863 10659
rect 12805 10619 12863 10625
rect 4249 10591 4307 10597
rect 4249 10557 4261 10591
rect 4295 10557 4307 10591
rect 4249 10551 4307 10557
rect 4433 10591 4491 10597
rect 4433 10557 4445 10591
rect 4479 10557 4491 10591
rect 4433 10551 4491 10557
rect 4709 10591 4767 10597
rect 4709 10557 4721 10591
rect 4755 10588 4767 10591
rect 5350 10588 5356 10600
rect 4755 10560 5356 10588
rect 4755 10557 4767 10560
rect 4709 10551 4767 10557
rect 4338 10520 4344 10532
rect 3344 10492 4344 10520
rect 4338 10480 4344 10492
rect 4396 10480 4402 10532
rect 4448 10520 4476 10551
rect 5350 10548 5356 10560
rect 5408 10548 5414 10600
rect 6270 10548 6276 10600
rect 6328 10588 6334 10600
rect 6549 10591 6607 10597
rect 6549 10588 6561 10591
rect 6328 10560 6561 10588
rect 6328 10548 6334 10560
rect 6549 10557 6561 10560
rect 6595 10557 6607 10591
rect 6549 10551 6607 10557
rect 7377 10591 7435 10597
rect 7377 10557 7389 10591
rect 7423 10588 7435 10591
rect 8386 10588 8392 10600
rect 7423 10560 8392 10588
rect 7423 10557 7435 10560
rect 7377 10551 7435 10557
rect 8386 10548 8392 10560
rect 8444 10548 8450 10600
rect 12360 10588 12388 10616
rect 12820 10588 12848 10619
rect 15470 10616 15476 10668
rect 15528 10656 15534 10668
rect 16117 10659 16175 10665
rect 16117 10656 16129 10659
rect 15528 10628 16129 10656
rect 15528 10616 15534 10628
rect 16117 10625 16129 10628
rect 16163 10625 16175 10659
rect 16117 10619 16175 10625
rect 16206 10616 16212 10668
rect 16264 10656 16270 10668
rect 16301 10659 16359 10665
rect 16301 10656 16313 10659
rect 16264 10628 16313 10656
rect 16264 10616 16270 10628
rect 16301 10625 16313 10628
rect 16347 10625 16359 10659
rect 16301 10619 16359 10625
rect 16482 10616 16488 10668
rect 16540 10656 16546 10668
rect 16853 10659 16911 10665
rect 16853 10656 16865 10659
rect 16540 10628 16865 10656
rect 16540 10616 16546 10628
rect 16853 10625 16865 10628
rect 16899 10625 16911 10659
rect 16853 10619 16911 10625
rect 17034 10616 17040 10668
rect 17092 10616 17098 10668
rect 17313 10659 17371 10665
rect 17313 10625 17325 10659
rect 17359 10625 17371 10659
rect 17313 10619 17371 10625
rect 12360 10560 12848 10588
rect 15378 10548 15384 10600
rect 15436 10588 15442 10600
rect 16224 10588 16252 10616
rect 15436 10560 16252 10588
rect 15436 10548 15442 10560
rect 16758 10548 16764 10600
rect 16816 10588 16822 10600
rect 17328 10588 17356 10619
rect 16816 10560 17356 10588
rect 17604 10588 17632 10696
rect 17770 10684 17776 10736
rect 17828 10733 17834 10736
rect 17828 10727 17857 10733
rect 17845 10693 17857 10727
rect 17828 10687 17857 10693
rect 17828 10684 17834 10687
rect 17954 10684 17960 10736
rect 18012 10733 18018 10736
rect 18012 10727 18031 10733
rect 18019 10693 18031 10727
rect 18012 10687 18031 10693
rect 18012 10684 18018 10687
rect 19702 10684 19708 10736
rect 19760 10724 19766 10736
rect 19981 10727 20039 10733
rect 19981 10724 19993 10727
rect 19760 10696 19993 10724
rect 19760 10684 19766 10696
rect 19981 10693 19993 10696
rect 20027 10693 20039 10727
rect 20181 10727 20239 10733
rect 20181 10724 20193 10727
rect 19981 10687 20039 10693
rect 20180 10693 20193 10724
rect 20227 10693 20239 10727
rect 20180 10687 20239 10693
rect 20441 10727 20499 10733
rect 20441 10693 20453 10727
rect 20487 10693 20499 10727
rect 20441 10687 20499 10693
rect 17678 10616 17684 10668
rect 17736 10616 17742 10668
rect 19613 10659 19671 10665
rect 19613 10625 19625 10659
rect 19659 10656 19671 10659
rect 19794 10656 19800 10668
rect 19659 10628 19800 10656
rect 19659 10625 19671 10628
rect 19613 10619 19671 10625
rect 19794 10616 19800 10628
rect 19852 10656 19858 10668
rect 20180 10656 20208 10687
rect 20456 10656 20484 10687
rect 19852 10628 20484 10656
rect 19852 10616 19858 10628
rect 20530 10616 20536 10668
rect 20588 10656 20594 10668
rect 21008 10665 21036 10764
rect 22189 10761 22201 10795
rect 22235 10792 22247 10795
rect 22235 10764 22784 10792
rect 22235 10761 22247 10764
rect 22189 10755 22247 10761
rect 20901 10659 20959 10665
rect 20901 10656 20913 10659
rect 20588 10628 20913 10656
rect 20588 10616 20594 10628
rect 20901 10625 20913 10628
rect 20947 10625 20959 10659
rect 20901 10619 20959 10625
rect 20993 10659 21051 10665
rect 20993 10625 21005 10659
rect 21039 10625 21051 10659
rect 20993 10619 21051 10625
rect 21082 10616 21088 10668
rect 21140 10656 21146 10668
rect 21450 10656 21456 10668
rect 21140 10628 21456 10656
rect 21140 10616 21146 10628
rect 21450 10616 21456 10628
rect 21508 10616 21514 10668
rect 22002 10616 22008 10668
rect 22060 10616 22066 10668
rect 22186 10616 22192 10668
rect 22244 10656 22250 10668
rect 22281 10659 22339 10665
rect 22281 10656 22293 10659
rect 22244 10628 22293 10656
rect 22244 10616 22250 10628
rect 22281 10625 22293 10628
rect 22327 10625 22339 10659
rect 22281 10619 22339 10625
rect 22465 10659 22523 10665
rect 22465 10625 22477 10659
rect 22511 10656 22523 10659
rect 22554 10656 22560 10668
rect 22511 10628 22560 10656
rect 22511 10625 22523 10628
rect 22465 10619 22523 10625
rect 22554 10616 22560 10628
rect 22612 10616 22618 10668
rect 22756 10665 22784 10764
rect 22925 10727 22983 10733
rect 22925 10693 22937 10727
rect 22971 10724 22983 10727
rect 22971 10696 24532 10724
rect 22971 10693 22983 10696
rect 22925 10687 22983 10693
rect 24504 10668 24532 10696
rect 25682 10684 25688 10736
rect 25740 10684 25746 10736
rect 22741 10659 22799 10665
rect 22741 10625 22753 10659
rect 22787 10656 22799 10659
rect 24210 10656 24216 10668
rect 22787 10628 24216 10656
rect 22787 10625 22799 10628
rect 22741 10619 22799 10625
rect 24210 10616 24216 10628
rect 24268 10616 24274 10668
rect 24302 10616 24308 10668
rect 24360 10616 24366 10668
rect 24486 10616 24492 10668
rect 24544 10616 24550 10668
rect 24670 10616 24676 10668
rect 24728 10616 24734 10668
rect 17604 10560 18138 10588
rect 16816 10548 16822 10560
rect 4985 10523 5043 10529
rect 4985 10520 4997 10523
rect 4448 10492 4997 10520
rect 4632 10464 4660 10492
rect 4985 10489 4997 10492
rect 5031 10489 5043 10523
rect 4985 10483 5043 10489
rect 12986 10480 12992 10532
rect 13044 10520 13050 10532
rect 13081 10523 13139 10529
rect 13081 10520 13093 10523
rect 13044 10492 13093 10520
rect 13044 10480 13050 10492
rect 13081 10489 13093 10492
rect 13127 10489 13139 10523
rect 13081 10483 13139 10489
rect 16117 10523 16175 10529
rect 16117 10489 16129 10523
rect 16163 10520 16175 10523
rect 17310 10520 17316 10532
rect 16163 10492 17316 10520
rect 16163 10489 16175 10492
rect 16117 10483 16175 10489
rect 17310 10480 17316 10492
rect 17368 10480 17374 10532
rect 4614 10412 4620 10464
rect 4672 10412 4678 10464
rect 7190 10412 7196 10464
rect 7248 10452 7254 10464
rect 7745 10455 7803 10461
rect 7745 10452 7757 10455
rect 7248 10424 7757 10452
rect 7248 10412 7254 10424
rect 7745 10421 7757 10424
rect 7791 10421 7803 10455
rect 7745 10415 7803 10421
rect 9677 10455 9735 10461
rect 9677 10421 9689 10455
rect 9723 10452 9735 10455
rect 9858 10452 9864 10464
rect 9723 10424 9864 10452
rect 9723 10421 9735 10424
rect 9677 10415 9735 10421
rect 9858 10412 9864 10424
rect 9916 10412 9922 10464
rect 11790 10412 11796 10464
rect 11848 10452 11854 10464
rect 12161 10455 12219 10461
rect 12161 10452 12173 10455
rect 11848 10424 12173 10452
rect 11848 10412 11854 10424
rect 12161 10421 12173 10424
rect 12207 10421 12219 10455
rect 12161 10415 12219 10421
rect 17494 10412 17500 10464
rect 17552 10452 17558 10464
rect 17917 10455 17975 10461
rect 17917 10452 17929 10455
rect 17552 10424 17929 10452
rect 17552 10412 17558 10424
rect 17917 10421 17929 10424
rect 17963 10421 17975 10455
rect 18110 10452 18138 10560
rect 19334 10548 19340 10600
rect 19392 10588 19398 10600
rect 19429 10591 19487 10597
rect 19429 10588 19441 10591
rect 19392 10560 19441 10588
rect 19392 10548 19398 10560
rect 19429 10557 19441 10560
rect 19475 10588 19487 10591
rect 19886 10588 19892 10600
rect 19475 10560 19892 10588
rect 19475 10557 19487 10560
rect 19429 10551 19487 10557
rect 19886 10548 19892 10560
rect 19944 10588 19950 10600
rect 19944 10560 20208 10588
rect 19944 10548 19950 10560
rect 20180 10520 20208 10560
rect 20548 10520 20576 10616
rect 21174 10548 21180 10600
rect 21232 10548 21238 10600
rect 21818 10548 21824 10600
rect 21876 10548 21882 10600
rect 22649 10591 22707 10597
rect 22649 10557 22661 10591
rect 22695 10588 22707 10591
rect 22830 10588 22836 10600
rect 22695 10560 22836 10588
rect 22695 10557 22707 10560
rect 22649 10551 22707 10557
rect 22830 10548 22836 10560
rect 22888 10548 22894 10600
rect 24397 10591 24455 10597
rect 24397 10557 24409 10591
rect 24443 10588 24455 10591
rect 24780 10588 24808 10642
rect 24443 10560 24808 10588
rect 24443 10557 24455 10560
rect 24397 10551 24455 10557
rect 20180 10492 20576 10520
rect 21085 10523 21143 10529
rect 19518 10452 19524 10464
rect 18110 10424 19524 10452
rect 17917 10415 17975 10421
rect 19518 10412 19524 10424
rect 19576 10412 19582 10464
rect 19797 10455 19855 10461
rect 19797 10421 19809 10455
rect 19843 10452 19855 10455
rect 19978 10452 19984 10464
rect 19843 10424 19984 10452
rect 19843 10421 19855 10424
rect 19797 10415 19855 10421
rect 19978 10412 19984 10424
rect 20036 10412 20042 10464
rect 20180 10461 20208 10492
rect 21085 10489 21097 10523
rect 21131 10520 21143 10523
rect 22557 10523 22615 10529
rect 22557 10520 22569 10523
rect 21131 10492 22569 10520
rect 21131 10489 21143 10492
rect 21085 10483 21143 10489
rect 22557 10489 22569 10492
rect 22603 10489 22615 10523
rect 22557 10483 22615 10489
rect 20165 10455 20223 10461
rect 20165 10421 20177 10455
rect 20211 10421 20223 10455
rect 20165 10415 20223 10421
rect 20349 10455 20407 10461
rect 20349 10421 20361 10455
rect 20395 10452 20407 10455
rect 20438 10452 20444 10464
rect 20395 10424 20444 10452
rect 20395 10421 20407 10424
rect 20349 10415 20407 10421
rect 20438 10412 20444 10424
rect 20496 10412 20502 10464
rect 20622 10412 20628 10464
rect 20680 10412 20686 10464
rect 21634 10412 21640 10464
rect 21692 10452 21698 10464
rect 22278 10452 22284 10464
rect 21692 10424 22284 10452
rect 21692 10412 21698 10424
rect 22278 10412 22284 10424
rect 22336 10412 22342 10464
rect 1104 10362 27876 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 27876 10362
rect 1104 10288 27876 10310
rect 6270 10208 6276 10260
rect 6328 10208 6334 10260
rect 11882 10208 11888 10260
rect 11940 10208 11946 10260
rect 15013 10251 15071 10257
rect 15013 10217 15025 10251
rect 15059 10248 15071 10251
rect 15102 10248 15108 10260
rect 15059 10220 15108 10248
rect 15059 10217 15071 10220
rect 15013 10211 15071 10217
rect 15102 10208 15108 10220
rect 15160 10208 15166 10260
rect 15470 10208 15476 10260
rect 15528 10208 15534 10260
rect 16025 10251 16083 10257
rect 16025 10248 16037 10251
rect 15580 10220 16037 10248
rect 15580 10124 15608 10220
rect 16025 10217 16037 10220
rect 16071 10217 16083 10251
rect 16025 10211 16083 10217
rect 16040 10180 16068 10211
rect 16758 10208 16764 10260
rect 16816 10208 16822 10260
rect 16853 10251 16911 10257
rect 16853 10217 16865 10251
rect 16899 10248 16911 10251
rect 17034 10248 17040 10260
rect 16899 10220 17040 10248
rect 16899 10217 16911 10220
rect 16853 10211 16911 10217
rect 17034 10208 17040 10220
rect 17092 10208 17098 10260
rect 19518 10208 19524 10260
rect 19576 10248 19582 10260
rect 21266 10248 21272 10260
rect 19576 10220 21272 10248
rect 19576 10208 19582 10220
rect 21266 10208 21272 10220
rect 21324 10248 21330 10260
rect 21361 10251 21419 10257
rect 21361 10248 21373 10251
rect 21324 10220 21373 10248
rect 21324 10208 21330 10220
rect 21361 10217 21373 10220
rect 21407 10217 21419 10251
rect 21361 10211 21419 10217
rect 21818 10208 21824 10260
rect 21876 10248 21882 10260
rect 21876 10220 22140 10248
rect 21876 10208 21882 10220
rect 17497 10183 17555 10189
rect 16040 10152 16252 10180
rect 5534 10112 5540 10124
rect 5460 10084 5540 10112
rect 4706 10004 4712 10056
rect 4764 10044 4770 10056
rect 5460 10053 5488 10084
rect 5534 10072 5540 10084
rect 5592 10112 5598 10124
rect 7466 10112 7472 10124
rect 5592 10084 7472 10112
rect 5592 10072 5598 10084
rect 5445 10047 5503 10053
rect 5445 10044 5457 10047
rect 4764 10016 5457 10044
rect 4764 10004 4770 10016
rect 5445 10013 5457 10016
rect 5491 10013 5503 10047
rect 5445 10007 5503 10013
rect 5629 10047 5687 10053
rect 5629 10013 5641 10047
rect 5675 10013 5687 10047
rect 5629 10007 5687 10013
rect 5721 10047 5779 10053
rect 5721 10013 5733 10047
rect 5767 10044 5779 10047
rect 5902 10044 5908 10056
rect 5767 10016 5908 10044
rect 5767 10013 5779 10016
rect 5721 10007 5779 10013
rect 5644 9976 5672 10007
rect 5902 10004 5908 10016
rect 5960 10004 5966 10056
rect 6472 10053 6500 10084
rect 7466 10072 7472 10084
rect 7524 10072 7530 10124
rect 9306 10072 9312 10124
rect 9364 10072 9370 10124
rect 14292 10084 15516 10112
rect 6457 10047 6515 10053
rect 6457 10013 6469 10047
rect 6503 10013 6515 10047
rect 6457 10007 6515 10013
rect 6822 10004 6828 10056
rect 6880 10004 6886 10056
rect 8021 10047 8079 10053
rect 8021 10013 8033 10047
rect 8067 10013 8079 10047
rect 8021 10007 8079 10013
rect 6178 9976 6184 9988
rect 5644 9948 6184 9976
rect 6178 9936 6184 9948
rect 6236 9976 6242 9988
rect 6546 9976 6552 9988
rect 6236 9948 6552 9976
rect 6236 9936 6242 9948
rect 6546 9936 6552 9948
rect 6604 9936 6610 9988
rect 6638 9936 6644 9988
rect 6696 9936 6702 9988
rect 8036 9976 8064 10007
rect 8202 10004 8208 10056
rect 8260 10044 8266 10056
rect 9217 10047 9275 10053
rect 9217 10044 9229 10047
rect 8260 10016 9229 10044
rect 8260 10004 8266 10016
rect 9217 10013 9229 10016
rect 9263 10013 9275 10047
rect 9217 10007 9275 10013
rect 9490 10004 9496 10056
rect 9548 10044 9554 10056
rect 10413 10047 10471 10053
rect 10413 10044 10425 10047
rect 9548 10016 10425 10044
rect 9548 10004 9554 10016
rect 10413 10013 10425 10016
rect 10459 10013 10471 10047
rect 10413 10007 10471 10013
rect 10778 10004 10784 10056
rect 10836 10004 10842 10056
rect 13906 10004 13912 10056
rect 13964 10044 13970 10056
rect 14292 10053 14320 10084
rect 14277 10047 14335 10053
rect 14277 10044 14289 10047
rect 13964 10016 14289 10044
rect 13964 10004 13970 10016
rect 14277 10013 14289 10016
rect 14323 10013 14335 10047
rect 14277 10007 14335 10013
rect 14366 10004 14372 10056
rect 14424 10044 14430 10056
rect 14553 10047 14611 10053
rect 14553 10044 14565 10047
rect 14424 10016 14565 10044
rect 14424 10004 14430 10016
rect 14553 10013 14565 10016
rect 14599 10013 14611 10047
rect 14553 10007 14611 10013
rect 15194 10004 15200 10056
rect 15252 10004 15258 10056
rect 15378 10004 15384 10056
rect 15436 10004 15442 10056
rect 15488 10044 15516 10084
rect 15562 10072 15568 10124
rect 15620 10072 15626 10124
rect 16114 10072 16120 10124
rect 16172 10072 16178 10124
rect 15749 10047 15807 10053
rect 15749 10044 15761 10047
rect 15488 10016 15761 10044
rect 15749 10013 15761 10016
rect 15795 10013 15807 10047
rect 15749 10007 15807 10013
rect 16022 10004 16028 10056
rect 16080 10004 16086 10056
rect 16224 10044 16252 10152
rect 17497 10149 17509 10183
rect 17543 10180 17555 10183
rect 17678 10180 17684 10192
rect 17543 10152 17684 10180
rect 17543 10149 17555 10152
rect 17497 10143 17555 10149
rect 17678 10140 17684 10152
rect 17736 10180 17742 10192
rect 18509 10183 18567 10189
rect 17736 10152 18092 10180
rect 17736 10140 17742 10152
rect 18064 10121 18092 10152
rect 18509 10149 18521 10183
rect 18555 10180 18567 10183
rect 19702 10180 19708 10192
rect 18555 10152 19708 10180
rect 18555 10149 18567 10152
rect 18509 10143 18567 10149
rect 19702 10140 19708 10152
rect 19760 10140 19766 10192
rect 20947 10183 21005 10189
rect 20947 10149 20959 10183
rect 20993 10180 21005 10183
rect 21082 10180 21088 10192
rect 20993 10152 21088 10180
rect 20993 10149 21005 10152
rect 20947 10143 21005 10149
rect 21082 10140 21088 10152
rect 21140 10140 21146 10192
rect 21177 10183 21235 10189
rect 21177 10149 21189 10183
rect 21223 10180 21235 10183
rect 22002 10180 22008 10192
rect 21223 10152 22008 10180
rect 21223 10149 21235 10152
rect 21177 10143 21235 10149
rect 22002 10140 22008 10152
rect 22060 10140 22066 10192
rect 18049 10115 18107 10121
rect 16776 10084 17908 10112
rect 16482 10044 16488 10056
rect 16224 10016 16488 10044
rect 16482 10004 16488 10016
rect 16540 10044 16546 10056
rect 16776 10053 16804 10084
rect 16577 10047 16635 10053
rect 16577 10044 16589 10047
rect 16540 10016 16589 10044
rect 16540 10004 16546 10016
rect 16577 10013 16589 10016
rect 16623 10013 16635 10047
rect 16577 10007 16635 10013
rect 16761 10047 16819 10053
rect 16761 10013 16773 10047
rect 16807 10013 16819 10047
rect 16761 10007 16819 10013
rect 8294 9976 8300 9988
rect 8036 9948 8300 9976
rect 8294 9936 8300 9948
rect 8352 9976 8358 9988
rect 8754 9976 8760 9988
rect 8352 9948 8760 9976
rect 8352 9936 8358 9948
rect 8754 9936 8760 9948
rect 8812 9936 8818 9988
rect 5261 9911 5319 9917
rect 5261 9877 5273 9911
rect 5307 9908 5319 9911
rect 5350 9908 5356 9920
rect 5307 9880 5356 9908
rect 5307 9877 5319 9880
rect 5261 9871 5319 9877
rect 5350 9868 5356 9880
rect 5408 9868 5414 9920
rect 5810 9868 5816 9920
rect 5868 9868 5874 9920
rect 7466 9868 7472 9920
rect 7524 9908 7530 9920
rect 7837 9911 7895 9917
rect 7837 9908 7849 9911
rect 7524 9880 7849 9908
rect 7524 9868 7530 9880
rect 7837 9877 7849 9880
rect 7883 9908 7895 9911
rect 8110 9908 8116 9920
rect 7883 9880 8116 9908
rect 7883 9877 7895 9880
rect 7837 9871 7895 9877
rect 8110 9868 8116 9880
rect 8168 9868 8174 9920
rect 8202 9868 8208 9920
rect 8260 9908 8266 9920
rect 9508 9908 9536 10004
rect 14737 9979 14795 9985
rect 14737 9945 14749 9979
rect 14783 9976 14795 9979
rect 14918 9976 14924 9988
rect 14783 9948 14924 9976
rect 14783 9945 14795 9948
rect 14737 9939 14795 9945
rect 14918 9936 14924 9948
rect 14976 9936 14982 9988
rect 15289 9979 15347 9985
rect 15289 9945 15301 9979
rect 15335 9976 15347 9979
rect 15473 9979 15531 9985
rect 15473 9976 15485 9979
rect 15335 9948 15485 9976
rect 15335 9945 15347 9948
rect 15289 9939 15347 9945
rect 15473 9945 15485 9948
rect 15519 9945 15531 9979
rect 16040 9976 16068 10004
rect 16776 9976 16804 10007
rect 17034 10004 17040 10056
rect 17092 10004 17098 10056
rect 17129 10047 17187 10053
rect 17129 10013 17141 10047
rect 17175 10044 17187 10047
rect 17218 10044 17224 10056
rect 17175 10016 17224 10044
rect 17175 10013 17187 10016
rect 17129 10007 17187 10013
rect 17218 10004 17224 10016
rect 17276 10004 17282 10056
rect 17310 10004 17316 10056
rect 17368 10004 17374 10056
rect 17420 10053 17448 10084
rect 17405 10047 17463 10053
rect 17405 10013 17417 10047
rect 17451 10013 17463 10047
rect 17773 10047 17831 10053
rect 17773 10044 17785 10047
rect 17405 10007 17463 10013
rect 17604 10016 17785 10044
rect 16040 9948 16804 9976
rect 15473 9939 15531 9945
rect 8260 9880 9536 9908
rect 8260 9868 8266 9880
rect 10042 9868 10048 9920
rect 10100 9868 10106 9920
rect 14090 9868 14096 9920
rect 14148 9868 14154 9920
rect 14458 9868 14464 9920
rect 14516 9868 14522 9920
rect 15933 9911 15991 9917
rect 15933 9877 15945 9911
rect 15979 9908 15991 9911
rect 16206 9908 16212 9920
rect 15979 9880 16212 9908
rect 15979 9877 15991 9880
rect 15933 9871 15991 9877
rect 16206 9868 16212 9880
rect 16264 9868 16270 9920
rect 16390 9868 16396 9920
rect 16448 9868 16454 9920
rect 17052 9908 17080 10004
rect 17328 9976 17356 10004
rect 17497 9979 17555 9985
rect 17497 9976 17509 9979
rect 17328 9948 17509 9976
rect 17497 9945 17509 9948
rect 17543 9945 17555 9979
rect 17497 9939 17555 9945
rect 17604 9920 17632 10016
rect 17773 10013 17785 10016
rect 17819 10013 17831 10047
rect 17880 10044 17908 10084
rect 18049 10081 18061 10115
rect 18095 10081 18107 10115
rect 18049 10075 18107 10081
rect 19978 10072 19984 10124
rect 20036 10072 20042 10124
rect 20622 10112 20628 10124
rect 20180 10084 20628 10112
rect 20180 10056 20208 10084
rect 20622 10072 20628 10084
rect 20680 10072 20686 10124
rect 20824 10084 21404 10112
rect 18141 10047 18199 10053
rect 18141 10044 18153 10047
rect 17880 10016 18153 10044
rect 17773 10007 17831 10013
rect 18141 10013 18153 10016
rect 18187 10013 18199 10047
rect 18141 10007 18199 10013
rect 19702 10004 19708 10056
rect 19760 10004 19766 10056
rect 20162 10004 20168 10056
rect 20220 10004 20226 10056
rect 20346 10004 20352 10056
rect 20404 10004 20410 10056
rect 20438 10004 20444 10056
rect 20496 10044 20502 10056
rect 20824 10053 20852 10084
rect 20809 10047 20867 10053
rect 20809 10044 20821 10047
rect 20496 10016 20821 10044
rect 20496 10004 20502 10016
rect 20809 10013 20821 10016
rect 20855 10013 20867 10047
rect 20809 10007 20867 10013
rect 21082 10004 21088 10056
rect 21140 10004 21146 10056
rect 21266 10004 21272 10056
rect 21324 10004 21330 10056
rect 21376 10044 21404 10084
rect 21450 10072 21456 10124
rect 21508 10072 21514 10124
rect 21634 10044 21640 10056
rect 21376 10016 21640 10044
rect 21634 10004 21640 10016
rect 21692 10004 21698 10056
rect 22021 10053 22049 10140
rect 21920 10047 21978 10053
rect 21920 10013 21932 10047
rect 21966 10013 21978 10047
rect 21920 10007 21978 10013
rect 22006 10047 22064 10053
rect 22006 10013 22018 10047
rect 22052 10013 22064 10047
rect 22112 10044 22140 10220
rect 22554 10208 22560 10260
rect 22612 10208 22618 10260
rect 25958 10208 25964 10260
rect 26016 10208 26022 10260
rect 26326 10208 26332 10260
rect 26384 10208 26390 10260
rect 26418 10208 26424 10260
rect 26476 10208 26482 10260
rect 23845 10183 23903 10189
rect 23845 10149 23857 10183
rect 23891 10180 23903 10183
rect 24394 10180 24400 10192
rect 23891 10152 24400 10180
rect 23891 10149 23903 10152
rect 23845 10143 23903 10149
rect 24394 10140 24400 10152
rect 24452 10140 24458 10192
rect 25682 10140 25688 10192
rect 25740 10180 25746 10192
rect 25740 10152 26648 10180
rect 25740 10140 25746 10152
rect 23566 10072 23572 10124
rect 23624 10072 23630 10124
rect 25516 10084 26096 10112
rect 25516 10056 25544 10084
rect 22189 10047 22247 10053
rect 22189 10044 22201 10047
rect 22112 10016 22201 10044
rect 22006 10007 22064 10013
rect 22189 10013 22201 10016
rect 22235 10013 22247 10047
rect 22189 10007 22247 10013
rect 19797 9979 19855 9985
rect 19797 9945 19809 9979
rect 19843 9976 19855 9979
rect 21174 9976 21180 9988
rect 19843 9948 21180 9976
rect 19843 9945 19855 9948
rect 19797 9939 19855 9945
rect 21174 9936 21180 9948
rect 21232 9936 21238 9988
rect 21358 9936 21364 9988
rect 21416 9936 21422 9988
rect 17586 9908 17592 9920
rect 17052 9880 17592 9908
rect 17586 9868 17592 9880
rect 17644 9868 17650 9920
rect 17678 9868 17684 9920
rect 17736 9868 17742 9920
rect 21192 9908 21220 9936
rect 21928 9908 21956 10007
rect 22278 10004 22284 10056
rect 22336 10004 22342 10056
rect 22370 10004 22376 10056
rect 22428 10053 22434 10056
rect 22428 10007 22436 10053
rect 22428 10004 22434 10007
rect 23474 10004 23480 10056
rect 23532 10004 23538 10056
rect 23934 10004 23940 10056
rect 23992 10004 23998 10056
rect 24121 10047 24179 10053
rect 24121 10013 24133 10047
rect 24167 10013 24179 10047
rect 24121 10007 24179 10013
rect 21192 9880 21956 9908
rect 22094 9868 22100 9920
rect 22152 9908 22158 9920
rect 22388 9908 22416 10004
rect 22922 9936 22928 9988
rect 22980 9976 22986 9988
rect 24136 9976 24164 10007
rect 25498 10004 25504 10056
rect 25556 10004 25562 10056
rect 25682 10004 25688 10056
rect 25740 10044 25746 10056
rect 26068 10053 26096 10084
rect 26418 10072 26424 10124
rect 26476 10072 26482 10124
rect 26620 10112 26648 10152
rect 26620 10084 26740 10112
rect 25777 10047 25835 10053
rect 25777 10044 25789 10047
rect 25740 10016 25789 10044
rect 25740 10004 25746 10016
rect 25777 10013 25789 10016
rect 25823 10013 25835 10047
rect 25777 10007 25835 10013
rect 26053 10047 26111 10053
rect 26053 10013 26065 10047
rect 26099 10013 26111 10047
rect 26053 10007 26111 10013
rect 26329 10047 26387 10053
rect 26329 10013 26341 10047
rect 26375 10044 26387 10047
rect 26436 10044 26464 10072
rect 26375 10016 26464 10044
rect 26375 10013 26387 10016
rect 26329 10007 26387 10013
rect 22980 9948 24164 9976
rect 26068 9976 26096 10007
rect 26510 10004 26516 10056
rect 26568 10044 26574 10056
rect 26712 10053 26740 10084
rect 26605 10047 26663 10053
rect 26605 10044 26617 10047
rect 26568 10016 26617 10044
rect 26568 10004 26574 10016
rect 26605 10013 26617 10016
rect 26651 10013 26663 10047
rect 26605 10007 26663 10013
rect 26697 10047 26755 10053
rect 26697 10013 26709 10047
rect 26743 10013 26755 10047
rect 26697 10007 26755 10013
rect 26421 9979 26479 9985
rect 26421 9976 26433 9979
rect 26068 9948 26433 9976
rect 22980 9936 22986 9948
rect 26421 9945 26433 9948
rect 26467 9945 26479 9979
rect 26421 9939 26479 9945
rect 22152 9880 22416 9908
rect 22152 9868 22158 9880
rect 24026 9868 24032 9920
rect 24084 9868 24090 9920
rect 25593 9911 25651 9917
rect 25593 9877 25605 9911
rect 25639 9908 25651 9911
rect 26145 9911 26203 9917
rect 26145 9908 26157 9911
rect 25639 9880 26157 9908
rect 25639 9877 25651 9880
rect 25593 9871 25651 9877
rect 26145 9877 26157 9880
rect 26191 9908 26203 9911
rect 26528 9908 26556 10004
rect 26191 9880 26556 9908
rect 26191 9877 26203 9880
rect 26145 9871 26203 9877
rect 1104 9818 27876 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 27876 9818
rect 1104 9744 27876 9766
rect 3712 9676 3924 9704
rect 3589 9639 3647 9645
rect 3589 9605 3601 9639
rect 3635 9636 3647 9639
rect 3712 9636 3740 9676
rect 3635 9608 3740 9636
rect 3789 9639 3847 9645
rect 3635 9605 3647 9608
rect 3589 9599 3647 9605
rect 3789 9605 3801 9639
rect 3835 9605 3847 9639
rect 3896 9636 3924 9676
rect 4706 9664 4712 9716
rect 4764 9704 4770 9716
rect 5350 9704 5356 9716
rect 4764 9676 5356 9704
rect 4764 9664 4770 9676
rect 5350 9664 5356 9676
rect 5408 9704 5414 9716
rect 8202 9704 8208 9716
rect 5408 9676 8208 9704
rect 5408 9664 5414 9676
rect 8202 9664 8208 9676
rect 8260 9664 8266 9716
rect 9306 9664 9312 9716
rect 9364 9664 9370 9716
rect 17218 9664 17224 9716
rect 17276 9704 17282 9716
rect 17678 9704 17684 9716
rect 17276 9676 17684 9704
rect 17276 9664 17282 9676
rect 17678 9664 17684 9676
rect 17736 9664 17742 9716
rect 23477 9707 23535 9713
rect 23477 9673 23489 9707
rect 23523 9704 23535 9707
rect 23566 9704 23572 9716
rect 23523 9676 23572 9704
rect 23523 9673 23535 9676
rect 23477 9667 23535 9673
rect 23566 9664 23572 9676
rect 23624 9664 23630 9716
rect 3896 9608 4200 9636
rect 3789 9599 3847 9605
rect 3804 9568 3832 9599
rect 3878 9568 3884 9580
rect 3804 9540 3884 9568
rect 3878 9528 3884 9540
rect 3936 9528 3942 9580
rect 4172 9577 4200 9608
rect 6546 9596 6552 9648
rect 6604 9636 6610 9648
rect 6733 9639 6791 9645
rect 6733 9636 6745 9639
rect 6604 9608 6745 9636
rect 6604 9596 6610 9608
rect 6733 9605 6745 9608
rect 6779 9636 6791 9639
rect 6779 9608 7328 9636
rect 6779 9605 6791 9608
rect 6733 9599 6791 9605
rect 4065 9571 4123 9577
rect 4065 9537 4077 9571
rect 4111 9537 4123 9571
rect 4065 9531 4123 9537
rect 4157 9571 4215 9577
rect 4157 9537 4169 9571
rect 4203 9537 4215 9571
rect 4157 9531 4215 9537
rect 4433 9571 4491 9577
rect 4433 9537 4445 9571
rect 4479 9568 4491 9571
rect 5169 9571 5227 9577
rect 4479 9540 4844 9568
rect 4479 9537 4491 9540
rect 4433 9531 4491 9537
rect 4080 9432 4108 9531
rect 4172 9500 4200 9531
rect 4614 9500 4620 9512
rect 4172 9472 4620 9500
rect 4614 9460 4620 9472
rect 4672 9460 4678 9512
rect 4706 9460 4712 9512
rect 4764 9460 4770 9512
rect 4816 9509 4844 9540
rect 5169 9537 5181 9571
rect 5215 9568 5227 9571
rect 5350 9568 5356 9580
rect 5215 9540 5356 9568
rect 5215 9537 5227 9540
rect 5169 9531 5227 9537
rect 5350 9528 5356 9540
rect 5408 9528 5414 9580
rect 5445 9571 5503 9577
rect 5445 9537 5457 9571
rect 5491 9568 5503 9571
rect 5534 9568 5540 9580
rect 5491 9540 5540 9568
rect 5491 9537 5503 9540
rect 5445 9531 5503 9537
rect 5534 9528 5540 9540
rect 5592 9528 5598 9580
rect 5626 9528 5632 9580
rect 5684 9577 5690 9580
rect 5684 9571 5697 9577
rect 5685 9537 5697 9571
rect 5684 9531 5697 9537
rect 6365 9571 6423 9577
rect 6365 9537 6377 9571
rect 6411 9568 6423 9571
rect 6638 9568 6644 9580
rect 6411 9540 6644 9568
rect 6411 9537 6423 9540
rect 6365 9531 6423 9537
rect 5684 9528 5690 9531
rect 6638 9528 6644 9540
rect 6696 9528 6702 9580
rect 6825 9571 6883 9577
rect 6825 9537 6837 9571
rect 6871 9568 6883 9571
rect 7190 9568 7196 9580
rect 6871 9540 7196 9568
rect 6871 9537 6883 9540
rect 6825 9531 6883 9537
rect 7190 9528 7196 9540
rect 7248 9528 7254 9580
rect 7300 9577 7328 9608
rect 7466 9596 7472 9648
rect 7524 9596 7530 9648
rect 7576 9608 8156 9636
rect 7285 9571 7343 9577
rect 7285 9537 7297 9571
rect 7331 9568 7343 9571
rect 7576 9568 7604 9608
rect 7331 9540 7604 9568
rect 7929 9571 7987 9577
rect 7331 9537 7343 9540
rect 7285 9531 7343 9537
rect 7929 9537 7941 9571
rect 7975 9537 7987 9571
rect 8128 9568 8156 9608
rect 8754 9596 8760 9648
rect 8812 9596 8818 9648
rect 11882 9596 11888 9648
rect 11940 9636 11946 9648
rect 19702 9636 19708 9648
rect 11940 9608 13032 9636
rect 11940 9596 11946 9608
rect 9309 9571 9367 9577
rect 9309 9568 9321 9571
rect 8128 9540 9321 9568
rect 7929 9531 7987 9537
rect 9309 9537 9321 9540
rect 9355 9568 9367 9571
rect 10318 9568 10324 9580
rect 9355 9540 10324 9568
rect 9355 9537 9367 9540
rect 9309 9531 9367 9537
rect 4801 9503 4859 9509
rect 4801 9469 4813 9503
rect 4847 9469 4859 9503
rect 4801 9463 4859 9469
rect 4982 9460 4988 9512
rect 5040 9460 5046 9512
rect 5077 9503 5135 9509
rect 5077 9469 5089 9503
rect 5123 9500 5135 9503
rect 5261 9503 5319 9509
rect 5123 9472 5212 9500
rect 5123 9469 5135 9472
rect 5077 9463 5135 9469
rect 5184 9432 5212 9472
rect 5261 9469 5273 9503
rect 5307 9500 5319 9503
rect 7745 9503 7803 9509
rect 5307 9472 5488 9500
rect 5307 9469 5319 9472
rect 5261 9463 5319 9469
rect 3620 9404 5212 9432
rect 5460 9432 5488 9472
rect 7745 9469 7757 9503
rect 7791 9469 7803 9503
rect 7745 9463 7803 9469
rect 5810 9432 5816 9444
rect 5460 9404 5816 9432
rect 3418 9324 3424 9376
rect 3476 9324 3482 9376
rect 3620 9373 3648 9404
rect 3605 9367 3663 9373
rect 3605 9333 3617 9367
rect 3651 9333 3663 9367
rect 3605 9327 3663 9333
rect 3786 9324 3792 9376
rect 3844 9364 3850 9376
rect 3881 9367 3939 9373
rect 3881 9364 3893 9367
rect 3844 9336 3893 9364
rect 3844 9324 3850 9336
rect 3881 9333 3893 9336
rect 3927 9333 3939 9367
rect 3881 9327 3939 9333
rect 4249 9367 4307 9373
rect 4249 9333 4261 9367
rect 4295 9364 4307 9367
rect 4706 9364 4712 9376
rect 4295 9336 4712 9364
rect 4295 9333 4307 9336
rect 4249 9327 4307 9333
rect 4706 9324 4712 9336
rect 4764 9324 4770 9376
rect 5184 9364 5212 9404
rect 5810 9392 5816 9404
rect 5868 9392 5874 9444
rect 7469 9435 7527 9441
rect 7469 9401 7481 9435
rect 7515 9432 7527 9435
rect 7760 9432 7788 9463
rect 7834 9460 7840 9512
rect 7892 9500 7898 9512
rect 7944 9500 7972 9531
rect 10318 9528 10324 9540
rect 10376 9528 10382 9580
rect 11698 9528 11704 9580
rect 11756 9528 11762 9580
rect 12802 9528 12808 9580
rect 12860 9528 12866 9580
rect 13004 9577 13032 9608
rect 19628 9608 19708 9636
rect 12989 9571 13047 9577
rect 12989 9537 13001 9571
rect 13035 9537 13047 9571
rect 12989 9531 13047 9537
rect 13906 9528 13912 9580
rect 13964 9568 13970 9580
rect 14829 9571 14887 9577
rect 14829 9568 14841 9571
rect 13964 9540 14841 9568
rect 13964 9528 13970 9540
rect 14829 9537 14841 9540
rect 14875 9537 14887 9571
rect 14829 9531 14887 9537
rect 15194 9528 15200 9580
rect 15252 9568 15258 9580
rect 15470 9568 15476 9580
rect 15252 9540 15476 9568
rect 15252 9528 15258 9540
rect 15470 9528 15476 9540
rect 15528 9528 15534 9580
rect 16482 9528 16488 9580
rect 16540 9568 16546 9580
rect 17037 9571 17095 9577
rect 17037 9568 17049 9571
rect 16540 9540 17049 9568
rect 16540 9528 16546 9540
rect 17037 9537 17049 9540
rect 17083 9537 17095 9571
rect 17037 9531 17095 9537
rect 17313 9571 17371 9577
rect 17313 9537 17325 9571
rect 17359 9568 17371 9571
rect 17402 9568 17408 9580
rect 17359 9540 17408 9568
rect 17359 9537 17371 9540
rect 17313 9531 17371 9537
rect 17402 9528 17408 9540
rect 17460 9528 17466 9580
rect 19518 9528 19524 9580
rect 19576 9528 19582 9580
rect 19628 9577 19656 9608
rect 19702 9596 19708 9608
rect 19760 9596 19766 9648
rect 24578 9636 24584 9648
rect 23676 9608 24584 9636
rect 19613 9571 19671 9577
rect 19613 9537 19625 9571
rect 19659 9537 19671 9571
rect 19613 9531 19671 9537
rect 19794 9528 19800 9580
rect 19852 9528 19858 9580
rect 23676 9577 23704 9608
rect 24578 9596 24584 9608
rect 24636 9596 24642 9648
rect 23661 9571 23719 9577
rect 23661 9537 23673 9571
rect 23707 9537 23719 9571
rect 23661 9531 23719 9537
rect 23750 9528 23756 9580
rect 23808 9528 23814 9580
rect 23842 9528 23848 9580
rect 23900 9568 23906 9580
rect 23937 9571 23995 9577
rect 23937 9568 23949 9571
rect 23900 9540 23949 9568
rect 23900 9528 23906 9540
rect 23937 9537 23949 9540
rect 23983 9537 23995 9571
rect 23937 9531 23995 9537
rect 24026 9528 24032 9580
rect 24084 9528 24090 9580
rect 7892 9472 7972 9500
rect 7892 9460 7898 9472
rect 8570 9460 8576 9512
rect 8628 9460 8634 9512
rect 9398 9460 9404 9512
rect 9456 9460 9462 9512
rect 11790 9460 11796 9512
rect 11848 9460 11854 9512
rect 14458 9460 14464 9512
rect 14516 9500 14522 9512
rect 15105 9503 15163 9509
rect 15105 9500 15117 9503
rect 14516 9472 15117 9500
rect 14516 9460 14522 9472
rect 15105 9469 15117 9472
rect 15151 9469 15163 9503
rect 15381 9503 15439 9509
rect 15381 9500 15393 9503
rect 15105 9463 15163 9469
rect 15212 9472 15393 9500
rect 9416 9432 9444 9460
rect 7515 9404 7788 9432
rect 7944 9404 9444 9432
rect 7515 9401 7527 9404
rect 7469 9395 7527 9401
rect 5534 9364 5540 9376
rect 5184 9336 5540 9364
rect 5534 9324 5540 9336
rect 5592 9324 5598 9376
rect 6546 9324 6552 9376
rect 6604 9324 6610 9376
rect 7190 9324 7196 9376
rect 7248 9364 7254 9376
rect 7944 9364 7972 9404
rect 12066 9392 12072 9444
rect 12124 9392 12130 9444
rect 13630 9392 13636 9444
rect 13688 9432 13694 9444
rect 14553 9435 14611 9441
rect 14553 9432 14565 9435
rect 13688 9404 14565 9432
rect 13688 9392 13694 9404
rect 14553 9401 14565 9404
rect 14599 9401 14611 9435
rect 14553 9395 14611 9401
rect 7248 9336 7972 9364
rect 7248 9324 7254 9336
rect 14182 9324 14188 9376
rect 14240 9364 14246 9376
rect 15212 9364 15240 9472
rect 15381 9469 15393 9472
rect 15427 9469 15439 9503
rect 15381 9463 15439 9469
rect 16022 9460 16028 9512
rect 16080 9500 16086 9512
rect 17129 9503 17187 9509
rect 17129 9500 17141 9503
rect 16080 9472 17141 9500
rect 16080 9460 16086 9472
rect 17129 9469 17141 9472
rect 17175 9469 17187 9503
rect 17129 9463 17187 9469
rect 19705 9503 19763 9509
rect 19705 9469 19717 9503
rect 19751 9500 19763 9503
rect 19886 9500 19892 9512
rect 19751 9472 19892 9500
rect 19751 9469 19763 9472
rect 19705 9463 19763 9469
rect 19886 9460 19892 9472
rect 19944 9460 19950 9512
rect 23768 9500 23796 9528
rect 25774 9500 25780 9512
rect 23768 9472 25780 9500
rect 25774 9460 25780 9472
rect 25832 9460 25838 9512
rect 17221 9435 17279 9441
rect 17221 9401 17233 9435
rect 17267 9432 17279 9435
rect 17310 9432 17316 9444
rect 17267 9404 17316 9432
rect 17267 9401 17279 9404
rect 17221 9395 17279 9401
rect 17310 9392 17316 9404
rect 17368 9392 17374 9444
rect 14240 9336 15240 9364
rect 14240 9324 14246 9336
rect 16850 9324 16856 9376
rect 16908 9324 16914 9376
rect 19518 9324 19524 9376
rect 19576 9364 19582 9376
rect 19981 9367 20039 9373
rect 19981 9364 19993 9367
rect 19576 9336 19993 9364
rect 19576 9324 19582 9336
rect 19981 9333 19993 9336
rect 20027 9333 20039 9367
rect 19981 9327 20039 9333
rect 1104 9274 27876 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 27876 9274
rect 1104 9200 27876 9222
rect 8113 9163 8171 9169
rect 8113 9129 8125 9163
rect 8159 9160 8171 9163
rect 8202 9160 8208 9172
rect 8159 9132 8208 9160
rect 8159 9129 8171 9132
rect 8113 9123 8171 9129
rect 8202 9120 8208 9132
rect 8260 9120 8266 9172
rect 12802 9120 12808 9172
rect 12860 9120 12866 9172
rect 16209 9163 16267 9169
rect 16209 9129 16221 9163
rect 16255 9160 16267 9163
rect 16390 9160 16396 9172
rect 16255 9132 16396 9160
rect 16255 9129 16267 9132
rect 16209 9123 16267 9129
rect 16390 9120 16396 9132
rect 16448 9120 16454 9172
rect 19705 9163 19763 9169
rect 19705 9129 19717 9163
rect 19751 9160 19763 9163
rect 20162 9160 20168 9172
rect 19751 9132 20168 9160
rect 19751 9129 19763 9132
rect 19705 9123 19763 9129
rect 20162 9120 20168 9132
rect 20220 9120 20226 9172
rect 21450 9120 21456 9172
rect 21508 9160 21514 9172
rect 21634 9160 21640 9172
rect 21508 9132 21640 9160
rect 21508 9120 21514 9132
rect 21634 9120 21640 9132
rect 21692 9160 21698 9172
rect 21821 9163 21879 9169
rect 21821 9160 21833 9163
rect 21692 9132 21833 9160
rect 21692 9120 21698 9132
rect 21821 9129 21833 9132
rect 21867 9129 21879 9163
rect 21821 9123 21879 9129
rect 4982 9052 4988 9104
rect 5040 9092 5046 9104
rect 5258 9092 5264 9104
rect 5040 9064 5264 9092
rect 5040 9052 5046 9064
rect 5258 9052 5264 9064
rect 5316 9092 5322 9104
rect 11333 9095 11391 9101
rect 5316 9064 5948 9092
rect 5316 9052 5322 9064
rect 3418 8984 3424 9036
rect 3476 9024 3482 9036
rect 5353 9027 5411 9033
rect 3476 8996 4016 9024
rect 3476 8984 3482 8996
rect 3786 8916 3792 8968
rect 3844 8916 3850 8968
rect 3988 8965 4016 8996
rect 5353 8993 5365 9027
rect 5399 9024 5411 9027
rect 5813 9027 5871 9033
rect 5813 9024 5825 9027
rect 5399 8996 5825 9024
rect 5399 8993 5411 8996
rect 5353 8987 5411 8993
rect 5813 8993 5825 8996
rect 5859 8993 5871 9027
rect 5813 8987 5871 8993
rect 3973 8959 4031 8965
rect 3973 8925 3985 8959
rect 4019 8925 4031 8959
rect 3973 8919 4031 8925
rect 5261 8959 5319 8965
rect 5261 8925 5273 8959
rect 5307 8956 5319 8959
rect 5442 8956 5448 8968
rect 5307 8928 5448 8956
rect 5307 8925 5319 8928
rect 5261 8919 5319 8925
rect 5442 8916 5448 8928
rect 5500 8916 5506 8968
rect 5534 8916 5540 8968
rect 5592 8956 5598 8968
rect 5920 8965 5948 9064
rect 11333 9061 11345 9095
rect 11379 9092 11391 9095
rect 11422 9092 11428 9104
rect 11379 9064 11428 9092
rect 11379 9061 11391 9064
rect 11333 9055 11391 9061
rect 11422 9052 11428 9064
rect 11480 9052 11486 9104
rect 19889 9095 19947 9101
rect 19889 9061 19901 9095
rect 19935 9061 19947 9095
rect 19889 9055 19947 9061
rect 21545 9095 21603 9101
rect 21545 9061 21557 9095
rect 21591 9092 21603 9095
rect 22094 9092 22100 9104
rect 21591 9064 22100 9092
rect 21591 9061 21603 9064
rect 21545 9055 21603 9061
rect 6546 8984 6552 9036
rect 6604 8984 6610 9036
rect 9766 8984 9772 9036
rect 9824 9024 9830 9036
rect 10045 9027 10103 9033
rect 9824 8996 9996 9024
rect 9824 8984 9830 8996
rect 5721 8959 5779 8965
rect 5721 8956 5733 8959
rect 5592 8928 5733 8956
rect 5592 8916 5598 8928
rect 5721 8925 5733 8928
rect 5767 8925 5779 8959
rect 5721 8919 5779 8925
rect 5905 8959 5963 8965
rect 5905 8925 5917 8959
rect 5951 8925 5963 8959
rect 5905 8919 5963 8925
rect 6730 8916 6736 8968
rect 6788 8916 6794 8968
rect 7834 8916 7840 8968
rect 7892 8956 7898 8968
rect 7929 8959 7987 8965
rect 7929 8956 7941 8959
rect 7892 8928 7941 8956
rect 7892 8916 7898 8928
rect 7929 8925 7941 8928
rect 7975 8925 7987 8959
rect 7929 8919 7987 8925
rect 8110 8916 8116 8968
rect 8168 8916 8174 8968
rect 9968 8942 9996 8996
rect 10045 8993 10057 9027
rect 10091 9024 10103 9027
rect 10134 9024 10140 9036
rect 10091 8996 10140 9024
rect 10091 8993 10103 8996
rect 10045 8987 10103 8993
rect 10134 8984 10140 8996
rect 10192 9024 10198 9036
rect 11238 9024 11244 9036
rect 10192 8996 11244 9024
rect 10192 8984 10198 8996
rect 11238 8984 11244 8996
rect 11296 8984 11302 9036
rect 13630 8984 13636 9036
rect 13688 8984 13694 9036
rect 13814 8984 13820 9036
rect 13872 9024 13878 9036
rect 15102 9024 15108 9036
rect 13872 8996 15108 9024
rect 13872 8984 13878 8996
rect 15102 8984 15108 8996
rect 15160 8984 15166 9036
rect 15289 9027 15347 9033
rect 15289 8993 15301 9027
rect 15335 9024 15347 9027
rect 15562 9024 15568 9036
rect 15335 8996 15568 9024
rect 15335 8993 15347 8996
rect 15289 8987 15347 8993
rect 15562 8984 15568 8996
rect 15620 8984 15626 9036
rect 16850 8984 16856 9036
rect 16908 8984 16914 9036
rect 17589 9027 17647 9033
rect 17589 8993 17601 9027
rect 17635 9024 17647 9027
rect 19904 9024 19932 9055
rect 22094 9052 22100 9064
rect 22152 9052 22158 9104
rect 22189 9095 22247 9101
rect 22189 9061 22201 9095
rect 22235 9061 22247 9095
rect 22189 9055 22247 9061
rect 20165 9027 20223 9033
rect 20165 9024 20177 9027
rect 17635 8996 19840 9024
rect 19904 8996 20177 9024
rect 17635 8993 17647 8996
rect 17589 8987 17647 8993
rect 11054 8916 11060 8968
rect 11112 8916 11118 8968
rect 11146 8916 11152 8968
rect 11204 8956 11210 8968
rect 11333 8959 11391 8965
rect 11333 8956 11345 8959
rect 11204 8928 11345 8956
rect 11204 8916 11210 8928
rect 11333 8925 11345 8928
rect 11379 8956 11391 8959
rect 11606 8956 11612 8968
rect 11379 8928 11612 8956
rect 11379 8925 11391 8928
rect 11333 8919 11391 8925
rect 11606 8916 11612 8928
rect 11664 8916 11670 8968
rect 12342 8916 12348 8968
rect 12400 8916 12406 8968
rect 12618 8916 12624 8968
rect 12676 8916 12682 8968
rect 13541 8959 13599 8965
rect 13541 8925 13553 8959
rect 13587 8956 13599 8959
rect 13832 8956 13860 8984
rect 13587 8928 13860 8956
rect 13909 8959 13967 8965
rect 13587 8925 13599 8928
rect 13541 8919 13599 8925
rect 13909 8925 13921 8959
rect 13955 8956 13967 8959
rect 14090 8956 14096 8968
rect 13955 8928 14096 8956
rect 13955 8925 13967 8928
rect 13909 8919 13967 8925
rect 14090 8916 14096 8928
rect 14148 8916 14154 8968
rect 14274 8916 14280 8968
rect 14332 8916 14338 8968
rect 14458 8916 14464 8968
rect 14516 8916 14522 8968
rect 16761 8959 16819 8965
rect 16761 8956 16773 8959
rect 16040 8928 16773 8956
rect 10873 8891 10931 8897
rect 10873 8857 10885 8891
rect 10919 8888 10931 8891
rect 11238 8888 11244 8900
rect 10919 8860 11244 8888
rect 10919 8857 10931 8860
rect 10873 8851 10931 8857
rect 11238 8848 11244 8860
rect 11296 8848 11302 8900
rect 16040 8897 16068 8928
rect 16761 8925 16773 8928
rect 16807 8956 16819 8959
rect 17034 8956 17040 8968
rect 16807 8928 17040 8956
rect 16807 8925 16819 8928
rect 16761 8919 16819 8925
rect 17034 8916 17040 8928
rect 17092 8916 17098 8968
rect 17678 8916 17684 8968
rect 17736 8916 17742 8968
rect 17862 8916 17868 8968
rect 17920 8916 17926 8968
rect 17957 8959 18015 8965
rect 17957 8925 17969 8959
rect 18003 8925 18015 8959
rect 17957 8919 18015 8925
rect 13817 8891 13875 8897
rect 13817 8857 13829 8891
rect 13863 8888 13875 8891
rect 16025 8891 16083 8897
rect 16025 8888 16037 8891
rect 13863 8860 16037 8888
rect 13863 8857 13875 8860
rect 13817 8851 13875 8857
rect 16025 8857 16037 8860
rect 16071 8857 16083 8891
rect 16025 8851 16083 8857
rect 16206 8848 16212 8900
rect 16264 8897 16270 8900
rect 16264 8891 16283 8897
rect 16271 8857 16283 8891
rect 17972 8888 18000 8919
rect 18138 8916 18144 8968
rect 18196 8916 18202 8968
rect 19812 8956 19840 8996
rect 20165 8993 20177 8996
rect 20211 8993 20223 9027
rect 22204 9024 22232 9055
rect 24578 9052 24584 9104
rect 24636 9092 24642 9104
rect 25590 9092 25596 9104
rect 24636 9064 25596 9092
rect 24636 9052 24642 9064
rect 25590 9052 25596 9064
rect 25648 9092 25654 9104
rect 25648 9064 25912 9092
rect 25648 9052 25654 9064
rect 22278 9024 22284 9036
rect 20165 8987 20223 8993
rect 21560 8996 21864 9024
rect 22204 8996 22284 9024
rect 20254 8956 20260 8968
rect 19812 8928 20260 8956
rect 20254 8916 20260 8928
rect 20312 8916 20318 8968
rect 21358 8916 21364 8968
rect 21416 8956 21422 8968
rect 21560 8965 21588 8996
rect 21545 8959 21603 8965
rect 21545 8956 21557 8959
rect 21416 8928 21557 8956
rect 21416 8916 21422 8928
rect 21545 8925 21557 8928
rect 21591 8925 21603 8959
rect 21545 8919 21603 8925
rect 21634 8916 21640 8968
rect 21692 8956 21698 8968
rect 21836 8965 21864 8996
rect 22278 8984 22284 8996
rect 22336 9024 22342 9036
rect 22336 8996 22876 9024
rect 22336 8984 22342 8996
rect 21729 8959 21787 8965
rect 21729 8956 21741 8959
rect 21692 8928 21741 8956
rect 21692 8916 21698 8928
rect 21729 8925 21741 8928
rect 21775 8925 21787 8959
rect 21729 8919 21787 8925
rect 21821 8959 21879 8965
rect 21821 8925 21833 8959
rect 21867 8956 21879 8959
rect 21910 8956 21916 8968
rect 21867 8928 21916 8956
rect 21867 8925 21879 8928
rect 21821 8919 21879 8925
rect 21910 8916 21916 8928
rect 21968 8916 21974 8968
rect 22002 8916 22008 8968
rect 22060 8916 22066 8968
rect 22186 8956 22192 8968
rect 22112 8928 22192 8956
rect 16264 8851 16283 8857
rect 16408 8860 18000 8888
rect 16264 8848 16270 8851
rect 4157 8823 4215 8829
rect 4157 8789 4169 8823
rect 4203 8820 4215 8823
rect 4798 8820 4804 8832
rect 4203 8792 4804 8820
rect 4203 8789 4215 8792
rect 4157 8783 4215 8789
rect 4798 8780 4804 8792
rect 4856 8780 4862 8832
rect 5629 8823 5687 8829
rect 5629 8789 5641 8823
rect 5675 8820 5687 8823
rect 5902 8820 5908 8832
rect 5675 8792 5908 8820
rect 5675 8789 5687 8792
rect 5629 8783 5687 8789
rect 5902 8780 5908 8792
rect 5960 8780 5966 8832
rect 7466 8780 7472 8832
rect 7524 8780 7530 8832
rect 7742 8780 7748 8832
rect 7800 8780 7806 8832
rect 11054 8780 11060 8832
rect 11112 8820 11118 8832
rect 16408 8829 16436 8860
rect 17880 8832 17908 8860
rect 19518 8848 19524 8900
rect 19576 8848 19582 8900
rect 21085 8891 21143 8897
rect 21085 8857 21097 8891
rect 21131 8888 21143 8891
rect 22112 8888 22140 8928
rect 22186 8916 22192 8928
rect 22244 8916 22250 8968
rect 22370 8916 22376 8968
rect 22428 8916 22434 8968
rect 22848 8965 22876 8996
rect 23842 8984 23848 9036
rect 23900 9024 23906 9036
rect 24765 9027 24823 9033
rect 24765 9024 24777 9027
rect 23900 8996 24777 9024
rect 23900 8984 23906 8996
rect 24765 8993 24777 8996
rect 24811 8993 24823 9027
rect 24765 8987 24823 8993
rect 24872 8996 25544 9024
rect 22833 8959 22891 8965
rect 22833 8925 22845 8959
rect 22879 8956 22891 8959
rect 23290 8956 23296 8968
rect 22879 8928 23296 8956
rect 22879 8925 22891 8928
rect 22833 8919 22891 8925
rect 23290 8916 23296 8928
rect 23348 8916 23354 8968
rect 24029 8959 24087 8965
rect 24029 8925 24041 8959
rect 24075 8925 24087 8959
rect 24029 8919 24087 8925
rect 24044 8888 24072 8919
rect 24210 8916 24216 8968
rect 24268 8916 24274 8968
rect 24394 8916 24400 8968
rect 24452 8916 24458 8968
rect 24670 8916 24676 8968
rect 24728 8956 24734 8968
rect 24872 8956 24900 8996
rect 25516 8965 25544 8996
rect 24728 8928 24900 8956
rect 24949 8959 25007 8965
rect 24728 8916 24734 8928
rect 24949 8925 24961 8959
rect 24995 8925 25007 8959
rect 25133 8959 25191 8965
rect 25133 8956 25145 8959
rect 24949 8919 25007 8925
rect 25056 8928 25145 8956
rect 24964 8888 24992 8919
rect 21131 8860 22140 8888
rect 22204 8860 24072 8888
rect 24136 8860 24992 8888
rect 25056 8888 25084 8928
rect 25133 8925 25145 8928
rect 25179 8925 25191 8959
rect 25133 8919 25191 8925
rect 25501 8959 25559 8965
rect 25501 8925 25513 8959
rect 25547 8925 25559 8959
rect 25501 8919 25559 8925
rect 25685 8959 25743 8965
rect 25685 8925 25697 8959
rect 25731 8956 25743 8959
rect 25774 8956 25780 8968
rect 25731 8928 25780 8956
rect 25731 8925 25743 8928
rect 25685 8919 25743 8925
rect 25774 8916 25780 8928
rect 25832 8916 25838 8968
rect 25884 8965 25912 9064
rect 25869 8959 25927 8965
rect 25869 8925 25881 8959
rect 25915 8925 25927 8959
rect 25869 8919 25927 8925
rect 25593 8891 25651 8897
rect 25593 8888 25605 8891
rect 25056 8860 25605 8888
rect 21131 8857 21143 8860
rect 21085 8851 21143 8857
rect 22204 8832 22232 8860
rect 24136 8832 24164 8860
rect 11149 8823 11207 8829
rect 11149 8820 11161 8823
rect 11112 8792 11161 8820
rect 11112 8780 11118 8792
rect 11149 8789 11161 8792
rect 11195 8820 11207 8823
rect 12437 8823 12495 8829
rect 12437 8820 12449 8823
rect 11195 8792 12449 8820
rect 11195 8789 11207 8792
rect 11149 8783 11207 8789
rect 12437 8789 12449 8792
rect 12483 8789 12495 8823
rect 12437 8783 12495 8789
rect 16393 8823 16451 8829
rect 16393 8789 16405 8823
rect 16439 8789 16451 8823
rect 16393 8783 16451 8789
rect 17402 8780 17408 8832
rect 17460 8820 17466 8832
rect 17681 8823 17739 8829
rect 17681 8820 17693 8823
rect 17460 8792 17693 8820
rect 17460 8780 17466 8792
rect 17681 8789 17693 8792
rect 17727 8789 17739 8823
rect 17681 8783 17739 8789
rect 17862 8780 17868 8832
rect 17920 8780 17926 8832
rect 18046 8780 18052 8832
rect 18104 8780 18110 8832
rect 19702 8780 19708 8832
rect 19760 8829 19766 8832
rect 19760 8823 19779 8829
rect 19767 8820 19779 8823
rect 20346 8820 20352 8832
rect 19767 8792 20352 8820
rect 19767 8789 19779 8792
rect 19760 8783 19779 8789
rect 19760 8780 19766 8783
rect 20346 8780 20352 8792
rect 20404 8780 20410 8832
rect 20438 8780 20444 8832
rect 20496 8820 20502 8832
rect 22186 8820 22192 8832
rect 20496 8792 22192 8820
rect 20496 8780 20502 8792
rect 22186 8780 22192 8792
rect 22244 8780 22250 8832
rect 22646 8780 22652 8832
rect 22704 8780 22710 8832
rect 22738 8780 22744 8832
rect 22796 8780 22802 8832
rect 24118 8780 24124 8832
rect 24176 8780 24182 8832
rect 24486 8780 24492 8832
rect 24544 8820 24550 8832
rect 25056 8820 25084 8860
rect 25593 8857 25605 8860
rect 25639 8857 25651 8891
rect 25593 8851 25651 8857
rect 24544 8792 25084 8820
rect 24544 8780 24550 8792
rect 25130 8780 25136 8832
rect 25188 8820 25194 8832
rect 25317 8823 25375 8829
rect 25317 8820 25329 8823
rect 25188 8792 25329 8820
rect 25188 8780 25194 8792
rect 25317 8789 25329 8792
rect 25363 8789 25375 8823
rect 25317 8783 25375 8789
rect 1104 8730 27876 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 27876 8730
rect 1104 8656 27876 8678
rect 4709 8619 4767 8625
rect 4709 8585 4721 8619
rect 4755 8616 4767 8619
rect 4890 8616 4896 8628
rect 4755 8588 4896 8616
rect 4755 8585 4767 8588
rect 4709 8579 4767 8585
rect 4890 8576 4896 8588
rect 4948 8576 4954 8628
rect 10134 8576 10140 8628
rect 10192 8576 10198 8628
rect 15470 8616 15476 8628
rect 14936 8588 15476 8616
rect 6733 8551 6791 8557
rect 6733 8517 6745 8551
rect 6779 8548 6791 8551
rect 6822 8548 6828 8560
rect 6779 8520 6828 8548
rect 6779 8517 6791 8520
rect 6733 8511 6791 8517
rect 6822 8508 6828 8520
rect 6880 8548 6886 8560
rect 6880 8520 12112 8548
rect 6880 8508 6886 8520
rect 3510 8440 3516 8492
rect 3568 8440 3574 8492
rect 4614 8440 4620 8492
rect 4672 8440 4678 8492
rect 4706 8440 4712 8492
rect 4764 8440 4770 8492
rect 4893 8483 4951 8489
rect 4893 8449 4905 8483
rect 4939 8480 4951 8483
rect 5074 8480 5080 8492
rect 4939 8452 5080 8480
rect 4939 8449 4951 8452
rect 4893 8443 4951 8449
rect 5074 8440 5080 8452
rect 5132 8480 5138 8492
rect 6549 8483 6607 8489
rect 6549 8480 6561 8483
rect 5132 8452 6561 8480
rect 5132 8440 5138 8452
rect 6549 8449 6561 8452
rect 6595 8480 6607 8483
rect 9493 8483 9551 8489
rect 6595 8452 6868 8480
rect 6595 8449 6607 8452
rect 6549 8443 6607 8449
rect 3418 8372 3424 8424
rect 3476 8372 3482 8424
rect 4724 8412 4752 8440
rect 4982 8412 4988 8424
rect 4724 8384 4988 8412
rect 4982 8372 4988 8384
rect 5040 8372 5046 8424
rect 6365 8415 6423 8421
rect 6365 8381 6377 8415
rect 6411 8412 6423 8415
rect 6730 8412 6736 8424
rect 6411 8384 6736 8412
rect 6411 8381 6423 8384
rect 6365 8375 6423 8381
rect 6730 8372 6736 8384
rect 6788 8372 6794 8424
rect 3881 8347 3939 8353
rect 3881 8313 3893 8347
rect 3927 8344 3939 8347
rect 4706 8344 4712 8356
rect 3927 8316 4712 8344
rect 3927 8313 3939 8316
rect 3881 8307 3939 8313
rect 4706 8304 4712 8316
rect 4764 8304 4770 8356
rect 4893 8279 4951 8285
rect 4893 8245 4905 8279
rect 4939 8276 4951 8279
rect 5258 8276 5264 8288
rect 4939 8248 5264 8276
rect 4939 8245 4951 8248
rect 4893 8239 4951 8245
rect 5258 8236 5264 8248
rect 5316 8236 5322 8288
rect 6840 8276 6868 8452
rect 9493 8449 9505 8483
rect 9539 8480 9551 8483
rect 10134 8480 10140 8492
rect 9539 8452 10140 8480
rect 9539 8449 9551 8452
rect 9493 8443 9551 8449
rect 10134 8440 10140 8452
rect 10192 8440 10198 8492
rect 11057 8483 11115 8489
rect 11057 8449 11069 8483
rect 11103 8480 11115 8483
rect 11146 8480 11152 8492
rect 11103 8452 11152 8480
rect 11103 8449 11115 8452
rect 11057 8443 11115 8449
rect 11146 8440 11152 8452
rect 11204 8440 11210 8492
rect 11238 8440 11244 8492
rect 11296 8440 11302 8492
rect 12084 8489 12112 8520
rect 12069 8483 12127 8489
rect 12069 8449 12081 8483
rect 12115 8449 12127 8483
rect 12069 8443 12127 8449
rect 12618 8440 12624 8492
rect 12676 8440 12682 8492
rect 14001 8483 14059 8489
rect 14001 8449 14013 8483
rect 14047 8449 14059 8483
rect 14001 8443 14059 8449
rect 9585 8415 9643 8421
rect 9585 8381 9597 8415
rect 9631 8412 9643 8415
rect 9766 8412 9772 8424
rect 9631 8384 9772 8412
rect 9631 8381 9643 8384
rect 9585 8375 9643 8381
rect 9766 8372 9772 8384
rect 9824 8372 9830 8424
rect 9858 8372 9864 8424
rect 9916 8412 9922 8424
rect 10505 8415 10563 8421
rect 10505 8412 10517 8415
rect 9916 8384 10517 8412
rect 9916 8372 9922 8384
rect 10505 8381 10517 8384
rect 10551 8381 10563 8415
rect 10505 8375 10563 8381
rect 13909 8415 13967 8421
rect 13909 8381 13921 8415
rect 13955 8412 13967 8415
rect 14016 8412 14044 8443
rect 14182 8440 14188 8492
rect 14240 8440 14246 8492
rect 14936 8489 14964 8588
rect 15470 8576 15476 8588
rect 15528 8576 15534 8628
rect 20254 8576 20260 8628
rect 20312 8576 20318 8628
rect 21634 8576 21640 8628
rect 21692 8616 21698 8628
rect 21692 8588 22140 8616
rect 21692 8576 21698 8588
rect 15933 8551 15991 8557
rect 15933 8517 15945 8551
rect 15979 8548 15991 8551
rect 16022 8548 16028 8560
rect 15979 8520 16028 8548
rect 15979 8517 15991 8520
rect 15933 8511 15991 8517
rect 16022 8508 16028 8520
rect 16080 8508 16086 8560
rect 18138 8548 18144 8560
rect 17144 8520 18144 8548
rect 15016 8492 15068 8498
rect 14921 8483 14979 8489
rect 14921 8449 14933 8483
rect 14967 8449 14979 8483
rect 14921 8443 14979 8449
rect 14936 8412 14964 8443
rect 16390 8440 16396 8492
rect 16448 8480 16454 8492
rect 16945 8483 17003 8489
rect 16945 8480 16957 8483
rect 16448 8452 16957 8480
rect 16448 8440 16454 8452
rect 16945 8449 16957 8452
rect 16991 8449 17003 8483
rect 16945 8443 17003 8449
rect 17034 8440 17040 8492
rect 17092 8440 17098 8492
rect 15016 8434 15068 8440
rect 17144 8424 17172 8520
rect 18138 8508 18144 8520
rect 18196 8548 18202 8560
rect 20272 8548 20300 8576
rect 21545 8551 21603 8557
rect 18196 8520 18644 8548
rect 20272 8520 21496 8548
rect 18196 8508 18202 8520
rect 17497 8483 17555 8489
rect 17497 8449 17509 8483
rect 17543 8480 17555 8483
rect 17586 8480 17592 8492
rect 17543 8452 17592 8480
rect 17543 8449 17555 8452
rect 17497 8443 17555 8449
rect 17586 8440 17592 8452
rect 17644 8440 17650 8492
rect 18616 8489 18644 8520
rect 17681 8483 17739 8489
rect 17681 8449 17693 8483
rect 17727 8449 17739 8483
rect 17681 8443 17739 8449
rect 17957 8483 18015 8489
rect 17957 8449 17969 8483
rect 18003 8480 18015 8483
rect 18233 8483 18291 8489
rect 18233 8480 18245 8483
rect 18003 8452 18245 8480
rect 18003 8449 18015 8452
rect 17957 8443 18015 8449
rect 18233 8449 18245 8452
rect 18279 8449 18291 8483
rect 18233 8443 18291 8449
rect 18601 8483 18659 8489
rect 18601 8449 18613 8483
rect 18647 8449 18659 8483
rect 18601 8443 18659 8449
rect 13955 8384 14964 8412
rect 13955 8381 13967 8384
rect 13909 8375 13967 8381
rect 16206 8372 16212 8424
rect 16264 8412 16270 8424
rect 16853 8415 16911 8421
rect 16853 8412 16865 8415
rect 16264 8384 16865 8412
rect 16264 8372 16270 8384
rect 16853 8381 16865 8384
rect 16899 8381 16911 8415
rect 16853 8375 16911 8381
rect 17126 8372 17132 8424
rect 17184 8372 17190 8424
rect 17696 8412 17724 8443
rect 19518 8440 19524 8492
rect 19576 8480 19582 8492
rect 20165 8483 20223 8489
rect 20165 8480 20177 8483
rect 19576 8452 20177 8480
rect 19576 8440 19582 8452
rect 20165 8449 20177 8452
rect 20211 8449 20223 8483
rect 20165 8443 20223 8449
rect 17512 8384 17724 8412
rect 17512 8356 17540 8384
rect 17862 8372 17868 8424
rect 17920 8412 17926 8424
rect 18049 8415 18107 8421
rect 18049 8412 18061 8415
rect 17920 8384 18061 8412
rect 17920 8372 17926 8384
rect 18049 8381 18061 8384
rect 18095 8381 18107 8415
rect 20180 8412 20208 8443
rect 20346 8440 20352 8492
rect 20404 8480 20410 8492
rect 20441 8483 20499 8489
rect 20441 8480 20453 8483
rect 20404 8452 20453 8480
rect 20404 8440 20410 8452
rect 20441 8449 20453 8452
rect 20487 8449 20499 8483
rect 20441 8443 20499 8449
rect 20530 8440 20536 8492
rect 20588 8480 20594 8492
rect 20824 8489 20852 8520
rect 20717 8483 20775 8489
rect 20717 8480 20729 8483
rect 20588 8452 20729 8480
rect 20588 8440 20594 8452
rect 20717 8449 20729 8452
rect 20763 8449 20775 8483
rect 20717 8443 20775 8449
rect 20809 8483 20867 8489
rect 20809 8449 20821 8483
rect 20855 8449 20867 8483
rect 20809 8443 20867 8449
rect 20993 8483 21051 8489
rect 20993 8449 21005 8483
rect 21039 8480 21051 8483
rect 21361 8483 21419 8489
rect 21361 8480 21373 8483
rect 21039 8452 21373 8480
rect 21039 8449 21051 8452
rect 20993 8443 21051 8449
rect 21361 8449 21373 8452
rect 21407 8449 21419 8483
rect 21361 8443 21419 8449
rect 21008 8412 21036 8443
rect 20180 8384 21036 8412
rect 21177 8415 21235 8421
rect 18049 8375 18107 8381
rect 21177 8381 21189 8415
rect 21223 8412 21235 8415
rect 21468 8412 21496 8520
rect 21545 8517 21557 8551
rect 21591 8548 21603 8551
rect 21591 8520 22048 8548
rect 21591 8517 21603 8520
rect 21545 8511 21603 8517
rect 22020 8492 22048 8520
rect 21821 8483 21879 8489
rect 21821 8449 21833 8483
rect 21867 8449 21879 8483
rect 21821 8443 21879 8449
rect 21223 8384 21496 8412
rect 21836 8412 21864 8443
rect 22002 8440 22008 8492
rect 22060 8440 22066 8492
rect 22112 8489 22140 8588
rect 22370 8576 22376 8628
rect 22428 8616 22434 8628
rect 22557 8619 22615 8625
rect 22557 8616 22569 8619
rect 22428 8588 22569 8616
rect 22428 8576 22434 8588
rect 22557 8585 22569 8588
rect 22603 8585 22615 8619
rect 22557 8579 22615 8585
rect 24216 8560 24268 8566
rect 24670 8548 24676 8560
rect 24268 8520 24676 8548
rect 24670 8508 24676 8520
rect 24728 8508 24734 8560
rect 24216 8502 24268 8508
rect 22097 8483 22155 8489
rect 22097 8449 22109 8483
rect 22143 8449 22155 8483
rect 22097 8443 22155 8449
rect 22186 8440 22192 8492
rect 22244 8480 22250 8492
rect 22281 8483 22339 8489
rect 22281 8480 22293 8483
rect 22244 8452 22293 8480
rect 22244 8440 22250 8452
rect 22281 8449 22293 8452
rect 22327 8449 22339 8483
rect 22281 8443 22339 8449
rect 22738 8440 22744 8492
rect 22796 8440 22802 8492
rect 23290 8440 23296 8492
rect 23348 8440 23354 8492
rect 24394 8440 24400 8492
rect 24452 8480 24458 8492
rect 25041 8483 25099 8489
rect 25041 8480 25053 8483
rect 24452 8452 25053 8480
rect 24452 8440 24458 8452
rect 25041 8449 25053 8452
rect 25087 8449 25099 8483
rect 25041 8443 25099 8449
rect 22756 8412 22784 8440
rect 21836 8384 22784 8412
rect 21223 8381 21235 8384
rect 21177 8375 21235 8381
rect 9214 8304 9220 8356
rect 9272 8344 9278 8356
rect 9953 8347 10011 8353
rect 9953 8344 9965 8347
rect 9272 8316 9965 8344
rect 9272 8304 9278 8316
rect 9953 8313 9965 8316
rect 9999 8313 10011 8347
rect 9953 8307 10011 8313
rect 16298 8304 16304 8356
rect 16356 8344 16362 8356
rect 16669 8347 16727 8353
rect 16669 8344 16681 8347
rect 16356 8316 16681 8344
rect 16356 8304 16362 8316
rect 16669 8313 16681 8316
rect 16715 8313 16727 8347
rect 16669 8307 16727 8313
rect 17494 8304 17500 8356
rect 17552 8304 17558 8356
rect 20625 8347 20683 8353
rect 20625 8313 20637 8347
rect 20671 8344 20683 8347
rect 20714 8344 20720 8356
rect 20671 8316 20720 8344
rect 20671 8313 20683 8316
rect 20625 8307 20683 8313
rect 20714 8304 20720 8316
rect 20772 8304 20778 8356
rect 21836 8344 21864 8384
rect 25130 8372 25136 8424
rect 25188 8372 25194 8424
rect 20824 8316 21864 8344
rect 8294 8276 8300 8288
rect 6840 8248 8300 8276
rect 8294 8236 8300 8248
rect 8352 8236 8358 8288
rect 9766 8236 9772 8288
rect 9824 8236 9830 8288
rect 10042 8236 10048 8288
rect 10100 8276 10106 8288
rect 10137 8279 10195 8285
rect 10137 8276 10149 8279
rect 10100 8248 10149 8276
rect 10100 8236 10106 8248
rect 10137 8245 10149 8248
rect 10183 8245 10195 8279
rect 10137 8239 10195 8245
rect 11057 8279 11115 8285
rect 11057 8245 11069 8279
rect 11103 8276 11115 8279
rect 11238 8276 11244 8288
rect 11103 8248 11244 8276
rect 11103 8245 11115 8248
rect 11057 8239 11115 8245
rect 11238 8236 11244 8248
rect 11296 8236 11302 8288
rect 13998 8236 14004 8288
rect 14056 8236 14062 8288
rect 19794 8236 19800 8288
rect 19852 8276 19858 8288
rect 20073 8279 20131 8285
rect 20073 8276 20085 8279
rect 19852 8248 20085 8276
rect 19852 8236 19858 8248
rect 20073 8245 20085 8248
rect 20119 8276 20131 8279
rect 20824 8276 20852 8316
rect 21910 8304 21916 8356
rect 21968 8344 21974 8356
rect 22189 8347 22247 8353
rect 22189 8344 22201 8347
rect 21968 8316 22201 8344
rect 21968 8304 21974 8316
rect 22189 8313 22201 8316
rect 22235 8313 22247 8347
rect 22189 8307 22247 8313
rect 23382 8304 23388 8356
rect 23440 8344 23446 8356
rect 24673 8347 24731 8353
rect 24673 8344 24685 8347
rect 23440 8316 24685 8344
rect 23440 8304 23446 8316
rect 24673 8313 24685 8316
rect 24719 8313 24731 8347
rect 24673 8307 24731 8313
rect 20119 8248 20852 8276
rect 20119 8245 20131 8248
rect 20073 8239 20131 8245
rect 1104 8186 27876 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 27876 8186
rect 1104 8112 27876 8134
rect 4985 8075 5043 8081
rect 4985 8041 4997 8075
rect 5031 8072 5043 8075
rect 5031 8044 6040 8072
rect 5031 8041 5043 8044
rect 4985 8035 5043 8041
rect 4706 8004 4712 8016
rect 4356 7976 4712 8004
rect 4356 7945 4384 7976
rect 4706 7964 4712 7976
rect 4764 8004 4770 8016
rect 4764 7976 5120 8004
rect 4764 7964 4770 7976
rect 4341 7939 4399 7945
rect 4341 7905 4353 7939
rect 4387 7905 4399 7939
rect 4341 7899 4399 7905
rect 4614 7896 4620 7948
rect 4672 7936 4678 7948
rect 5092 7945 5120 7976
rect 5442 7964 5448 8016
rect 5500 7964 5506 8016
rect 6012 8004 6040 8044
rect 7834 8032 7840 8084
rect 7892 8072 7898 8084
rect 8938 8072 8944 8084
rect 7892 8044 8944 8072
rect 7892 8032 7898 8044
rect 8938 8032 8944 8044
rect 8996 8072 9002 8084
rect 11146 8072 11152 8084
rect 8996 8044 11152 8072
rect 8996 8032 9002 8044
rect 11146 8032 11152 8044
rect 11204 8032 11210 8084
rect 12713 8075 12771 8081
rect 12713 8041 12725 8075
rect 12759 8072 12771 8075
rect 12894 8072 12900 8084
rect 12759 8044 12900 8072
rect 12759 8041 12771 8044
rect 12713 8035 12771 8041
rect 12894 8032 12900 8044
rect 12952 8032 12958 8084
rect 13170 8032 13176 8084
rect 13228 8072 13234 8084
rect 14182 8072 14188 8084
rect 13228 8044 14188 8072
rect 13228 8032 13234 8044
rect 14182 8032 14188 8044
rect 14240 8032 14246 8084
rect 15197 8075 15255 8081
rect 15197 8041 15209 8075
rect 15243 8072 15255 8075
rect 17126 8072 17132 8084
rect 15243 8044 17132 8072
rect 15243 8041 15255 8044
rect 15197 8035 15255 8041
rect 17126 8032 17132 8044
rect 17184 8032 17190 8084
rect 19429 8075 19487 8081
rect 19429 8041 19441 8075
rect 19475 8072 19487 8075
rect 20346 8072 20352 8084
rect 19475 8044 20352 8072
rect 19475 8041 19487 8044
rect 19429 8035 19487 8041
rect 20346 8032 20352 8044
rect 20404 8072 20410 8084
rect 21266 8072 21272 8084
rect 20404 8044 21272 8072
rect 20404 8032 20410 8044
rect 21266 8032 21272 8044
rect 21324 8032 21330 8084
rect 22741 8075 22799 8081
rect 22741 8041 22753 8075
rect 22787 8072 22799 8075
rect 24029 8075 24087 8081
rect 24029 8072 24041 8075
rect 22787 8044 24041 8072
rect 22787 8041 22799 8044
rect 22741 8035 22799 8041
rect 24029 8041 24041 8044
rect 24075 8072 24087 8075
rect 24394 8072 24400 8084
rect 24075 8044 24400 8072
rect 24075 8041 24087 8044
rect 24029 8035 24087 8041
rect 24394 8032 24400 8044
rect 24452 8032 24458 8084
rect 12434 8004 12440 8016
rect 6012 7976 12440 8004
rect 4801 7939 4859 7945
rect 4801 7936 4813 7939
rect 4672 7908 4813 7936
rect 4672 7896 4678 7908
rect 4801 7905 4813 7908
rect 4847 7905 4859 7939
rect 4801 7899 4859 7905
rect 5077 7939 5135 7945
rect 5077 7905 5089 7939
rect 5123 7905 5135 7939
rect 5077 7899 5135 7905
rect 4709 7871 4767 7877
rect 4709 7837 4721 7871
rect 4755 7837 4767 7871
rect 4709 7831 4767 7837
rect 4724 7800 4752 7831
rect 5258 7828 5264 7880
rect 5316 7828 5322 7880
rect 6012 7877 6040 7976
rect 12434 7964 12440 7976
rect 12492 7964 12498 8016
rect 13725 8007 13783 8013
rect 13725 7973 13737 8007
rect 13771 8004 13783 8007
rect 14274 8004 14280 8016
rect 13771 7976 14280 8004
rect 13771 7973 13783 7976
rect 13725 7967 13783 7973
rect 14274 7964 14280 7976
rect 14332 7964 14338 8016
rect 9214 7936 9220 7948
rect 7760 7908 9220 7936
rect 5997 7871 6055 7877
rect 5997 7837 6009 7871
rect 6043 7837 6055 7871
rect 5997 7831 6055 7837
rect 7650 7828 7656 7880
rect 7708 7828 7714 7880
rect 7760 7877 7788 7908
rect 7745 7871 7803 7877
rect 7745 7837 7757 7871
rect 7791 7837 7803 7871
rect 7745 7831 7803 7837
rect 7834 7828 7840 7880
rect 7892 7828 7898 7880
rect 8110 7828 8116 7880
rect 8168 7868 8174 7880
rect 8389 7871 8447 7877
rect 8389 7868 8401 7871
rect 8168 7840 8401 7868
rect 8168 7828 8174 7840
rect 8389 7837 8401 7840
rect 8435 7837 8447 7871
rect 8389 7831 8447 7837
rect 8478 7828 8484 7880
rect 8536 7828 8542 7880
rect 8570 7828 8576 7880
rect 8628 7828 8634 7880
rect 8938 7828 8944 7880
rect 8996 7828 9002 7880
rect 9140 7877 9168 7908
rect 9214 7896 9220 7908
rect 9272 7896 9278 7948
rect 11422 7896 11428 7948
rect 11480 7896 11486 7948
rect 13081 7939 13139 7945
rect 13081 7936 13093 7939
rect 12728 7908 13093 7936
rect 9125 7871 9183 7877
rect 9125 7837 9137 7871
rect 9171 7837 9183 7871
rect 9125 7831 9183 7837
rect 9766 7828 9772 7880
rect 9824 7828 9830 7880
rect 9858 7828 9864 7880
rect 9916 7828 9922 7880
rect 9953 7871 10011 7877
rect 9953 7837 9965 7871
rect 9999 7837 10011 7871
rect 9953 7831 10011 7837
rect 4890 7800 4896 7812
rect 4724 7772 4896 7800
rect 4890 7760 4896 7772
rect 4948 7800 4954 7812
rect 5350 7800 5356 7812
rect 4948 7772 5356 7800
rect 4948 7760 4954 7772
rect 5350 7760 5356 7772
rect 5408 7760 5414 7812
rect 5626 7760 5632 7812
rect 5684 7800 5690 7812
rect 6730 7800 6736 7812
rect 5684 7772 6736 7800
rect 5684 7760 5690 7772
rect 4430 7692 4436 7744
rect 4488 7732 4494 7744
rect 4982 7732 4988 7744
rect 4488 7704 4988 7732
rect 4488 7692 4494 7704
rect 4982 7692 4988 7704
rect 5040 7692 5046 7744
rect 5074 7692 5080 7744
rect 5132 7732 5138 7744
rect 5258 7732 5264 7744
rect 5132 7704 5264 7732
rect 5132 7692 5138 7704
rect 5258 7692 5264 7704
rect 5316 7692 5322 7744
rect 5828 7741 5856 7772
rect 6730 7760 6736 7772
rect 6788 7760 6794 7812
rect 7929 7803 7987 7809
rect 7929 7769 7941 7803
rect 7975 7800 7987 7803
rect 8205 7803 8263 7809
rect 8205 7800 8217 7803
rect 7975 7772 8217 7800
rect 7975 7769 7987 7772
rect 7929 7763 7987 7769
rect 8205 7769 8217 7772
rect 8251 7769 8263 7803
rect 8588 7800 8616 7828
rect 9582 7800 9588 7812
rect 8588 7772 9588 7800
rect 8205 7763 8263 7769
rect 9582 7760 9588 7772
rect 9640 7800 9646 7812
rect 9968 7800 9996 7831
rect 10042 7828 10048 7880
rect 10100 7868 10106 7880
rect 10137 7871 10195 7877
rect 10137 7868 10149 7871
rect 10100 7840 10149 7868
rect 10100 7828 10106 7840
rect 10137 7837 10149 7840
rect 10183 7837 10195 7871
rect 10137 7831 10195 7837
rect 11330 7828 11336 7880
rect 11388 7828 11394 7880
rect 9640 7772 9996 7800
rect 9640 7760 9646 7772
rect 12526 7760 12532 7812
rect 12584 7760 12590 7812
rect 12728 7809 12756 7908
rect 13081 7905 13093 7908
rect 13127 7936 13139 7939
rect 13446 7936 13452 7948
rect 13127 7908 13452 7936
rect 13127 7905 13139 7908
rect 13081 7899 13139 7905
rect 13446 7896 13452 7908
rect 13504 7896 13510 7948
rect 13817 7939 13875 7945
rect 13817 7905 13829 7939
rect 13863 7936 13875 7939
rect 13998 7936 14004 7948
rect 13863 7908 14004 7936
rect 13863 7905 13875 7908
rect 13817 7899 13875 7905
rect 13998 7896 14004 7908
rect 14056 7896 14062 7948
rect 20438 7936 20444 7948
rect 19628 7908 20444 7936
rect 19628 7880 19656 7908
rect 20438 7896 20444 7908
rect 20496 7896 20502 7948
rect 24121 7939 24179 7945
rect 24121 7905 24133 7939
rect 24167 7936 24179 7939
rect 24210 7936 24216 7948
rect 24167 7908 24216 7936
rect 24167 7905 24179 7908
rect 24121 7899 24179 7905
rect 24210 7896 24216 7908
rect 24268 7896 24274 7948
rect 12894 7828 12900 7880
rect 12952 7868 12958 7880
rect 13173 7871 13231 7877
rect 13173 7868 13185 7871
rect 12952 7840 13185 7868
rect 12952 7828 12958 7840
rect 13173 7837 13185 7840
rect 13219 7837 13231 7871
rect 13173 7831 13231 7837
rect 13357 7871 13415 7877
rect 13357 7837 13369 7871
rect 13403 7837 13415 7871
rect 13357 7831 13415 7837
rect 12728 7803 12787 7809
rect 12728 7772 12741 7803
rect 12729 7769 12741 7772
rect 12775 7769 12787 7803
rect 13262 7800 13268 7812
rect 12729 7763 12787 7769
rect 12820 7772 13268 7800
rect 5813 7735 5871 7741
rect 5813 7701 5825 7735
rect 5859 7701 5871 7735
rect 5813 7695 5871 7701
rect 6546 7692 6552 7744
rect 6604 7732 6610 7744
rect 8113 7735 8171 7741
rect 8113 7732 8125 7735
rect 6604 7704 8125 7732
rect 6604 7692 6610 7704
rect 8113 7701 8125 7704
rect 8159 7701 8171 7735
rect 8113 7695 8171 7701
rect 8662 7692 8668 7744
rect 8720 7732 8726 7744
rect 8941 7735 8999 7741
rect 8941 7732 8953 7735
rect 8720 7704 8953 7732
rect 8720 7692 8726 7704
rect 8941 7701 8953 7704
rect 8987 7701 8999 7735
rect 8941 7695 8999 7701
rect 9490 7692 9496 7744
rect 9548 7692 9554 7744
rect 12069 7735 12127 7741
rect 12069 7701 12081 7735
rect 12115 7732 12127 7735
rect 12158 7732 12164 7744
rect 12115 7704 12164 7732
rect 12115 7701 12127 7704
rect 12069 7695 12127 7701
rect 12158 7692 12164 7704
rect 12216 7692 12222 7744
rect 12544 7732 12572 7760
rect 12820 7732 12848 7772
rect 13262 7760 13268 7772
rect 13320 7800 13326 7812
rect 13372 7800 13400 7831
rect 13630 7828 13636 7880
rect 13688 7868 13694 7880
rect 14185 7871 14243 7877
rect 14185 7868 14197 7871
rect 13688 7840 14197 7868
rect 13688 7828 13694 7840
rect 14185 7837 14197 7840
rect 14231 7837 14243 7871
rect 14185 7831 14243 7837
rect 14553 7871 14611 7877
rect 14553 7837 14565 7871
rect 14599 7868 14611 7871
rect 14645 7871 14703 7877
rect 14645 7868 14657 7871
rect 14599 7840 14657 7868
rect 14599 7837 14611 7840
rect 14553 7831 14611 7837
rect 14645 7837 14657 7840
rect 14691 7837 14703 7871
rect 14921 7871 14979 7877
rect 14921 7868 14933 7871
rect 14645 7831 14703 7837
rect 14752 7840 14933 7868
rect 13320 7772 13400 7800
rect 13320 7760 13326 7772
rect 13722 7760 13728 7812
rect 13780 7800 13786 7812
rect 14369 7803 14427 7809
rect 14369 7800 14381 7803
rect 13780 7772 14381 7800
rect 13780 7760 13786 7772
rect 14369 7769 14381 7772
rect 14415 7800 14427 7803
rect 14752 7800 14780 7840
rect 14921 7837 14933 7840
rect 14967 7837 14979 7871
rect 14921 7831 14979 7837
rect 15018 7871 15076 7877
rect 15018 7837 15030 7871
rect 15064 7837 15076 7871
rect 15018 7831 15076 7837
rect 14415 7772 14780 7800
rect 14415 7769 14427 7772
rect 14369 7763 14427 7769
rect 14826 7760 14832 7812
rect 14884 7760 14890 7812
rect 12544 7704 12848 7732
rect 12897 7735 12955 7741
rect 12897 7701 12909 7735
rect 12943 7732 12955 7735
rect 14918 7732 14924 7744
rect 12943 7704 14924 7732
rect 12943 7701 12955 7704
rect 12897 7695 12955 7701
rect 14918 7692 14924 7704
rect 14976 7732 14982 7744
rect 15028 7732 15056 7831
rect 17586 7828 17592 7880
rect 17644 7828 17650 7880
rect 17865 7871 17923 7877
rect 17865 7837 17877 7871
rect 17911 7868 17923 7871
rect 18046 7868 18052 7880
rect 17911 7840 18052 7868
rect 17911 7837 17923 7840
rect 17865 7831 17923 7837
rect 18046 7828 18052 7840
rect 18104 7828 18110 7880
rect 19610 7828 19616 7880
rect 19668 7828 19674 7880
rect 19794 7828 19800 7880
rect 19852 7828 19858 7880
rect 21266 7828 21272 7880
rect 21324 7868 21330 7880
rect 22097 7871 22155 7877
rect 22097 7868 22109 7871
rect 21324 7840 22109 7868
rect 21324 7828 21330 7840
rect 22097 7837 22109 7840
rect 22143 7837 22155 7871
rect 22097 7831 22155 7837
rect 22278 7828 22284 7880
rect 22336 7828 22342 7880
rect 22370 7828 22376 7880
rect 22428 7868 22434 7880
rect 22557 7871 22615 7877
rect 22557 7868 22569 7871
rect 22428 7840 22569 7868
rect 22428 7828 22434 7840
rect 22557 7837 22569 7840
rect 22603 7837 22615 7871
rect 22557 7831 22615 7837
rect 23474 7828 23480 7880
rect 23532 7868 23538 7880
rect 23661 7871 23719 7877
rect 23661 7868 23673 7871
rect 23532 7840 23673 7868
rect 23532 7828 23538 7840
rect 23661 7837 23673 7840
rect 23707 7837 23719 7871
rect 23661 7831 23719 7837
rect 17310 7760 17316 7812
rect 17368 7800 17374 7812
rect 17494 7800 17500 7812
rect 17368 7772 17500 7800
rect 17368 7760 17374 7772
rect 17494 7760 17500 7772
rect 17552 7800 17558 7812
rect 17681 7803 17739 7809
rect 17681 7800 17693 7803
rect 17552 7772 17693 7800
rect 17552 7760 17558 7772
rect 17681 7769 17693 7772
rect 17727 7769 17739 7803
rect 17681 7763 17739 7769
rect 20073 7803 20131 7809
rect 20073 7769 20085 7803
rect 20119 7800 20131 7803
rect 21082 7800 21088 7812
rect 20119 7772 21088 7800
rect 20119 7769 20131 7772
rect 20073 7763 20131 7769
rect 21082 7760 21088 7772
rect 21140 7760 21146 7812
rect 23385 7803 23443 7809
rect 23385 7769 23397 7803
rect 23431 7800 23443 7803
rect 24302 7800 24308 7812
rect 23431 7772 24308 7800
rect 23431 7769 23443 7772
rect 23385 7763 23443 7769
rect 24302 7760 24308 7772
rect 24360 7760 24366 7812
rect 14976 7704 15056 7732
rect 14976 7692 14982 7704
rect 18046 7692 18052 7744
rect 18104 7692 18110 7744
rect 19978 7692 19984 7744
rect 20036 7692 20042 7744
rect 22922 7692 22928 7744
rect 22980 7732 22986 7744
rect 23753 7735 23811 7741
rect 23753 7732 23765 7735
rect 22980 7704 23765 7732
rect 22980 7692 22986 7704
rect 23753 7701 23765 7704
rect 23799 7701 23811 7735
rect 23753 7695 23811 7701
rect 23842 7692 23848 7744
rect 23900 7692 23906 7744
rect 1104 7642 27876 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 27876 7642
rect 1104 7568 27876 7590
rect 4525 7531 4583 7537
rect 4525 7497 4537 7531
rect 4571 7528 4583 7531
rect 4614 7528 4620 7540
rect 4571 7500 4620 7528
rect 4571 7497 4583 7500
rect 4525 7491 4583 7497
rect 4614 7488 4620 7500
rect 4672 7488 4678 7540
rect 4893 7531 4951 7537
rect 4893 7497 4905 7531
rect 4939 7528 4951 7531
rect 5258 7528 5264 7540
rect 4939 7500 5264 7528
rect 4939 7497 4951 7500
rect 4893 7491 4951 7497
rect 5258 7488 5264 7500
rect 5316 7488 5322 7540
rect 6638 7528 6644 7540
rect 5828 7500 6644 7528
rect 4154 7420 4160 7472
rect 4212 7460 4218 7472
rect 5828 7469 5856 7500
rect 6638 7488 6644 7500
rect 6696 7528 6702 7540
rect 6733 7531 6791 7537
rect 6733 7528 6745 7531
rect 6696 7500 6745 7528
rect 6696 7488 6702 7500
rect 6733 7497 6745 7500
rect 6779 7497 6791 7531
rect 11054 7528 11060 7540
rect 6733 7491 6791 7497
rect 7300 7500 11060 7528
rect 5813 7463 5871 7469
rect 4212 7432 4752 7460
rect 4212 7420 4218 7432
rect 4430 7352 4436 7404
rect 4488 7352 4494 7404
rect 4614 7352 4620 7404
rect 4672 7352 4678 7404
rect 4724 7401 4752 7432
rect 5813 7429 5825 7463
rect 5859 7429 5871 7463
rect 5813 7423 5871 7429
rect 5905 7463 5963 7469
rect 5905 7429 5917 7463
rect 5951 7460 5963 7463
rect 7193 7463 7251 7469
rect 7193 7460 7205 7463
rect 5951 7432 7205 7460
rect 5951 7429 5963 7432
rect 5905 7423 5963 7429
rect 4709 7395 4767 7401
rect 4709 7361 4721 7395
rect 4755 7361 4767 7395
rect 4709 7355 4767 7361
rect 5537 7395 5595 7401
rect 5537 7361 5549 7395
rect 5583 7361 5595 7395
rect 5537 7355 5595 7361
rect 5629 7395 5687 7401
rect 5629 7361 5641 7395
rect 5675 7392 5687 7395
rect 5718 7392 5724 7404
rect 5675 7364 5724 7392
rect 5675 7361 5687 7364
rect 5629 7355 5687 7361
rect 4448 7256 4476 7352
rect 4724 7324 4752 7355
rect 5552 7324 5580 7355
rect 5718 7352 5724 7364
rect 5776 7352 5782 7404
rect 6380 7401 6408 7432
rect 7193 7429 7205 7432
rect 7239 7429 7251 7463
rect 7193 7423 7251 7429
rect 5997 7395 6055 7401
rect 5997 7361 6009 7395
rect 6043 7361 6055 7395
rect 5997 7355 6055 7361
rect 6365 7395 6423 7401
rect 6365 7361 6377 7395
rect 6411 7361 6423 7395
rect 6365 7355 6423 7361
rect 5810 7324 5816 7336
rect 4724 7296 5304 7324
rect 5552 7296 5816 7324
rect 4706 7256 4712 7268
rect 4448 7228 4712 7256
rect 4706 7216 4712 7228
rect 4764 7216 4770 7268
rect 5276 7188 5304 7296
rect 5810 7284 5816 7296
rect 5868 7284 5874 7336
rect 6012 7324 6040 7355
rect 6546 7352 6552 7404
rect 6604 7352 6610 7404
rect 6641 7395 6699 7401
rect 6641 7361 6653 7395
rect 6687 7361 6699 7395
rect 6641 7355 6699 7361
rect 6564 7324 6592 7352
rect 6012 7296 6592 7324
rect 5350 7216 5356 7268
rect 5408 7256 5414 7268
rect 6181 7259 6239 7265
rect 6181 7256 6193 7259
rect 5408 7228 6193 7256
rect 5408 7216 5414 7228
rect 6181 7225 6193 7228
rect 6227 7225 6239 7259
rect 6181 7219 6239 7225
rect 6270 7216 6276 7268
rect 6328 7256 6334 7268
rect 6457 7259 6515 7265
rect 6457 7256 6469 7259
rect 6328 7228 6469 7256
rect 6328 7216 6334 7228
rect 6457 7225 6469 7228
rect 6503 7225 6515 7259
rect 6457 7219 6515 7225
rect 6546 7216 6552 7268
rect 6604 7256 6610 7268
rect 6656 7256 6684 7355
rect 6730 7352 6736 7404
rect 6788 7392 6794 7404
rect 7300 7392 7328 7500
rect 7837 7463 7895 7469
rect 7837 7460 7849 7463
rect 7392 7432 7849 7460
rect 7392 7401 7420 7432
rect 7837 7429 7849 7432
rect 7883 7429 7895 7463
rect 8386 7460 8392 7472
rect 7837 7423 7895 7429
rect 7944 7432 8392 7460
rect 6788 7364 7328 7392
rect 7377 7395 7435 7401
rect 6788 7352 6794 7364
rect 7377 7361 7389 7395
rect 7423 7361 7435 7395
rect 7377 7355 7435 7361
rect 7466 7352 7472 7404
rect 7524 7392 7530 7404
rect 7944 7401 7972 7432
rect 8386 7420 8392 7432
rect 8444 7420 8450 7472
rect 8496 7469 8524 7500
rect 11054 7488 11060 7500
rect 11112 7488 11118 7540
rect 13633 7531 13691 7537
rect 13633 7497 13645 7531
rect 13679 7528 13691 7531
rect 15010 7528 15016 7540
rect 13679 7500 15016 7528
rect 13679 7497 13691 7500
rect 13633 7491 13691 7497
rect 15010 7488 15016 7500
rect 15068 7488 15074 7540
rect 17586 7488 17592 7540
rect 17644 7488 17650 7540
rect 18785 7531 18843 7537
rect 18785 7497 18797 7531
rect 18831 7528 18843 7531
rect 19610 7528 19616 7540
rect 18831 7500 19616 7528
rect 18831 7497 18843 7500
rect 18785 7491 18843 7497
rect 19610 7488 19616 7500
rect 19668 7488 19674 7540
rect 21174 7488 21180 7540
rect 21232 7488 21238 7540
rect 22370 7488 22376 7540
rect 22428 7528 22434 7540
rect 23017 7531 23075 7537
rect 23017 7528 23029 7531
rect 22428 7500 23029 7528
rect 22428 7488 22434 7500
rect 23017 7497 23029 7500
rect 23063 7528 23075 7531
rect 23474 7528 23480 7540
rect 23063 7500 23480 7528
rect 23063 7497 23075 7500
rect 23017 7491 23075 7497
rect 23474 7488 23480 7500
rect 23532 7488 23538 7540
rect 24946 7488 24952 7540
rect 25004 7488 25010 7540
rect 25685 7531 25743 7537
rect 25685 7497 25697 7531
rect 25731 7528 25743 7531
rect 25774 7528 25780 7540
rect 25731 7500 25780 7528
rect 25731 7497 25743 7500
rect 25685 7491 25743 7497
rect 25774 7488 25780 7500
rect 25832 7488 25838 7540
rect 8481 7463 8539 7469
rect 8481 7429 8493 7463
rect 8527 7429 8539 7463
rect 8481 7423 8539 7429
rect 8573 7463 8631 7469
rect 8573 7429 8585 7463
rect 8619 7460 8631 7463
rect 9490 7460 9496 7472
rect 8619 7432 9496 7460
rect 8619 7429 8631 7432
rect 8573 7423 8631 7429
rect 7745 7395 7803 7401
rect 7745 7392 7757 7395
rect 7524 7364 7757 7392
rect 7524 7352 7530 7364
rect 7745 7361 7757 7364
rect 7791 7361 7803 7395
rect 7745 7355 7803 7361
rect 7929 7395 7987 7401
rect 7929 7361 7941 7395
rect 7975 7361 7987 7395
rect 7929 7355 7987 7361
rect 7650 7284 7656 7336
rect 7708 7284 7714 7336
rect 7760 7324 7788 7355
rect 8294 7352 8300 7404
rect 8352 7352 8358 7404
rect 8110 7324 8116 7336
rect 7760 7296 8116 7324
rect 8110 7284 8116 7296
rect 8168 7284 8174 7336
rect 6604 7228 6684 7256
rect 7561 7259 7619 7265
rect 6604 7216 6610 7228
rect 7561 7225 7573 7259
rect 7607 7256 7619 7259
rect 8588 7256 8616 7423
rect 9490 7420 9496 7432
rect 9548 7420 9554 7472
rect 9858 7420 9864 7472
rect 9916 7460 9922 7472
rect 11238 7460 11244 7472
rect 9916 7432 10732 7460
rect 9916 7420 9922 7432
rect 8662 7352 8668 7404
rect 8720 7352 8726 7404
rect 9953 7395 10011 7401
rect 9953 7361 9965 7395
rect 9999 7392 10011 7395
rect 10042 7392 10048 7404
rect 9999 7364 10048 7392
rect 9999 7361 10011 7364
rect 9953 7355 10011 7361
rect 10042 7352 10048 7364
rect 10100 7352 10106 7404
rect 10704 7401 10732 7432
rect 10888 7432 11244 7460
rect 10888 7401 10916 7432
rect 11238 7420 11244 7432
rect 11296 7420 11302 7472
rect 12986 7420 12992 7472
rect 13044 7460 13050 7472
rect 13044 7432 13676 7460
rect 13044 7420 13050 7432
rect 13648 7404 13676 7432
rect 14826 7420 14832 7472
rect 14884 7420 14890 7472
rect 17604 7460 17632 7488
rect 17236 7432 17632 7460
rect 20809 7463 20867 7469
rect 10689 7395 10747 7401
rect 10689 7361 10701 7395
rect 10735 7361 10747 7395
rect 10689 7355 10747 7361
rect 10873 7395 10931 7401
rect 10873 7361 10885 7395
rect 10919 7361 10931 7395
rect 10873 7355 10931 7361
rect 10704 7324 10732 7355
rect 10962 7352 10968 7404
rect 11020 7352 11026 7404
rect 11793 7395 11851 7401
rect 11793 7392 11805 7395
rect 11072 7364 11805 7392
rect 11072 7324 11100 7364
rect 11793 7361 11805 7364
rect 11839 7361 11851 7395
rect 11793 7355 11851 7361
rect 12066 7352 12072 7404
rect 12124 7392 12130 7404
rect 12713 7395 12771 7401
rect 12713 7392 12725 7395
rect 12124 7364 12725 7392
rect 12124 7352 12130 7364
rect 12713 7361 12725 7364
rect 12759 7361 12771 7395
rect 12713 7355 12771 7361
rect 13170 7352 13176 7404
rect 13228 7352 13234 7404
rect 13262 7352 13268 7404
rect 13320 7352 13326 7404
rect 13357 7395 13415 7401
rect 13357 7361 13369 7395
rect 13403 7392 13415 7395
rect 13538 7392 13544 7404
rect 13403 7364 13544 7392
rect 13403 7361 13415 7364
rect 13357 7355 13415 7361
rect 11701 7327 11759 7333
rect 11701 7324 11713 7327
rect 10704 7296 11100 7324
rect 11256 7296 11713 7324
rect 10962 7256 10968 7268
rect 7607 7228 8616 7256
rect 8772 7228 10968 7256
rect 7607 7225 7619 7228
rect 7561 7219 7619 7225
rect 8772 7188 8800 7228
rect 10962 7216 10968 7228
rect 11020 7216 11026 7268
rect 11256 7265 11284 7296
rect 11701 7293 11713 7296
rect 11747 7293 11759 7327
rect 11701 7287 11759 7293
rect 12621 7327 12679 7333
rect 12621 7293 12633 7327
rect 12667 7293 12679 7327
rect 12621 7287 12679 7293
rect 11241 7259 11299 7265
rect 11241 7225 11253 7259
rect 11287 7225 11299 7259
rect 12636 7256 12664 7287
rect 12894 7284 12900 7336
rect 12952 7324 12958 7336
rect 13372 7324 13400 7355
rect 13538 7352 13544 7364
rect 13596 7352 13602 7404
rect 13630 7352 13636 7404
rect 13688 7392 13694 7404
rect 14277 7395 14335 7401
rect 14277 7392 14289 7395
rect 13688 7364 14289 7392
rect 13688 7352 13694 7364
rect 14277 7361 14289 7364
rect 14323 7361 14335 7395
rect 14277 7355 14335 7361
rect 14461 7395 14519 7401
rect 14461 7361 14473 7395
rect 14507 7361 14519 7395
rect 14461 7355 14519 7361
rect 14737 7395 14795 7401
rect 14737 7361 14749 7395
rect 14783 7392 14795 7395
rect 14844 7392 14872 7420
rect 17236 7404 17264 7432
rect 20809 7429 20821 7463
rect 20855 7460 20867 7463
rect 20855 7432 22094 7460
rect 20855 7429 20867 7432
rect 20809 7423 20867 7429
rect 15197 7395 15255 7401
rect 15197 7392 15209 7395
rect 14783 7364 15209 7392
rect 14783 7361 14795 7364
rect 14737 7355 14795 7361
rect 15197 7361 15209 7364
rect 15243 7361 15255 7395
rect 15197 7355 15255 7361
rect 15381 7395 15439 7401
rect 15381 7361 15393 7395
rect 15427 7361 15439 7395
rect 15381 7355 15439 7361
rect 12952 7296 13400 7324
rect 12952 7284 12958 7296
rect 13446 7284 13452 7336
rect 13504 7284 13510 7336
rect 13722 7284 13728 7336
rect 13780 7324 13786 7336
rect 14476 7324 14504 7355
rect 13780 7296 14504 7324
rect 14829 7327 14887 7333
rect 13780 7284 13786 7296
rect 14829 7293 14841 7327
rect 14875 7324 14887 7327
rect 14918 7324 14924 7336
rect 14875 7296 14924 7324
rect 14875 7293 14887 7296
rect 14829 7287 14887 7293
rect 14918 7284 14924 7296
rect 14976 7284 14982 7336
rect 12710 7256 12716 7268
rect 12636 7228 12716 7256
rect 11241 7219 11299 7225
rect 12710 7216 12716 7228
rect 12768 7216 12774 7268
rect 13262 7216 13268 7268
rect 13320 7256 13326 7268
rect 15396 7256 15424 7355
rect 17218 7352 17224 7404
rect 17276 7352 17282 7404
rect 17310 7352 17316 7404
rect 17368 7352 17374 7404
rect 17497 7395 17555 7401
rect 17497 7361 17509 7395
rect 17543 7361 17555 7395
rect 17497 7355 17555 7361
rect 17589 7395 17647 7401
rect 17589 7361 17601 7395
rect 17635 7392 17647 7395
rect 17862 7392 17868 7404
rect 17635 7364 17868 7392
rect 17635 7361 17647 7364
rect 17589 7355 17647 7361
rect 16114 7284 16120 7336
rect 16172 7324 16178 7336
rect 16209 7327 16267 7333
rect 16209 7324 16221 7327
rect 16172 7296 16221 7324
rect 16172 7284 16178 7296
rect 16209 7293 16221 7296
rect 16255 7324 16267 7327
rect 17512 7324 17540 7355
rect 17862 7352 17868 7364
rect 17920 7352 17926 7404
rect 17957 7395 18015 7401
rect 17957 7361 17969 7395
rect 18003 7361 18015 7395
rect 17957 7355 18015 7361
rect 17972 7324 18000 7355
rect 19794 7352 19800 7404
rect 19852 7352 19858 7404
rect 19978 7352 19984 7404
rect 20036 7352 20042 7404
rect 21082 7352 21088 7404
rect 21140 7401 21146 7404
rect 21140 7395 21173 7401
rect 21161 7361 21173 7395
rect 21140 7355 21173 7361
rect 21499 7395 21557 7401
rect 21499 7361 21511 7395
rect 21545 7392 21557 7395
rect 22066 7392 22094 7432
rect 22646 7420 22652 7472
rect 22704 7460 22710 7472
rect 22833 7463 22891 7469
rect 22833 7460 22845 7463
rect 22704 7432 22845 7460
rect 22704 7420 22710 7432
rect 22833 7429 22845 7432
rect 22879 7429 22891 7463
rect 22833 7423 22891 7429
rect 22922 7420 22928 7472
rect 22980 7460 22986 7472
rect 23109 7463 23167 7469
rect 23109 7460 23121 7463
rect 22980 7432 23121 7460
rect 22980 7420 22986 7432
rect 23109 7429 23121 7432
rect 23155 7429 23167 7463
rect 23109 7423 23167 7429
rect 25222 7420 25228 7472
rect 25280 7460 25286 7472
rect 25869 7463 25927 7469
rect 25869 7460 25881 7463
rect 25280 7432 25881 7460
rect 25280 7420 25286 7432
rect 25869 7429 25881 7432
rect 25915 7429 25927 7463
rect 25869 7423 25927 7429
rect 22940 7392 22968 7420
rect 23201 7395 23259 7401
rect 23201 7392 23213 7395
rect 21545 7364 21864 7392
rect 22066 7364 22968 7392
rect 23032 7364 23213 7392
rect 21545 7361 21557 7364
rect 21499 7355 21557 7361
rect 21140 7352 21146 7355
rect 16255 7296 18000 7324
rect 16255 7293 16267 7296
rect 16209 7287 16267 7293
rect 18046 7284 18052 7336
rect 18104 7284 18110 7336
rect 21634 7284 21640 7336
rect 21692 7284 21698 7336
rect 13320 7228 15424 7256
rect 20993 7259 21051 7265
rect 13320 7216 13326 7228
rect 20993 7225 21005 7259
rect 21039 7256 21051 7259
rect 21836 7256 21864 7364
rect 22094 7256 22100 7268
rect 21039 7228 21680 7256
rect 21836 7228 22100 7256
rect 21039 7225 21051 7228
rect 20993 7219 21051 7225
rect 5276 7160 8800 7188
rect 8846 7148 8852 7200
rect 8904 7148 8910 7200
rect 10045 7191 10103 7197
rect 10045 7157 10057 7191
rect 10091 7188 10103 7191
rect 10686 7188 10692 7200
rect 10091 7160 10692 7188
rect 10091 7157 10103 7160
rect 10045 7151 10103 7157
rect 10686 7148 10692 7160
rect 10744 7148 10750 7200
rect 10870 7148 10876 7200
rect 10928 7148 10934 7200
rect 12805 7191 12863 7197
rect 12805 7157 12817 7191
rect 12851 7188 12863 7191
rect 13170 7188 13176 7200
rect 12851 7160 13176 7188
rect 12851 7157 12863 7160
rect 12805 7151 12863 7157
rect 13170 7148 13176 7160
rect 13228 7188 13234 7200
rect 13722 7188 13728 7200
rect 13228 7160 13728 7188
rect 13228 7148 13234 7160
rect 13722 7148 13728 7160
rect 13780 7148 13786 7200
rect 17034 7148 17040 7200
rect 17092 7148 17098 7200
rect 21652 7188 21680 7228
rect 22094 7216 22100 7228
rect 22152 7256 22158 7268
rect 22278 7256 22284 7268
rect 22152 7228 22284 7256
rect 22152 7216 22158 7228
rect 22278 7216 22284 7228
rect 22336 7216 22342 7268
rect 23032 7188 23060 7364
rect 23201 7361 23213 7364
rect 23247 7392 23259 7395
rect 23842 7392 23848 7404
rect 23247 7364 23848 7392
rect 23247 7361 23259 7364
rect 23201 7355 23259 7361
rect 23842 7352 23848 7364
rect 23900 7352 23906 7404
rect 24118 7352 24124 7404
rect 24176 7352 24182 7404
rect 24302 7352 24308 7404
rect 24360 7352 24366 7404
rect 25130 7352 25136 7404
rect 25188 7392 25194 7404
rect 25317 7395 25375 7401
rect 25317 7392 25329 7395
rect 25188 7364 25329 7392
rect 25188 7352 25194 7364
rect 25317 7361 25329 7364
rect 25363 7361 25375 7395
rect 25317 7355 25375 7361
rect 25590 7352 25596 7404
rect 25648 7352 25654 7404
rect 23750 7284 23756 7336
rect 23808 7324 23814 7336
rect 24029 7327 24087 7333
rect 24029 7324 24041 7327
rect 23808 7296 24041 7324
rect 23808 7284 23814 7296
rect 24029 7293 24041 7296
rect 24075 7324 24087 7327
rect 24486 7324 24492 7336
rect 24075 7296 24492 7324
rect 24075 7293 24087 7296
rect 24029 7287 24087 7293
rect 24486 7284 24492 7296
rect 24544 7284 24550 7336
rect 25409 7327 25467 7333
rect 25409 7293 25421 7327
rect 25455 7324 25467 7327
rect 25455 7296 25912 7324
rect 25455 7293 25467 7296
rect 25409 7287 25467 7293
rect 25884 7268 25912 7296
rect 25866 7216 25872 7268
rect 25924 7216 25930 7268
rect 21652 7160 23060 7188
rect 23382 7148 23388 7200
rect 23440 7148 23446 7200
rect 24489 7191 24547 7197
rect 24489 7157 24501 7191
rect 24535 7188 24547 7191
rect 25222 7188 25228 7200
rect 24535 7160 25228 7188
rect 24535 7157 24547 7160
rect 24489 7151 24547 7157
rect 25222 7148 25228 7160
rect 25280 7148 25286 7200
rect 1104 7098 27876 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 27876 7098
rect 1104 7024 27876 7046
rect 21085 6987 21143 6993
rect 21085 6953 21097 6987
rect 21131 6984 21143 6987
rect 21174 6984 21180 6996
rect 21131 6956 21180 6984
rect 21131 6953 21143 6956
rect 21085 6947 21143 6953
rect 21174 6944 21180 6956
rect 21232 6944 21238 6996
rect 21542 6944 21548 6996
rect 21600 6944 21606 6996
rect 23750 6944 23756 6996
rect 23808 6944 23814 6996
rect 25038 6944 25044 6996
rect 25096 6984 25102 6996
rect 25590 6984 25596 6996
rect 25096 6956 25596 6984
rect 25096 6944 25102 6956
rect 25590 6944 25596 6956
rect 25648 6944 25654 6996
rect 6270 6876 6276 6928
rect 6328 6876 6334 6928
rect 8294 6876 8300 6928
rect 8352 6916 8358 6928
rect 8352 6888 10364 6916
rect 8352 6876 8358 6888
rect 6288 6848 6316 6876
rect 10336 6848 10364 6888
rect 10410 6876 10416 6928
rect 10468 6916 10474 6928
rect 11054 6916 11060 6928
rect 10468 6888 11060 6916
rect 10468 6876 10474 6888
rect 11054 6876 11060 6888
rect 11112 6876 11118 6928
rect 12158 6876 12164 6928
rect 12216 6916 12222 6928
rect 13262 6916 13268 6928
rect 12216 6888 13268 6916
rect 12216 6876 12222 6888
rect 13262 6876 13268 6888
rect 13320 6876 13326 6928
rect 17129 6919 17187 6925
rect 17129 6885 17141 6919
rect 17175 6916 17187 6919
rect 21634 6916 21640 6928
rect 17175 6888 21640 6916
rect 17175 6885 17187 6888
rect 17129 6879 17187 6885
rect 6012 6820 6500 6848
rect 6012 6789 6040 6820
rect 5997 6783 6055 6789
rect 5997 6749 6009 6783
rect 6043 6749 6055 6783
rect 5997 6743 6055 6749
rect 6181 6783 6239 6789
rect 6181 6749 6193 6783
rect 6227 6780 6239 6783
rect 6273 6783 6331 6789
rect 6273 6780 6285 6783
rect 6227 6752 6285 6780
rect 6227 6749 6239 6752
rect 6181 6743 6239 6749
rect 6273 6749 6285 6752
rect 6319 6780 6331 6783
rect 6362 6780 6368 6792
rect 6319 6752 6368 6780
rect 6319 6749 6331 6752
rect 6273 6743 6331 6749
rect 6362 6740 6368 6752
rect 6420 6740 6426 6792
rect 6472 6789 6500 6820
rect 10336 6820 11100 6848
rect 6457 6783 6515 6789
rect 6457 6749 6469 6783
rect 6503 6749 6515 6783
rect 6457 6743 6515 6749
rect 8846 6740 8852 6792
rect 8904 6780 8910 6792
rect 10336 6789 10364 6820
rect 9033 6783 9091 6789
rect 9033 6780 9045 6783
rect 8904 6752 9045 6780
rect 8904 6740 8910 6752
rect 9033 6749 9045 6752
rect 9079 6749 9091 6783
rect 9033 6743 9091 6749
rect 9217 6783 9275 6789
rect 9217 6749 9229 6783
rect 9263 6749 9275 6783
rect 9217 6743 9275 6749
rect 10321 6783 10379 6789
rect 10321 6749 10333 6783
rect 10367 6749 10379 6783
rect 10321 6743 10379 6749
rect 7650 6672 7656 6724
rect 7708 6712 7714 6724
rect 9232 6712 9260 6743
rect 10410 6740 10416 6792
rect 10468 6740 10474 6792
rect 10597 6783 10655 6789
rect 10597 6749 10609 6783
rect 10643 6749 10655 6783
rect 10597 6743 10655 6749
rect 7708 6684 9260 6712
rect 7708 6672 7714 6684
rect 9766 6672 9772 6724
rect 9824 6712 9830 6724
rect 10137 6715 10195 6721
rect 10137 6712 10149 6715
rect 9824 6684 10149 6712
rect 9824 6672 9830 6684
rect 10137 6681 10149 6684
rect 10183 6681 10195 6715
rect 10612 6712 10640 6743
rect 10686 6740 10692 6792
rect 10744 6740 10750 6792
rect 10781 6783 10839 6789
rect 10781 6749 10793 6783
rect 10827 6780 10839 6783
rect 10870 6780 10876 6792
rect 10827 6752 10876 6780
rect 10827 6749 10839 6752
rect 10781 6743 10839 6749
rect 10796 6712 10824 6743
rect 10870 6740 10876 6752
rect 10928 6740 10934 6792
rect 11072 6789 11100 6820
rect 15948 6820 16804 6848
rect 15948 6792 15976 6820
rect 11057 6783 11115 6789
rect 11057 6749 11069 6783
rect 11103 6780 11115 6783
rect 12342 6780 12348 6792
rect 11103 6752 12348 6780
rect 11103 6749 11115 6752
rect 11057 6743 11115 6749
rect 12342 6740 12348 6752
rect 12400 6740 12406 6792
rect 15930 6740 15936 6792
rect 15988 6740 15994 6792
rect 16114 6740 16120 6792
rect 16172 6740 16178 6792
rect 16298 6740 16304 6792
rect 16356 6740 16362 6792
rect 16776 6789 16804 6820
rect 16393 6783 16451 6789
rect 16393 6749 16405 6783
rect 16439 6749 16451 6783
rect 16393 6743 16451 6749
rect 16761 6783 16819 6789
rect 16761 6749 16773 6783
rect 16807 6749 16819 6783
rect 16761 6743 16819 6749
rect 10612 6684 10824 6712
rect 16025 6715 16083 6721
rect 10137 6675 10195 6681
rect 16025 6681 16037 6715
rect 16071 6712 16083 6715
rect 16408 6712 16436 6743
rect 17034 6740 17040 6792
rect 17092 6740 17098 6792
rect 17221 6783 17279 6789
rect 17221 6749 17233 6783
rect 17267 6749 17279 6783
rect 17221 6743 17279 6749
rect 16071 6684 16436 6712
rect 16577 6715 16635 6721
rect 16071 6681 16083 6684
rect 16025 6675 16083 6681
rect 16132 6656 16160 6684
rect 16577 6681 16589 6715
rect 16623 6712 16635 6715
rect 16850 6712 16856 6724
rect 16623 6684 16856 6712
rect 16623 6681 16635 6684
rect 16577 6675 16635 6681
rect 16850 6672 16856 6684
rect 16908 6712 16914 6724
rect 17236 6712 17264 6743
rect 17402 6740 17408 6792
rect 17460 6740 17466 6792
rect 18598 6740 18604 6792
rect 18656 6780 18662 6792
rect 19245 6783 19303 6789
rect 19245 6780 19257 6783
rect 18656 6752 19257 6780
rect 18656 6740 18662 6752
rect 19245 6749 19257 6752
rect 19291 6749 19303 6783
rect 19245 6743 19303 6749
rect 19610 6740 19616 6792
rect 19668 6780 19674 6792
rect 19705 6783 19763 6789
rect 19705 6780 19717 6783
rect 19668 6752 19717 6780
rect 19668 6740 19674 6752
rect 19705 6749 19717 6752
rect 19751 6749 19763 6783
rect 19705 6743 19763 6749
rect 19886 6740 19892 6792
rect 19944 6740 19950 6792
rect 20180 6789 20208 6888
rect 21634 6876 21640 6888
rect 21692 6876 21698 6928
rect 21729 6919 21787 6925
rect 21729 6885 21741 6919
rect 21775 6885 21787 6919
rect 21729 6879 21787 6885
rect 21358 6808 21364 6860
rect 21416 6808 21422 6860
rect 21744 6848 21772 6879
rect 22370 6876 22376 6928
rect 22428 6876 22434 6928
rect 25774 6916 25780 6928
rect 25240 6888 25780 6916
rect 21913 6851 21971 6857
rect 21913 6848 21925 6851
rect 21744 6820 21925 6848
rect 21913 6817 21925 6820
rect 21959 6817 21971 6851
rect 21913 6811 21971 6817
rect 24946 6808 24952 6860
rect 25004 6848 25010 6860
rect 25240 6848 25268 6888
rect 25774 6876 25780 6888
rect 25832 6876 25838 6928
rect 26237 6851 26295 6857
rect 26237 6848 26249 6851
rect 25004 6820 25268 6848
rect 25424 6820 26249 6848
rect 25004 6808 25010 6820
rect 20165 6783 20223 6789
rect 20165 6749 20177 6783
rect 20211 6749 20223 6783
rect 20165 6743 20223 6749
rect 20254 6740 20260 6792
rect 20312 6780 20318 6792
rect 21545 6783 21603 6789
rect 21545 6780 21557 6783
rect 20312 6752 21557 6780
rect 20312 6740 20318 6752
rect 21545 6749 21557 6752
rect 21591 6749 21603 6783
rect 21545 6743 21603 6749
rect 22005 6783 22063 6789
rect 22005 6749 22017 6783
rect 22051 6749 22063 6783
rect 22005 6743 22063 6749
rect 23293 6783 23351 6789
rect 23293 6749 23305 6783
rect 23339 6780 23351 6783
rect 23382 6780 23388 6792
rect 23339 6752 23388 6780
rect 23339 6749 23351 6752
rect 23293 6743 23351 6749
rect 16908 6684 17264 6712
rect 16908 6672 16914 6684
rect 18690 6672 18696 6724
rect 18748 6712 18754 6724
rect 18748 6684 20484 6712
rect 18748 6672 18754 6684
rect 6178 6604 6184 6656
rect 6236 6604 6242 6656
rect 6365 6647 6423 6653
rect 6365 6613 6377 6647
rect 6411 6644 6423 6647
rect 6730 6644 6736 6656
rect 6411 6616 6736 6644
rect 6411 6613 6423 6616
rect 6365 6607 6423 6613
rect 6730 6604 6736 6616
rect 6788 6604 6794 6656
rect 10045 6647 10103 6653
rect 10045 6613 10057 6647
rect 10091 6644 10103 6647
rect 10226 6644 10232 6656
rect 10091 6616 10232 6644
rect 10091 6613 10103 6616
rect 10045 6607 10103 6613
rect 10226 6604 10232 6616
rect 10284 6604 10290 6656
rect 10410 6604 10416 6656
rect 10468 6644 10474 6656
rect 10879 6647 10937 6653
rect 10879 6644 10891 6647
rect 10468 6616 10891 6644
rect 10468 6604 10474 6616
rect 10879 6613 10891 6616
rect 10925 6613 10937 6647
rect 10879 6607 10937 6613
rect 10965 6647 11023 6653
rect 10965 6613 10977 6647
rect 11011 6644 11023 6647
rect 11054 6644 11060 6656
rect 11011 6616 11060 6644
rect 11011 6613 11023 6616
rect 10965 6607 11023 6613
rect 11054 6604 11060 6616
rect 11112 6604 11118 6656
rect 16114 6604 16120 6656
rect 16172 6604 16178 6656
rect 19337 6647 19395 6653
rect 19337 6613 19349 6647
rect 19383 6644 19395 6647
rect 19794 6644 19800 6656
rect 19383 6616 19800 6644
rect 19383 6613 19395 6616
rect 19337 6607 19395 6613
rect 19794 6604 19800 6616
rect 19852 6644 19858 6656
rect 20254 6644 20260 6656
rect 19852 6616 20260 6644
rect 19852 6604 19858 6616
rect 20254 6604 20260 6616
rect 20312 6604 20318 6656
rect 20346 6604 20352 6656
rect 20404 6604 20410 6656
rect 20456 6644 20484 6684
rect 20714 6672 20720 6724
rect 20772 6672 20778 6724
rect 20898 6672 20904 6724
rect 20956 6672 20962 6724
rect 20990 6672 20996 6724
rect 21048 6712 21054 6724
rect 21269 6715 21327 6721
rect 21269 6712 21281 6715
rect 21048 6684 21281 6712
rect 21048 6672 21054 6684
rect 21269 6681 21281 6684
rect 21315 6681 21327 6715
rect 21269 6675 21327 6681
rect 22020 6644 22048 6743
rect 23382 6740 23388 6752
rect 23440 6740 23446 6792
rect 23566 6740 23572 6792
rect 23624 6740 23630 6792
rect 23750 6740 23756 6792
rect 23808 6740 23814 6792
rect 25038 6740 25044 6792
rect 25096 6740 25102 6792
rect 25148 6789 25176 6820
rect 25133 6783 25191 6789
rect 25133 6749 25145 6783
rect 25179 6749 25191 6783
rect 25133 6743 25191 6749
rect 25222 6740 25228 6792
rect 25280 6780 25286 6792
rect 25424 6789 25452 6820
rect 26237 6817 26249 6820
rect 26283 6817 26295 6851
rect 26237 6811 26295 6817
rect 25317 6783 25375 6789
rect 25317 6780 25329 6783
rect 25280 6752 25329 6780
rect 25280 6740 25286 6752
rect 25317 6749 25329 6752
rect 25363 6749 25375 6783
rect 25317 6743 25375 6749
rect 25409 6783 25467 6789
rect 25409 6749 25421 6783
rect 25455 6749 25467 6783
rect 25409 6743 25467 6749
rect 25501 6783 25559 6789
rect 25501 6749 25513 6783
rect 25547 6780 25559 6783
rect 25590 6780 25596 6792
rect 25547 6752 25596 6780
rect 25547 6749 25559 6752
rect 25501 6743 25559 6749
rect 25590 6740 25596 6752
rect 25648 6740 25654 6792
rect 25866 6740 25872 6792
rect 25924 6740 25930 6792
rect 26145 6783 26203 6789
rect 26145 6780 26157 6783
rect 25976 6752 26157 6780
rect 24857 6715 24915 6721
rect 24857 6681 24869 6715
rect 24903 6712 24915 6715
rect 25685 6715 25743 6721
rect 25685 6712 25697 6715
rect 24903 6684 25697 6712
rect 24903 6681 24915 6684
rect 24857 6675 24915 6681
rect 25685 6681 25697 6684
rect 25731 6681 25743 6715
rect 25685 6675 25743 6681
rect 25774 6672 25780 6724
rect 25832 6672 25838 6724
rect 20456 6616 22048 6644
rect 23658 6604 23664 6656
rect 23716 6644 23722 6656
rect 23937 6647 23995 6653
rect 23937 6644 23949 6647
rect 23716 6616 23949 6644
rect 23716 6604 23722 6616
rect 23937 6613 23949 6616
rect 23983 6613 23995 6647
rect 23937 6607 23995 6613
rect 25130 6604 25136 6656
rect 25188 6644 25194 6656
rect 25976 6644 26004 6752
rect 26145 6749 26157 6752
rect 26191 6749 26203 6783
rect 26145 6743 26203 6749
rect 25188 6616 26004 6644
rect 26053 6647 26111 6653
rect 25188 6604 25194 6616
rect 26053 6613 26065 6647
rect 26099 6644 26111 6647
rect 26142 6644 26148 6656
rect 26099 6616 26148 6644
rect 26099 6613 26111 6616
rect 26053 6607 26111 6613
rect 26142 6604 26148 6616
rect 26200 6604 26206 6656
rect 1104 6554 27876 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 27876 6554
rect 1104 6480 27876 6502
rect 4985 6443 5043 6449
rect 4985 6409 4997 6443
rect 5031 6440 5043 6443
rect 5626 6440 5632 6452
rect 5031 6412 5632 6440
rect 5031 6409 5043 6412
rect 4985 6403 5043 6409
rect 5626 6400 5632 6412
rect 5684 6400 5690 6452
rect 6730 6440 6736 6452
rect 5828 6412 6736 6440
rect 5828 6381 5856 6412
rect 6730 6400 6736 6412
rect 6788 6400 6794 6452
rect 7650 6400 7656 6452
rect 7708 6440 7714 6452
rect 8297 6443 8355 6449
rect 8297 6440 8309 6443
rect 7708 6412 8309 6440
rect 7708 6400 7714 6412
rect 8297 6409 8309 6412
rect 8343 6409 8355 6443
rect 12986 6440 12992 6452
rect 8297 6403 8355 6409
rect 12728 6412 12992 6440
rect 5813 6375 5871 6381
rect 5813 6372 5825 6375
rect 5368 6344 5825 6372
rect 4982 6307 5040 6313
rect 4982 6273 4994 6307
rect 5028 6304 5040 6307
rect 5258 6304 5264 6316
rect 5028 6276 5264 6304
rect 5028 6273 5040 6276
rect 4982 6267 5040 6273
rect 5258 6264 5264 6276
rect 5316 6264 5322 6316
rect 5368 6313 5396 6344
rect 5813 6341 5825 6344
rect 5859 6341 5871 6375
rect 5813 6335 5871 6341
rect 6638 6332 6644 6384
rect 6696 6332 6702 6384
rect 12066 6372 12072 6384
rect 11808 6344 12072 6372
rect 5353 6307 5411 6313
rect 5353 6273 5365 6307
rect 5399 6273 5411 6307
rect 5353 6267 5411 6273
rect 5534 6264 5540 6316
rect 5592 6264 5598 6316
rect 5718 6264 5724 6316
rect 5776 6264 5782 6316
rect 6178 6264 6184 6316
rect 6236 6304 6242 6316
rect 6365 6307 6423 6313
rect 6365 6304 6377 6307
rect 6236 6276 6377 6304
rect 6236 6264 6242 6276
rect 6365 6273 6377 6276
rect 6411 6273 6423 6307
rect 6365 6267 6423 6273
rect 6549 6307 6607 6313
rect 6549 6273 6561 6307
rect 6595 6273 6607 6307
rect 6549 6267 6607 6273
rect 6733 6307 6791 6313
rect 6733 6273 6745 6307
rect 6779 6304 6791 6307
rect 6822 6304 6828 6316
rect 6779 6276 6828 6304
rect 6779 6273 6791 6276
rect 6733 6267 6791 6273
rect 5445 6239 5503 6245
rect 5445 6205 5457 6239
rect 5491 6236 5503 6239
rect 5736 6236 5764 6264
rect 5994 6236 6000 6248
rect 5491 6208 6000 6236
rect 5491 6205 5503 6208
rect 5445 6199 5503 6205
rect 5994 6196 6000 6208
rect 6052 6196 6058 6248
rect 5718 6128 5724 6180
rect 5776 6168 5782 6180
rect 5813 6171 5871 6177
rect 5813 6168 5825 6171
rect 5776 6140 5825 6168
rect 5776 6128 5782 6140
rect 5813 6137 5825 6140
rect 5859 6168 5871 6171
rect 6564 6168 6592 6267
rect 6822 6264 6828 6276
rect 6880 6264 6886 6316
rect 7558 6264 7564 6316
rect 7616 6264 7622 6316
rect 7742 6264 7748 6316
rect 7800 6264 7806 6316
rect 10042 6264 10048 6316
rect 10100 6304 10106 6316
rect 11808 6313 11836 6344
rect 12066 6332 12072 6344
rect 12124 6332 12130 6384
rect 10321 6307 10379 6313
rect 10321 6304 10333 6307
rect 10100 6276 10333 6304
rect 10100 6264 10106 6276
rect 10321 6273 10333 6276
rect 10367 6273 10379 6307
rect 10321 6267 10379 6273
rect 11793 6307 11851 6313
rect 11793 6273 11805 6307
rect 11839 6273 11851 6307
rect 11793 6267 11851 6273
rect 11974 6264 11980 6316
rect 12032 6304 12038 6316
rect 12253 6307 12311 6313
rect 12253 6304 12265 6307
rect 12032 6276 12265 6304
rect 12032 6264 12038 6276
rect 12253 6273 12265 6276
rect 12299 6273 12311 6307
rect 12253 6267 12311 6273
rect 12437 6307 12495 6313
rect 12437 6273 12449 6307
rect 12483 6304 12495 6307
rect 12618 6304 12624 6316
rect 12483 6276 12624 6304
rect 12483 6273 12495 6276
rect 12437 6267 12495 6273
rect 12618 6264 12624 6276
rect 12676 6264 12682 6316
rect 12728 6313 12756 6412
rect 12986 6400 12992 6412
rect 13044 6400 13050 6452
rect 13814 6400 13820 6452
rect 13872 6400 13878 6452
rect 14737 6443 14795 6449
rect 14737 6409 14749 6443
rect 14783 6440 14795 6443
rect 14826 6440 14832 6452
rect 14783 6412 14832 6440
rect 14783 6409 14795 6412
rect 14737 6403 14795 6409
rect 14826 6400 14832 6412
rect 14884 6400 14890 6452
rect 14921 6443 14979 6449
rect 14921 6409 14933 6443
rect 14967 6409 14979 6443
rect 14921 6403 14979 6409
rect 15565 6443 15623 6449
rect 15565 6409 15577 6443
rect 15611 6440 15623 6443
rect 15930 6440 15936 6452
rect 15611 6412 15936 6440
rect 15611 6409 15623 6412
rect 15565 6403 15623 6409
rect 13541 6375 13599 6381
rect 13541 6372 13553 6375
rect 12820 6344 13553 6372
rect 12713 6307 12771 6313
rect 12713 6273 12725 6307
rect 12759 6273 12771 6307
rect 12713 6267 12771 6273
rect 10410 6196 10416 6248
rect 10468 6196 10474 6248
rect 11882 6196 11888 6248
rect 11940 6196 11946 6248
rect 5859 6140 6592 6168
rect 6917 6171 6975 6177
rect 5859 6137 5871 6140
rect 5813 6131 5871 6137
rect 6917 6137 6929 6171
rect 6963 6168 6975 6171
rect 9950 6168 9956 6180
rect 6963 6140 9956 6168
rect 6963 6137 6975 6140
rect 6917 6131 6975 6137
rect 9950 6128 9956 6140
rect 10008 6128 10014 6180
rect 10689 6171 10747 6177
rect 10689 6137 10701 6171
rect 10735 6168 10747 6171
rect 12161 6171 12219 6177
rect 10735 6140 11928 6168
rect 10735 6137 10747 6140
rect 10689 6131 10747 6137
rect 4798 6060 4804 6112
rect 4856 6060 4862 6112
rect 11790 6060 11796 6112
rect 11848 6060 11854 6112
rect 11900 6100 11928 6140
rect 12161 6137 12173 6171
rect 12207 6168 12219 6171
rect 12529 6171 12587 6177
rect 12529 6168 12541 6171
rect 12207 6140 12541 6168
rect 12207 6137 12219 6140
rect 12161 6131 12219 6137
rect 12529 6137 12541 6140
rect 12575 6137 12587 6171
rect 12529 6131 12587 6137
rect 12621 6171 12679 6177
rect 12621 6137 12633 6171
rect 12667 6168 12679 6171
rect 12820 6168 12848 6344
rect 13541 6341 13553 6344
rect 13587 6341 13599 6375
rect 13832 6372 13860 6400
rect 14001 6375 14059 6381
rect 14001 6372 14013 6375
rect 13832 6344 14013 6372
rect 13541 6335 13599 6341
rect 14001 6341 14013 6344
rect 14047 6372 14059 6375
rect 14366 6372 14372 6384
rect 14047 6344 14372 6372
rect 14047 6341 14059 6344
rect 14001 6335 14059 6341
rect 14366 6332 14372 6344
rect 14424 6332 14430 6384
rect 14936 6372 14964 6403
rect 15930 6400 15936 6412
rect 15988 6400 15994 6452
rect 16025 6443 16083 6449
rect 16025 6409 16037 6443
rect 16071 6440 16083 6443
rect 16298 6440 16304 6452
rect 16071 6412 16304 6440
rect 16071 6409 16083 6412
rect 16025 6403 16083 6409
rect 16298 6400 16304 6412
rect 16356 6400 16362 6452
rect 20990 6400 20996 6452
rect 21048 6400 21054 6452
rect 23566 6400 23572 6452
rect 23624 6440 23630 6452
rect 23661 6443 23719 6449
rect 23661 6440 23673 6443
rect 23624 6412 23673 6440
rect 23624 6400 23630 6412
rect 23661 6409 23673 6412
rect 23707 6440 23719 6443
rect 25409 6443 25467 6449
rect 23707 6412 25360 6440
rect 23707 6409 23719 6412
rect 23661 6403 23719 6409
rect 14936 6344 15884 6372
rect 15856 6316 15884 6344
rect 18690 6332 18696 6384
rect 18748 6332 18754 6384
rect 20898 6372 20904 6384
rect 20640 6344 20904 6372
rect 12986 6264 12992 6316
rect 13044 6264 13050 6316
rect 13081 6307 13139 6313
rect 13081 6273 13093 6307
rect 13127 6304 13139 6307
rect 13170 6304 13176 6316
rect 13127 6276 13176 6304
rect 13127 6273 13139 6276
rect 13081 6267 13139 6273
rect 13170 6264 13176 6276
rect 13228 6264 13234 6316
rect 13262 6264 13268 6316
rect 13320 6264 13326 6316
rect 13357 6307 13415 6313
rect 13357 6273 13369 6307
rect 13403 6273 13415 6307
rect 13357 6267 13415 6273
rect 13817 6307 13875 6313
rect 13817 6273 13829 6307
rect 13863 6273 13875 6307
rect 13817 6267 13875 6273
rect 13372 6236 13400 6267
rect 13832 6236 13860 6267
rect 14090 6264 14096 6316
rect 14148 6304 14154 6316
rect 14740 6307 14798 6313
rect 14740 6304 14752 6307
rect 14148 6276 14752 6304
rect 14148 6264 14154 6276
rect 14740 6273 14752 6276
rect 14786 6273 14798 6307
rect 14740 6267 14798 6273
rect 15194 6264 15200 6316
rect 15252 6264 15258 6316
rect 15838 6264 15844 6316
rect 15896 6264 15902 6316
rect 16114 6264 16120 6316
rect 16172 6264 16178 6316
rect 18414 6264 18420 6316
rect 18472 6313 18478 6316
rect 18472 6307 18521 6313
rect 18472 6273 18475 6307
rect 18509 6273 18521 6307
rect 18472 6267 18521 6273
rect 18472 6264 18478 6267
rect 18598 6264 18604 6316
rect 18656 6264 18662 6316
rect 20640 6313 20668 6344
rect 20898 6332 20904 6344
rect 20956 6332 20962 6384
rect 18785 6307 18843 6313
rect 18785 6273 18797 6307
rect 18831 6273 18843 6307
rect 18785 6267 18843 6273
rect 20625 6307 20683 6313
rect 20625 6273 20637 6307
rect 20671 6273 20683 6307
rect 20625 6267 20683 6273
rect 14277 6239 14335 6245
rect 14277 6236 14289 6239
rect 13280 6208 13860 6236
rect 14108 6208 14289 6236
rect 13078 6168 13084 6180
rect 12667 6140 13084 6168
rect 12667 6137 12679 6140
rect 12621 6131 12679 6137
rect 13078 6128 13084 6140
rect 13136 6128 13142 6180
rect 13280 6177 13308 6208
rect 13265 6171 13323 6177
rect 13265 6137 13277 6171
rect 13311 6137 13323 6171
rect 13265 6131 13323 6137
rect 12802 6100 12808 6112
rect 11900 6072 12808 6100
rect 12802 6060 12808 6072
rect 12860 6060 12866 6112
rect 12894 6060 12900 6112
rect 12952 6060 12958 6112
rect 13722 6060 13728 6112
rect 13780 6100 13786 6112
rect 14108 6100 14136 6208
rect 14277 6205 14289 6208
rect 14323 6205 14335 6239
rect 14277 6199 14335 6205
rect 14366 6196 14372 6248
rect 14424 6196 14430 6248
rect 15105 6239 15163 6245
rect 15105 6205 15117 6239
rect 15151 6205 15163 6239
rect 15105 6199 15163 6205
rect 14185 6171 14243 6177
rect 14185 6137 14197 6171
rect 14231 6168 14243 6171
rect 14458 6168 14464 6180
rect 14231 6140 14464 6168
rect 14231 6137 14243 6140
rect 14185 6131 14243 6137
rect 14458 6128 14464 6140
rect 14516 6168 14522 6180
rect 15120 6168 15148 6199
rect 18322 6196 18328 6248
rect 18380 6196 18386 6248
rect 14516 6140 15148 6168
rect 14516 6128 14522 6140
rect 13780 6072 14136 6100
rect 13780 6060 13786 6072
rect 15562 6060 15568 6112
rect 15620 6100 15626 6112
rect 15657 6103 15715 6109
rect 15657 6100 15669 6103
rect 15620 6072 15669 6100
rect 15620 6060 15626 6072
rect 15657 6069 15669 6072
rect 15703 6069 15715 6103
rect 18800 6100 18828 6267
rect 20714 6264 20720 6316
rect 20772 6304 20778 6316
rect 20809 6307 20867 6313
rect 20809 6304 20821 6307
rect 20772 6276 20821 6304
rect 20772 6264 20778 6276
rect 20809 6273 20821 6276
rect 20855 6273 20867 6307
rect 21008 6304 21036 6400
rect 23293 6375 23351 6381
rect 23293 6372 23305 6375
rect 21192 6344 23305 6372
rect 21085 6307 21143 6313
rect 21085 6304 21097 6307
rect 21008 6276 21097 6304
rect 20809 6267 20867 6273
rect 21085 6273 21097 6276
rect 21131 6273 21143 6307
rect 21085 6267 21143 6273
rect 21192 6236 21220 6344
rect 23293 6341 23305 6344
rect 23339 6372 23351 6375
rect 23339 6344 23980 6372
rect 23339 6341 23351 6344
rect 23293 6335 23351 6341
rect 21361 6307 21419 6313
rect 21361 6273 21373 6307
rect 21407 6304 21419 6307
rect 21542 6304 21548 6316
rect 21407 6276 21548 6304
rect 21407 6273 21419 6276
rect 21361 6267 21419 6273
rect 21542 6264 21548 6276
rect 21600 6304 21606 6316
rect 21910 6304 21916 6316
rect 21600 6276 21916 6304
rect 21600 6264 21606 6276
rect 21910 6264 21916 6276
rect 21968 6264 21974 6316
rect 23198 6264 23204 6316
rect 23256 6264 23262 6316
rect 23474 6264 23480 6316
rect 23532 6264 23538 6316
rect 23952 6313 23980 6344
rect 25332 6313 25360 6412
rect 25409 6409 25421 6443
rect 25455 6440 25467 6443
rect 25774 6440 25780 6452
rect 25455 6412 25780 6440
rect 25455 6409 25467 6412
rect 25409 6403 25467 6409
rect 25774 6400 25780 6412
rect 25832 6400 25838 6452
rect 23753 6307 23811 6313
rect 23753 6273 23765 6307
rect 23799 6273 23811 6307
rect 23753 6267 23811 6273
rect 23937 6307 23995 6313
rect 23937 6273 23949 6307
rect 23983 6273 23995 6307
rect 23937 6267 23995 6273
rect 25317 6307 25375 6313
rect 25317 6273 25329 6307
rect 25363 6273 25375 6307
rect 25317 6267 25375 6273
rect 21100 6208 21220 6236
rect 23216 6236 23244 6264
rect 23768 6236 23796 6267
rect 23216 6208 23796 6236
rect 23845 6239 23903 6245
rect 18969 6171 19027 6177
rect 18969 6137 18981 6171
rect 19015 6168 19027 6171
rect 21100 6168 21128 6208
rect 23845 6205 23857 6239
rect 23891 6236 23903 6239
rect 25130 6236 25136 6248
rect 23891 6208 25136 6236
rect 23891 6205 23903 6208
rect 23845 6199 23903 6205
rect 25130 6196 25136 6208
rect 25188 6196 25194 6248
rect 19015 6140 21128 6168
rect 21177 6171 21235 6177
rect 19015 6137 19027 6140
rect 18969 6131 19027 6137
rect 21177 6137 21189 6171
rect 21223 6168 21235 6171
rect 21358 6168 21364 6180
rect 21223 6140 21364 6168
rect 21223 6137 21235 6140
rect 21177 6131 21235 6137
rect 21358 6128 21364 6140
rect 21416 6168 21422 6180
rect 21818 6168 21824 6180
rect 21416 6140 21824 6168
rect 21416 6128 21422 6140
rect 21818 6128 21824 6140
rect 21876 6128 21882 6180
rect 23474 6128 23480 6180
rect 23532 6168 23538 6180
rect 25590 6168 25596 6180
rect 23532 6140 25596 6168
rect 23532 6128 23538 6140
rect 25590 6128 25596 6140
rect 25648 6128 25654 6180
rect 21082 6100 21088 6112
rect 18800 6072 21088 6100
rect 15657 6063 15715 6069
rect 21082 6060 21088 6072
rect 21140 6060 21146 6112
rect 1104 6010 27876 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 27876 6010
rect 1104 5936 27876 5958
rect 11241 5899 11299 5905
rect 11241 5865 11253 5899
rect 11287 5896 11299 5899
rect 11974 5896 11980 5908
rect 11287 5868 11980 5896
rect 11287 5865 11299 5868
rect 11241 5859 11299 5865
rect 11974 5856 11980 5868
rect 12032 5856 12038 5908
rect 12618 5856 12624 5908
rect 12676 5856 12682 5908
rect 12710 5856 12716 5908
rect 12768 5856 12774 5908
rect 13078 5856 13084 5908
rect 13136 5856 13142 5908
rect 14826 5856 14832 5908
rect 14884 5856 14890 5908
rect 16298 5856 16304 5908
rect 16356 5896 16362 5908
rect 16356 5868 18276 5896
rect 16356 5856 16362 5868
rect 9953 5831 10011 5837
rect 9953 5797 9965 5831
rect 9999 5797 10011 5831
rect 9953 5791 10011 5797
rect 7469 5763 7527 5769
rect 7469 5729 7481 5763
rect 7515 5760 7527 5763
rect 7650 5760 7656 5772
rect 7515 5732 7656 5760
rect 7515 5729 7527 5732
rect 7469 5723 7527 5729
rect 7650 5720 7656 5732
rect 7708 5720 7714 5772
rect 7745 5763 7803 5769
rect 7745 5729 7757 5763
rect 7791 5760 7803 5763
rect 7926 5760 7932 5772
rect 7791 5732 7932 5760
rect 7791 5729 7803 5732
rect 7745 5723 7803 5729
rect 7926 5720 7932 5732
rect 7984 5720 7990 5772
rect 9493 5763 9551 5769
rect 9493 5729 9505 5763
rect 9539 5760 9551 5763
rect 9766 5760 9772 5772
rect 9539 5732 9772 5760
rect 9539 5729 9551 5732
rect 9493 5723 9551 5729
rect 9766 5720 9772 5732
rect 9824 5720 9830 5772
rect 5902 5652 5908 5704
rect 5960 5652 5966 5704
rect 6086 5652 6092 5704
rect 6144 5652 6150 5704
rect 7377 5695 7435 5701
rect 7377 5661 7389 5695
rect 7423 5692 7435 5695
rect 7558 5692 7564 5704
rect 7423 5664 7564 5692
rect 7423 5661 7435 5664
rect 7377 5655 7435 5661
rect 7558 5652 7564 5664
rect 7616 5652 7622 5704
rect 8754 5652 8760 5704
rect 8812 5692 8818 5704
rect 9582 5692 9588 5704
rect 8812 5664 9588 5692
rect 8812 5652 8818 5664
rect 9582 5652 9588 5664
rect 9640 5652 9646 5704
rect 9968 5692 9996 5791
rect 10226 5788 10232 5840
rect 10284 5828 10290 5840
rect 10962 5828 10968 5840
rect 10284 5800 10968 5828
rect 10284 5788 10290 5800
rect 10962 5788 10968 5800
rect 11020 5828 11026 5840
rect 11057 5831 11115 5837
rect 11057 5828 11069 5831
rect 11020 5800 11069 5828
rect 11020 5788 11026 5800
rect 11057 5797 11069 5800
rect 11103 5797 11115 5831
rect 11057 5791 11115 5797
rect 11790 5788 11796 5840
rect 11848 5828 11854 5840
rect 12158 5828 12164 5840
rect 11848 5800 12164 5828
rect 11848 5788 11854 5800
rect 12158 5788 12164 5800
rect 12216 5788 12222 5840
rect 12253 5831 12311 5837
rect 12253 5797 12265 5831
rect 12299 5828 12311 5831
rect 13170 5828 13176 5840
rect 12299 5800 13176 5828
rect 12299 5797 12311 5800
rect 12253 5791 12311 5797
rect 13170 5788 13176 5800
rect 13228 5788 13234 5840
rect 16850 5788 16856 5840
rect 16908 5828 16914 5840
rect 16908 5800 17816 5828
rect 16908 5788 16914 5800
rect 12526 5720 12532 5772
rect 12584 5720 12590 5772
rect 16945 5763 17003 5769
rect 16945 5760 16957 5763
rect 16684 5732 16957 5760
rect 11882 5692 11888 5704
rect 9968 5664 11888 5692
rect 11882 5652 11888 5664
rect 11940 5692 11946 5704
rect 12069 5695 12127 5701
rect 12069 5692 12081 5695
rect 11940 5664 12081 5692
rect 11940 5652 11946 5664
rect 12069 5661 12081 5664
rect 12115 5661 12127 5695
rect 12069 5655 12127 5661
rect 12342 5652 12348 5704
rect 12400 5652 12406 5704
rect 12802 5652 12808 5704
rect 12860 5692 12866 5704
rect 13265 5695 13323 5701
rect 13265 5692 13277 5695
rect 12860 5664 13277 5692
rect 12860 5652 12866 5664
rect 13265 5661 13277 5664
rect 13311 5692 13323 5695
rect 14090 5692 14096 5704
rect 13311 5664 14096 5692
rect 13311 5661 13323 5664
rect 13265 5655 13323 5661
rect 14090 5652 14096 5664
rect 14148 5652 14154 5704
rect 14458 5652 14464 5704
rect 14516 5652 14522 5704
rect 15838 5652 15844 5704
rect 15896 5692 15902 5704
rect 16684 5701 16712 5732
rect 16945 5729 16957 5732
rect 16991 5760 17003 5763
rect 16991 5732 17632 5760
rect 16991 5729 17003 5732
rect 16945 5723 17003 5729
rect 16669 5695 16727 5701
rect 16669 5692 16681 5695
rect 15896 5664 16681 5692
rect 15896 5652 15902 5664
rect 16669 5661 16681 5664
rect 16715 5661 16727 5695
rect 16669 5655 16727 5661
rect 16850 5652 16856 5704
rect 16908 5652 16914 5704
rect 17037 5695 17095 5701
rect 17037 5661 17049 5695
rect 17083 5692 17095 5695
rect 17310 5692 17316 5704
rect 17083 5664 17316 5692
rect 17083 5661 17095 5664
rect 17037 5655 17095 5661
rect 17310 5652 17316 5664
rect 17368 5652 17374 5704
rect 17408 5695 17466 5701
rect 17408 5661 17420 5695
rect 17454 5661 17466 5695
rect 17604 5692 17632 5732
rect 17681 5695 17739 5701
rect 17681 5692 17693 5695
rect 17604 5664 17693 5692
rect 17408 5655 17466 5661
rect 17681 5661 17693 5664
rect 17727 5661 17739 5695
rect 17788 5692 17816 5800
rect 17865 5695 17923 5701
rect 17865 5692 17877 5695
rect 17788 5664 17877 5692
rect 17681 5655 17739 5661
rect 17865 5661 17877 5664
rect 17911 5661 17923 5695
rect 17865 5655 17923 5661
rect 8386 5584 8392 5636
rect 8444 5624 8450 5636
rect 9030 5624 9036 5636
rect 8444 5596 9036 5624
rect 8444 5584 8450 5596
rect 9030 5584 9036 5596
rect 9088 5624 9094 5636
rect 10781 5627 10839 5633
rect 10781 5624 10793 5627
rect 9088 5596 10793 5624
rect 9088 5584 9094 5596
rect 10781 5593 10793 5596
rect 10827 5593 10839 5627
rect 10781 5587 10839 5593
rect 12710 5584 12716 5636
rect 12768 5624 12774 5636
rect 13449 5627 13507 5633
rect 13449 5624 13461 5627
rect 12768 5596 13461 5624
rect 12768 5584 12774 5596
rect 13449 5593 13461 5596
rect 13495 5624 13507 5627
rect 14645 5627 14703 5633
rect 14645 5624 14657 5627
rect 13495 5596 14657 5624
rect 13495 5593 13507 5596
rect 13449 5587 13507 5593
rect 14645 5593 14657 5596
rect 14691 5624 14703 5627
rect 15194 5624 15200 5636
rect 14691 5596 15200 5624
rect 14691 5593 14703 5596
rect 14645 5587 14703 5593
rect 15194 5584 15200 5596
rect 15252 5584 15258 5636
rect 17420 5624 17448 5655
rect 17954 5652 17960 5704
rect 18012 5652 18018 5704
rect 18248 5701 18276 5868
rect 18414 5856 18420 5908
rect 18472 5856 18478 5908
rect 20901 5899 20959 5905
rect 20901 5865 20913 5899
rect 20947 5896 20959 5899
rect 22005 5899 22063 5905
rect 20947 5868 21404 5896
rect 20947 5865 20959 5868
rect 20901 5859 20959 5865
rect 18690 5788 18696 5840
rect 18748 5788 18754 5840
rect 18877 5831 18935 5837
rect 18877 5797 18889 5831
rect 18923 5828 18935 5831
rect 20916 5828 20944 5859
rect 21266 5828 21272 5840
rect 18923 5800 20944 5828
rect 21100 5800 21272 5828
rect 18923 5797 18935 5800
rect 18877 5791 18935 5797
rect 18708 5760 18736 5788
rect 18708 5732 19012 5760
rect 18984 5701 19012 5732
rect 20254 5720 20260 5772
rect 20312 5720 20318 5772
rect 18233 5695 18291 5701
rect 18233 5661 18245 5695
rect 18279 5692 18291 5695
rect 18693 5695 18751 5701
rect 18693 5692 18705 5695
rect 18279 5664 18705 5692
rect 18279 5661 18291 5664
rect 18233 5655 18291 5661
rect 18693 5661 18705 5664
rect 18739 5661 18751 5695
rect 18693 5655 18751 5661
rect 18969 5695 19027 5701
rect 18969 5661 18981 5695
rect 19015 5661 19027 5695
rect 18969 5655 19027 5661
rect 19797 5695 19855 5701
rect 19797 5661 19809 5695
rect 19843 5661 19855 5695
rect 19797 5655 19855 5661
rect 17773 5627 17831 5633
rect 17773 5624 17785 5627
rect 17328 5596 17448 5624
rect 17512 5596 17785 5624
rect 17328 5568 17356 5596
rect 5994 5516 6000 5568
rect 6052 5556 6058 5568
rect 6638 5556 6644 5568
rect 6052 5528 6644 5556
rect 6052 5516 6058 5528
rect 6638 5516 6644 5528
rect 6696 5516 6702 5568
rect 11882 5516 11888 5568
rect 11940 5516 11946 5568
rect 16666 5516 16672 5568
rect 16724 5556 16730 5568
rect 16761 5559 16819 5565
rect 16761 5556 16773 5559
rect 16724 5528 16773 5556
rect 16724 5516 16730 5528
rect 16761 5525 16773 5528
rect 16807 5525 16819 5559
rect 16761 5519 16819 5525
rect 17310 5516 17316 5568
rect 17368 5516 17374 5568
rect 17405 5559 17463 5565
rect 17405 5525 17417 5559
rect 17451 5556 17463 5559
rect 17512 5556 17540 5596
rect 17773 5593 17785 5596
rect 17819 5593 17831 5627
rect 18598 5624 18604 5636
rect 17773 5587 17831 5593
rect 17972 5596 18604 5624
rect 17451 5528 17540 5556
rect 17589 5559 17647 5565
rect 17451 5525 17463 5528
rect 17405 5519 17463 5525
rect 17589 5525 17601 5559
rect 17635 5556 17647 5559
rect 17972 5556 18000 5596
rect 18598 5584 18604 5596
rect 18656 5624 18662 5636
rect 18785 5627 18843 5633
rect 18785 5624 18797 5627
rect 18656 5596 18797 5624
rect 18656 5584 18662 5596
rect 18785 5593 18797 5596
rect 18831 5593 18843 5627
rect 19812 5624 19840 5655
rect 20346 5652 20352 5704
rect 20404 5652 20410 5704
rect 20456 5701 20484 5800
rect 20714 5720 20720 5772
rect 20772 5760 20778 5772
rect 21100 5769 21128 5800
rect 21266 5788 21272 5800
rect 21324 5788 21330 5840
rect 21085 5763 21143 5769
rect 20772 5732 21036 5760
rect 20772 5720 20778 5732
rect 20441 5695 20499 5701
rect 20441 5661 20453 5695
rect 20487 5661 20499 5695
rect 20441 5655 20499 5661
rect 20908 5695 20966 5701
rect 20908 5661 20920 5695
rect 20954 5661 20966 5695
rect 21008 5692 21036 5732
rect 21085 5729 21097 5763
rect 21131 5729 21143 5763
rect 21085 5723 21143 5729
rect 21269 5695 21327 5701
rect 21269 5692 21281 5695
rect 21008 5664 21281 5692
rect 20908 5655 20966 5661
rect 21269 5661 21281 5664
rect 21315 5661 21327 5695
rect 21376 5692 21404 5868
rect 22005 5865 22017 5899
rect 22051 5896 22063 5899
rect 23198 5896 23204 5908
rect 22051 5868 23204 5896
rect 22051 5865 22063 5868
rect 22005 5859 22063 5865
rect 23198 5856 23204 5868
rect 23256 5856 23262 5908
rect 25409 5899 25467 5905
rect 25409 5896 25421 5899
rect 23860 5868 25421 5896
rect 21545 5831 21603 5837
rect 21545 5797 21557 5831
rect 21591 5797 21603 5831
rect 21545 5791 21603 5797
rect 21560 5760 21588 5791
rect 22186 5788 22192 5840
rect 22244 5828 22250 5840
rect 22370 5828 22376 5840
rect 22244 5800 22376 5828
rect 22244 5788 22250 5800
rect 22370 5788 22376 5800
rect 22428 5788 22434 5840
rect 23566 5788 23572 5840
rect 23624 5828 23630 5840
rect 23860 5837 23888 5868
rect 25409 5865 25421 5868
rect 25455 5865 25467 5899
rect 25409 5859 25467 5865
rect 23845 5831 23903 5837
rect 23845 5828 23857 5831
rect 23624 5800 23857 5828
rect 23624 5788 23630 5800
rect 23845 5797 23857 5800
rect 23891 5797 23903 5831
rect 23845 5791 23903 5797
rect 23937 5831 23995 5837
rect 23937 5797 23949 5831
rect 23983 5828 23995 5831
rect 24302 5828 24308 5840
rect 23983 5800 24308 5828
rect 23983 5797 23995 5800
rect 23937 5791 23995 5797
rect 24302 5788 24308 5800
rect 24360 5788 24366 5840
rect 22278 5760 22284 5772
rect 21560 5732 21956 5760
rect 21545 5695 21603 5701
rect 21545 5692 21557 5695
rect 21376 5664 21557 5692
rect 21269 5655 21327 5661
rect 21545 5661 21557 5664
rect 21591 5661 21603 5695
rect 21545 5655 21603 5661
rect 19886 5624 19892 5636
rect 19812 5596 19892 5624
rect 18785 5587 18843 5593
rect 19886 5584 19892 5596
rect 19944 5624 19950 5636
rect 20916 5624 20944 5655
rect 21634 5652 21640 5704
rect 21692 5652 21698 5704
rect 21928 5701 21956 5732
rect 22112 5732 22284 5760
rect 22112 5701 22140 5732
rect 22278 5720 22284 5732
rect 22336 5720 22342 5772
rect 25222 5720 25228 5772
rect 25280 5760 25286 5772
rect 25501 5763 25559 5769
rect 25501 5760 25513 5763
rect 25280 5732 25513 5760
rect 25280 5720 25286 5732
rect 25501 5729 25513 5732
rect 25547 5729 25559 5763
rect 25501 5723 25559 5729
rect 21913 5695 21971 5701
rect 21913 5661 21925 5695
rect 21959 5661 21971 5695
rect 21913 5655 21971 5661
rect 22097 5695 22155 5701
rect 22097 5661 22109 5695
rect 22143 5661 22155 5695
rect 22097 5655 22155 5661
rect 19944 5596 20944 5624
rect 19944 5584 19950 5596
rect 21174 5584 21180 5636
rect 21232 5584 21238 5636
rect 21361 5627 21419 5633
rect 21361 5593 21373 5627
rect 21407 5624 21419 5627
rect 21729 5627 21787 5633
rect 21729 5624 21741 5627
rect 21407 5596 21741 5624
rect 21407 5593 21419 5596
rect 21361 5587 21419 5593
rect 21729 5593 21741 5596
rect 21775 5593 21787 5627
rect 21928 5624 21956 5655
rect 22186 5652 22192 5704
rect 22244 5652 22250 5704
rect 22373 5695 22431 5701
rect 22373 5661 22385 5695
rect 22419 5692 22431 5695
rect 22922 5692 22928 5704
rect 22419 5664 22928 5692
rect 22419 5661 22431 5664
rect 22373 5655 22431 5661
rect 22922 5652 22928 5664
rect 22980 5652 22986 5704
rect 23750 5652 23756 5704
rect 23808 5652 23814 5704
rect 24026 5652 24032 5704
rect 24084 5652 24090 5704
rect 24946 5652 24952 5704
rect 25004 5701 25010 5704
rect 25004 5695 25040 5701
rect 25028 5661 25040 5695
rect 25004 5655 25040 5661
rect 25004 5652 25010 5655
rect 22554 5624 22560 5636
rect 21928 5596 22560 5624
rect 21729 5587 21787 5593
rect 17635 5528 18000 5556
rect 17635 5525 17647 5528
rect 17589 5519 17647 5525
rect 18046 5516 18052 5568
rect 18104 5516 18110 5568
rect 20438 5516 20444 5568
rect 20496 5556 20502 5568
rect 20717 5559 20775 5565
rect 20717 5556 20729 5559
rect 20496 5528 20729 5556
rect 20496 5516 20502 5528
rect 20717 5525 20729 5528
rect 20763 5525 20775 5559
rect 20717 5519 20775 5525
rect 20898 5516 20904 5568
rect 20956 5556 20962 5568
rect 21376 5556 21404 5587
rect 22554 5584 22560 5596
rect 22612 5584 22618 5636
rect 20956 5528 21404 5556
rect 22281 5559 22339 5565
rect 20956 5516 20962 5528
rect 22281 5525 22293 5559
rect 22327 5556 22339 5559
rect 23198 5556 23204 5568
rect 22327 5528 23204 5556
rect 22327 5525 22339 5528
rect 22281 5519 22339 5525
rect 23198 5516 23204 5528
rect 23256 5516 23262 5568
rect 23474 5516 23480 5568
rect 23532 5556 23538 5568
rect 23569 5559 23627 5565
rect 23569 5556 23581 5559
rect 23532 5528 23581 5556
rect 23532 5516 23538 5528
rect 23569 5525 23581 5528
rect 23615 5525 23627 5559
rect 23569 5519 23627 5525
rect 24854 5516 24860 5568
rect 24912 5516 24918 5568
rect 25038 5516 25044 5568
rect 25096 5516 25102 5568
rect 1104 5466 27876 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 27876 5466
rect 1104 5392 27876 5414
rect 5813 5355 5871 5361
rect 5813 5321 5825 5355
rect 5859 5352 5871 5355
rect 6086 5352 6092 5364
rect 5859 5324 6092 5352
rect 5859 5321 5871 5324
rect 5813 5315 5871 5321
rect 6086 5312 6092 5324
rect 6144 5312 6150 5364
rect 6917 5355 6975 5361
rect 6917 5321 6929 5355
rect 6963 5352 6975 5355
rect 10502 5352 10508 5364
rect 6963 5324 10508 5352
rect 6963 5321 6975 5324
rect 6917 5315 6975 5321
rect 10502 5312 10508 5324
rect 10560 5352 10566 5364
rect 11790 5352 11796 5364
rect 10560 5324 11796 5352
rect 10560 5312 10566 5324
rect 11790 5312 11796 5324
rect 11848 5312 11854 5364
rect 11882 5312 11888 5364
rect 11940 5352 11946 5364
rect 12066 5352 12072 5364
rect 11940 5324 12072 5352
rect 11940 5312 11946 5324
rect 12066 5312 12072 5324
rect 12124 5312 12130 5364
rect 17681 5355 17739 5361
rect 16500 5324 17632 5352
rect 4433 5287 4491 5293
rect 4433 5253 4445 5287
rect 4479 5284 4491 5287
rect 4798 5284 4804 5296
rect 4479 5256 4804 5284
rect 4479 5253 4491 5256
rect 4433 5247 4491 5253
rect 4798 5244 4804 5256
rect 4856 5244 4862 5296
rect 13817 5287 13875 5293
rect 13817 5284 13829 5287
rect 8312 5256 9628 5284
rect 4706 5176 4712 5228
rect 4764 5216 4770 5228
rect 4985 5219 5043 5225
rect 4985 5216 4997 5219
rect 4764 5188 4997 5216
rect 4764 5176 4770 5188
rect 4985 5185 4997 5188
rect 5031 5185 5043 5219
rect 4985 5179 5043 5185
rect 5718 5176 5724 5228
rect 5776 5176 5782 5228
rect 5902 5176 5908 5228
rect 5960 5216 5966 5228
rect 5997 5219 6055 5225
rect 5997 5216 6009 5219
rect 5960 5188 6009 5216
rect 5960 5176 5966 5188
rect 5997 5185 6009 5188
rect 6043 5185 6055 5219
rect 5997 5179 6055 5185
rect 6181 5219 6239 5225
rect 6181 5185 6193 5219
rect 6227 5216 6239 5219
rect 6457 5219 6515 5225
rect 6457 5216 6469 5219
rect 6227 5188 6469 5216
rect 6227 5185 6239 5188
rect 6181 5179 6239 5185
rect 6457 5185 6469 5188
rect 6503 5185 6515 5219
rect 6457 5179 6515 5185
rect 6638 5176 6644 5228
rect 6696 5176 6702 5228
rect 6730 5176 6736 5228
rect 6788 5176 6794 5228
rect 7926 5176 7932 5228
rect 7984 5176 7990 5228
rect 8312 5225 8340 5256
rect 8205 5219 8263 5225
rect 8205 5185 8217 5219
rect 8251 5185 8263 5219
rect 8205 5179 8263 5185
rect 8297 5219 8355 5225
rect 8297 5185 8309 5219
rect 8343 5185 8355 5219
rect 8297 5179 8355 5185
rect 4724 5089 4752 5176
rect 6549 5151 6607 5157
rect 6549 5117 6561 5151
rect 6595 5148 6607 5151
rect 6822 5148 6828 5160
rect 6595 5120 6828 5148
rect 6595 5117 6607 5120
rect 6549 5111 6607 5117
rect 6822 5108 6828 5120
rect 6880 5148 6886 5160
rect 8021 5151 8079 5157
rect 8021 5148 8033 5151
rect 6880 5120 8033 5148
rect 6880 5108 6886 5120
rect 8021 5117 8033 5120
rect 8067 5117 8079 5151
rect 8220 5148 8248 5179
rect 8754 5176 8760 5228
rect 8812 5176 8818 5228
rect 9600 5225 9628 5256
rect 11992 5256 12296 5284
rect 9125 5219 9183 5225
rect 9125 5185 9137 5219
rect 9171 5185 9183 5219
rect 9125 5179 9183 5185
rect 9585 5219 9643 5225
rect 9585 5185 9597 5219
rect 9631 5216 9643 5219
rect 9766 5216 9772 5228
rect 9631 5188 9772 5216
rect 9631 5185 9643 5188
rect 9585 5179 9643 5185
rect 8665 5151 8723 5157
rect 8665 5148 8677 5151
rect 8220 5120 8677 5148
rect 8021 5111 8079 5117
rect 8665 5117 8677 5120
rect 8711 5148 8723 5151
rect 9140 5148 9168 5179
rect 9766 5176 9772 5188
rect 9824 5176 9830 5228
rect 11698 5176 11704 5228
rect 11756 5176 11762 5228
rect 11992 5225 12020 5256
rect 11977 5219 12035 5225
rect 11977 5185 11989 5219
rect 12023 5185 12035 5219
rect 11977 5179 12035 5185
rect 12066 5176 12072 5228
rect 12124 5176 12130 5228
rect 12268 5225 12296 5256
rect 13464 5256 13829 5284
rect 12253 5219 12311 5225
rect 12253 5185 12265 5219
rect 12299 5216 12311 5219
rect 12894 5216 12900 5228
rect 12299 5188 12900 5216
rect 12299 5185 12311 5188
rect 12253 5179 12311 5185
rect 12894 5176 12900 5188
rect 12952 5176 12958 5228
rect 8711 5120 9168 5148
rect 9953 5151 10011 5157
rect 8711 5117 8723 5120
rect 8665 5111 8723 5117
rect 9953 5117 9965 5151
rect 9999 5148 10011 5151
rect 9999 5120 12434 5148
rect 9999 5117 10011 5120
rect 9953 5111 10011 5117
rect 4709 5083 4767 5089
rect 4709 5049 4721 5083
rect 4755 5049 4767 5083
rect 4709 5043 4767 5049
rect 4798 5040 4804 5092
rect 4856 5080 4862 5092
rect 5261 5083 5319 5089
rect 5261 5080 5273 5083
rect 4856 5052 5273 5080
rect 4856 5040 4862 5052
rect 5261 5049 5273 5052
rect 5307 5049 5319 5083
rect 5261 5043 5319 5049
rect 11054 5040 11060 5092
rect 11112 5080 11118 5092
rect 12406 5080 12434 5120
rect 12526 5080 12532 5092
rect 11112 5052 12296 5080
rect 12406 5052 12532 5080
rect 11112 5040 11118 5052
rect 4890 4972 4896 5024
rect 4948 4972 4954 5024
rect 5442 4972 5448 5024
rect 5500 4972 5506 5024
rect 8478 4972 8484 5024
rect 8536 4972 8542 5024
rect 11514 4972 11520 5024
rect 11572 4972 11578 5024
rect 11882 4972 11888 5024
rect 11940 5012 11946 5024
rect 12161 5015 12219 5021
rect 12161 5012 12173 5015
rect 11940 4984 12173 5012
rect 11940 4972 11946 4984
rect 12161 4981 12173 4984
rect 12207 4981 12219 5015
rect 12268 5012 12296 5052
rect 12526 5040 12532 5052
rect 12584 5080 12590 5092
rect 13464 5080 13492 5256
rect 13817 5253 13829 5256
rect 13863 5284 13875 5287
rect 15933 5287 15991 5293
rect 13863 5256 15148 5284
rect 13863 5253 13875 5256
rect 13817 5247 13875 5253
rect 13722 5176 13728 5228
rect 13780 5176 13786 5228
rect 13906 5176 13912 5228
rect 13964 5216 13970 5228
rect 14001 5219 14059 5225
rect 14001 5216 14013 5219
rect 13964 5188 14013 5216
rect 13964 5176 13970 5188
rect 14001 5185 14013 5188
rect 14047 5216 14059 5219
rect 14277 5219 14335 5225
rect 14277 5216 14289 5219
rect 14047 5188 14289 5216
rect 14047 5185 14059 5188
rect 14001 5179 14059 5185
rect 14277 5185 14289 5188
rect 14323 5216 14335 5219
rect 14366 5216 14372 5228
rect 14323 5188 14372 5216
rect 14323 5185 14335 5188
rect 14277 5179 14335 5185
rect 14366 5176 14372 5188
rect 14424 5176 14430 5228
rect 15120 5225 15148 5256
rect 15933 5253 15945 5287
rect 15979 5284 15991 5287
rect 16500 5284 16528 5324
rect 17604 5284 17632 5324
rect 17681 5321 17693 5355
rect 17727 5352 17739 5355
rect 17954 5352 17960 5364
rect 17727 5324 17960 5352
rect 17727 5321 17739 5324
rect 17681 5315 17739 5321
rect 17954 5312 17960 5324
rect 18012 5352 18018 5364
rect 18012 5324 18184 5352
rect 18012 5312 18018 5324
rect 15979 5256 16528 5284
rect 15979 5253 15991 5256
rect 15933 5247 15991 5253
rect 15105 5219 15163 5225
rect 15105 5185 15117 5219
rect 15151 5185 15163 5219
rect 15105 5179 15163 5185
rect 16298 5176 16304 5228
rect 16356 5176 16362 5228
rect 16500 5225 16528 5256
rect 16684 5256 17356 5284
rect 17604 5256 17816 5284
rect 16684 5228 16712 5256
rect 16485 5219 16543 5225
rect 16485 5185 16497 5219
rect 16531 5185 16543 5219
rect 16485 5179 16543 5185
rect 16666 5176 16672 5228
rect 16724 5176 16730 5228
rect 16761 5219 16819 5225
rect 16761 5185 16773 5219
rect 16807 5185 16819 5219
rect 16761 5179 16819 5185
rect 16945 5219 17003 5225
rect 16945 5185 16957 5219
rect 16991 5185 17003 5219
rect 16945 5179 17003 5185
rect 17037 5219 17095 5225
rect 17037 5185 17049 5219
rect 17083 5216 17095 5219
rect 17218 5216 17224 5228
rect 17083 5188 17224 5216
rect 17083 5185 17095 5188
rect 17037 5179 17095 5185
rect 12584 5052 13492 5080
rect 13740 5080 13768 5176
rect 14737 5151 14795 5157
rect 14737 5117 14749 5151
rect 14783 5148 14795 5151
rect 15013 5151 15071 5157
rect 15013 5148 15025 5151
rect 14783 5120 15025 5148
rect 14783 5117 14795 5120
rect 14737 5111 14795 5117
rect 15013 5117 15025 5120
rect 15059 5117 15071 5151
rect 15013 5111 15071 5117
rect 16393 5151 16451 5157
rect 16393 5117 16405 5151
rect 16439 5148 16451 5151
rect 16776 5148 16804 5179
rect 16439 5120 16804 5148
rect 16960 5148 16988 5179
rect 17218 5176 17224 5188
rect 17276 5176 17282 5228
rect 17328 5225 17356 5256
rect 17313 5219 17371 5225
rect 17313 5185 17325 5219
rect 17359 5185 17371 5219
rect 17313 5179 17371 5185
rect 17586 5176 17592 5228
rect 17644 5216 17650 5228
rect 17681 5219 17739 5225
rect 17681 5216 17693 5219
rect 17644 5188 17693 5216
rect 17644 5176 17650 5188
rect 17681 5185 17693 5188
rect 17727 5185 17739 5219
rect 17788 5216 17816 5256
rect 17788 5214 18000 5216
rect 18046 5214 18052 5228
rect 17788 5188 18052 5214
rect 17972 5186 18052 5188
rect 17681 5179 17739 5185
rect 18046 5176 18052 5186
rect 18104 5176 18110 5228
rect 18156 5202 18184 5324
rect 18690 5312 18696 5364
rect 18748 5352 18754 5364
rect 18748 5324 18828 5352
rect 18748 5312 18754 5324
rect 18800 5293 18828 5324
rect 19886 5312 19892 5364
rect 19944 5312 19950 5364
rect 22094 5312 22100 5364
rect 22152 5352 22158 5364
rect 22152 5324 22876 5352
rect 22152 5312 22158 5324
rect 18785 5287 18843 5293
rect 18785 5253 18797 5287
rect 18831 5253 18843 5287
rect 18785 5247 18843 5253
rect 21910 5244 21916 5296
rect 21968 5284 21974 5296
rect 21968 5256 22692 5284
rect 21968 5244 21974 5256
rect 19794 5176 19800 5228
rect 19852 5176 19858 5228
rect 19978 5176 19984 5228
rect 20036 5176 20042 5228
rect 21453 5219 21511 5225
rect 21453 5185 21465 5219
rect 21499 5185 21511 5219
rect 21453 5179 21511 5185
rect 21545 5219 21603 5225
rect 21545 5185 21557 5219
rect 21591 5216 21603 5219
rect 22097 5219 22155 5225
rect 22097 5216 22109 5219
rect 21591 5188 22109 5216
rect 21591 5185 21603 5188
rect 21545 5179 21603 5185
rect 22097 5185 22109 5188
rect 22143 5216 22155 5219
rect 22370 5216 22376 5228
rect 22143 5188 22376 5216
rect 22143 5185 22155 5188
rect 22097 5179 22155 5185
rect 17236 5148 17264 5176
rect 17865 5151 17923 5157
rect 17865 5148 17877 5151
rect 16960 5120 17080 5148
rect 17236 5120 17877 5148
rect 16439 5117 16451 5120
rect 16393 5111 16451 5117
rect 16500 5092 16528 5120
rect 14553 5083 14611 5089
rect 14553 5080 14565 5083
rect 13740 5052 14565 5080
rect 12584 5040 12590 5052
rect 14553 5049 14565 5052
rect 14599 5049 14611 5083
rect 14553 5043 14611 5049
rect 16482 5040 16488 5092
rect 16540 5040 16546 5092
rect 13906 5012 13912 5024
rect 12268 4984 13912 5012
rect 12161 4975 12219 4981
rect 13906 4972 13912 4984
rect 13964 4972 13970 5024
rect 13998 4972 14004 5024
rect 14056 4972 14062 5024
rect 17052 5012 17080 5120
rect 17865 5117 17877 5120
rect 17911 5117 17923 5151
rect 19812 5148 19840 5176
rect 21468 5148 21496 5179
rect 22370 5176 22376 5188
rect 22428 5176 22434 5228
rect 22554 5176 22560 5228
rect 22612 5176 22618 5228
rect 22664 5225 22692 5256
rect 22649 5219 22707 5225
rect 22649 5185 22661 5219
rect 22695 5185 22707 5219
rect 22848 5216 22876 5324
rect 22922 5312 22928 5364
rect 22980 5312 22986 5364
rect 23661 5355 23719 5361
rect 23661 5321 23673 5355
rect 23707 5352 23719 5355
rect 24026 5352 24032 5364
rect 23707 5324 24032 5352
rect 23707 5321 23719 5324
rect 23661 5315 23719 5321
rect 24026 5312 24032 5324
rect 24084 5312 24090 5364
rect 25314 5312 25320 5364
rect 25372 5312 25378 5364
rect 23293 5219 23351 5225
rect 23293 5216 23305 5219
rect 22848 5188 23305 5216
rect 22649 5179 22707 5185
rect 23293 5185 23305 5188
rect 23339 5216 23351 5219
rect 23750 5216 23756 5228
rect 23339 5188 23756 5216
rect 23339 5185 23351 5188
rect 23293 5179 23351 5185
rect 23750 5176 23756 5188
rect 23808 5176 23814 5228
rect 24044 5216 24072 5312
rect 24673 5219 24731 5225
rect 24673 5216 24685 5219
rect 24044 5188 24685 5216
rect 24673 5185 24685 5188
rect 24719 5185 24731 5219
rect 24673 5179 24731 5185
rect 24854 5176 24860 5228
rect 24912 5176 24918 5228
rect 25130 5176 25136 5228
rect 25188 5176 25194 5228
rect 19812 5120 21496 5148
rect 22189 5151 22247 5157
rect 17865 5111 17923 5117
rect 22189 5117 22201 5151
rect 22235 5148 22247 5151
rect 22922 5148 22928 5160
rect 22235 5120 22928 5148
rect 22235 5117 22247 5120
rect 22189 5111 22247 5117
rect 22922 5108 22928 5120
rect 22980 5108 22986 5160
rect 23198 5108 23204 5160
rect 23256 5108 23262 5160
rect 17221 5083 17279 5089
rect 17221 5049 17233 5083
rect 17267 5080 17279 5083
rect 18322 5080 18328 5092
rect 17267 5052 18328 5080
rect 17267 5049 17279 5052
rect 17221 5043 17279 5049
rect 18322 5040 18328 5052
rect 18380 5040 18386 5092
rect 19978 5040 19984 5092
rect 20036 5080 20042 5092
rect 22094 5080 22100 5092
rect 20036 5052 22100 5080
rect 20036 5040 20042 5052
rect 22094 5040 22100 5052
rect 22152 5040 22158 5092
rect 22296 5052 22508 5080
rect 17586 5012 17592 5024
rect 17052 4984 17592 5012
rect 17586 4972 17592 4984
rect 17644 4972 17650 5024
rect 21818 4972 21824 5024
rect 21876 5012 21882 5024
rect 22296 5012 22324 5052
rect 21876 4984 22324 5012
rect 21876 4972 21882 4984
rect 22370 4972 22376 5024
rect 22428 4972 22434 5024
rect 22480 5012 22508 5052
rect 22557 5015 22615 5021
rect 22557 5012 22569 5015
rect 22480 4984 22569 5012
rect 22557 4981 22569 4984
rect 22603 4981 22615 5015
rect 22557 4975 22615 4981
rect 1104 4922 27876 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 27876 4922
rect 1104 4848 27876 4870
rect 7650 4768 7656 4820
rect 7708 4808 7714 4820
rect 10686 4808 10692 4820
rect 7708 4780 10692 4808
rect 7708 4768 7714 4780
rect 10686 4768 10692 4780
rect 10744 4768 10750 4820
rect 14645 4811 14703 4817
rect 14645 4777 14657 4811
rect 14691 4808 14703 4811
rect 16298 4808 16304 4820
rect 14691 4780 16304 4808
rect 14691 4777 14703 4780
rect 14645 4771 14703 4777
rect 16298 4768 16304 4780
rect 16356 4768 16362 4820
rect 18417 4811 18475 4817
rect 18417 4777 18429 4811
rect 18463 4808 18475 4811
rect 19794 4808 19800 4820
rect 18463 4780 19800 4808
rect 18463 4777 18475 4780
rect 18417 4771 18475 4777
rect 19794 4768 19800 4780
rect 19852 4768 19858 4820
rect 20438 4768 20444 4820
rect 20496 4768 20502 4820
rect 22370 4768 22376 4820
rect 22428 4808 22434 4820
rect 23566 4808 23572 4820
rect 22428 4780 23572 4808
rect 22428 4768 22434 4780
rect 23566 4768 23572 4780
rect 23624 4768 23630 4820
rect 24302 4768 24308 4820
rect 24360 4808 24366 4820
rect 24581 4811 24639 4817
rect 24581 4808 24593 4811
rect 24360 4780 24593 4808
rect 24360 4768 24366 4780
rect 24581 4777 24593 4780
rect 24627 4808 24639 4811
rect 25038 4808 25044 4820
rect 24627 4780 25044 4808
rect 24627 4777 24639 4780
rect 24581 4771 24639 4777
rect 25038 4768 25044 4780
rect 25096 4768 25102 4820
rect 6546 4700 6552 4752
rect 6604 4700 6610 4752
rect 10962 4740 10968 4752
rect 8496 4712 9168 4740
rect 4709 4675 4767 4681
rect 4709 4641 4721 4675
rect 4755 4672 4767 4675
rect 4755 4644 5488 4672
rect 4755 4641 4767 4644
rect 4709 4635 4767 4641
rect 5460 4616 5488 4644
rect 5718 4632 5724 4684
rect 5776 4672 5782 4684
rect 8496 4681 8524 4712
rect 9140 4681 9168 4712
rect 9232 4712 10968 4740
rect 9232 4681 9260 4712
rect 10962 4700 10968 4712
rect 11020 4740 11026 4752
rect 11020 4712 13400 4740
rect 11020 4700 11026 4712
rect 6089 4675 6147 4681
rect 6089 4672 6101 4675
rect 5776 4644 6101 4672
rect 5776 4632 5782 4644
rect 6089 4641 6101 4644
rect 6135 4641 6147 4675
rect 8481 4675 8539 4681
rect 6089 4635 6147 4641
rect 7484 4644 8432 4672
rect 7484 4616 7512 4644
rect 4614 4564 4620 4616
rect 4672 4604 4678 4616
rect 4801 4607 4859 4613
rect 4801 4604 4813 4607
rect 4672 4576 4813 4604
rect 4672 4564 4678 4576
rect 4801 4573 4813 4576
rect 4847 4573 4859 4607
rect 4801 4567 4859 4573
rect 4890 4564 4896 4616
rect 4948 4604 4954 4616
rect 5261 4607 5319 4613
rect 5261 4604 5273 4607
rect 4948 4576 5273 4604
rect 4948 4564 4954 4576
rect 5261 4573 5273 4576
rect 5307 4573 5319 4607
rect 5261 4567 5319 4573
rect 5442 4564 5448 4616
rect 5500 4564 5506 4616
rect 6178 4564 6184 4616
rect 6236 4564 6242 4616
rect 7466 4564 7472 4616
rect 7524 4564 7530 4616
rect 8404 4604 8432 4644
rect 8481 4641 8493 4675
rect 8527 4641 8539 4675
rect 8481 4635 8539 4641
rect 8665 4675 8723 4681
rect 8665 4641 8677 4675
rect 8711 4672 8723 4675
rect 9033 4675 9091 4681
rect 9033 4672 9045 4675
rect 8711 4644 9045 4672
rect 8711 4641 8723 4644
rect 8665 4635 8723 4641
rect 9033 4641 9045 4644
rect 9079 4641 9091 4675
rect 9033 4635 9091 4641
rect 9125 4675 9183 4681
rect 9125 4641 9137 4675
rect 9171 4641 9183 4675
rect 9125 4635 9183 4641
rect 9217 4675 9275 4681
rect 9217 4641 9229 4675
rect 9263 4641 9275 4675
rect 9217 4635 9275 4641
rect 9309 4675 9367 4681
rect 9309 4641 9321 4675
rect 9355 4672 9367 4675
rect 9355 4644 9536 4672
rect 9355 4641 9367 4644
rect 9309 4635 9367 4641
rect 8573 4607 8631 4613
rect 8573 4604 8585 4607
rect 5629 4539 5687 4545
rect 5629 4505 5641 4539
rect 5675 4536 5687 4539
rect 7650 4536 7656 4548
rect 5675 4508 7656 4536
rect 5675 4505 5687 4508
rect 5629 4499 5687 4505
rect 7650 4496 7656 4508
rect 7708 4496 7714 4548
rect 8128 4536 8156 4590
rect 8404 4576 8585 4604
rect 8573 4573 8585 4576
rect 8619 4573 8631 4607
rect 8573 4567 8631 4573
rect 8757 4607 8815 4613
rect 8757 4573 8769 4607
rect 8803 4573 8815 4607
rect 8757 4567 8815 4573
rect 8478 4536 8484 4548
rect 8128 4508 8484 4536
rect 8478 4496 8484 4508
rect 8536 4536 8542 4548
rect 8772 4536 8800 4567
rect 8536 4508 8800 4536
rect 9140 4536 9168 4635
rect 9508 4604 9536 4644
rect 9582 4632 9588 4684
rect 9640 4672 9646 4684
rect 12342 4672 12348 4684
rect 9640 4644 12348 4672
rect 9640 4632 9646 4644
rect 12342 4632 12348 4644
rect 12400 4672 12406 4684
rect 13372 4681 13400 4712
rect 21910 4700 21916 4752
rect 21968 4740 21974 4752
rect 22097 4743 22155 4749
rect 22097 4740 22109 4743
rect 21968 4712 22109 4740
rect 21968 4700 21974 4712
rect 22097 4709 22109 4712
rect 22143 4709 22155 4743
rect 22097 4703 22155 4709
rect 25317 4743 25375 4749
rect 25317 4709 25329 4743
rect 25363 4740 25375 4743
rect 25498 4740 25504 4752
rect 25363 4712 25504 4740
rect 25363 4709 25375 4712
rect 25317 4703 25375 4709
rect 25498 4700 25504 4712
rect 25556 4700 25562 4752
rect 12621 4675 12679 4681
rect 12400 4632 12434 4672
rect 12621 4641 12633 4675
rect 12667 4672 12679 4675
rect 12989 4675 13047 4681
rect 12989 4672 13001 4675
rect 12667 4644 13001 4672
rect 12667 4641 12679 4644
rect 12621 4635 12679 4641
rect 12989 4641 13001 4644
rect 13035 4641 13047 4675
rect 12989 4635 13047 4641
rect 13357 4675 13415 4681
rect 13357 4641 13369 4675
rect 13403 4672 13415 4675
rect 14369 4675 14427 4681
rect 13403 4644 14320 4672
rect 13403 4641 13415 4644
rect 13357 4635 13415 4641
rect 9508 4576 10456 4604
rect 9582 4536 9588 4548
rect 9140 4508 9588 4536
rect 8536 4496 8542 4508
rect 9582 4496 9588 4508
rect 9640 4496 9646 4548
rect 10428 4536 10456 4576
rect 10502 4564 10508 4616
rect 10560 4564 10566 4616
rect 10686 4564 10692 4616
rect 10744 4564 10750 4616
rect 12406 4604 12434 4632
rect 14292 4613 14320 4644
rect 14369 4641 14381 4675
rect 14415 4641 14427 4675
rect 16393 4675 16451 4681
rect 16393 4672 16405 4675
rect 14369 4635 14427 4641
rect 15672 4644 16405 4672
rect 12529 4607 12587 4613
rect 12529 4604 12541 4607
rect 12406 4576 12541 4604
rect 12529 4573 12541 4576
rect 12575 4573 12587 4607
rect 12529 4567 12587 4573
rect 13173 4607 13231 4613
rect 13173 4573 13185 4607
rect 13219 4573 13231 4607
rect 13173 4567 13231 4573
rect 14277 4607 14335 4613
rect 14277 4573 14289 4607
rect 14323 4573 14335 4607
rect 14277 4567 14335 4573
rect 13188 4536 13216 4567
rect 13998 4536 14004 4548
rect 10428 4508 14004 4536
rect 13998 4496 14004 4508
rect 14056 4536 14062 4548
rect 14384 4536 14412 4635
rect 15672 4616 15700 4644
rect 16393 4641 16405 4644
rect 16439 4641 16451 4675
rect 16393 4635 16451 4641
rect 18233 4675 18291 4681
rect 18233 4641 18245 4675
rect 18279 4672 18291 4675
rect 18322 4672 18328 4684
rect 18279 4644 18328 4672
rect 18279 4641 18291 4644
rect 18233 4635 18291 4641
rect 18322 4632 18328 4644
rect 18380 4632 18386 4684
rect 20530 4632 20536 4684
rect 20588 4632 20594 4684
rect 25041 4675 25099 4681
rect 25041 4641 25053 4675
rect 25087 4672 25099 4675
rect 25130 4672 25136 4684
rect 25087 4644 25136 4672
rect 25087 4641 25099 4644
rect 25041 4635 25099 4641
rect 25130 4632 25136 4644
rect 25188 4632 25194 4684
rect 15562 4564 15568 4616
rect 15620 4564 15626 4616
rect 15654 4564 15660 4616
rect 15712 4564 15718 4616
rect 16301 4607 16359 4613
rect 16301 4604 16313 4607
rect 15764 4576 16313 4604
rect 14056 4508 14412 4536
rect 14056 4496 14062 4508
rect 5169 4471 5227 4477
rect 5169 4437 5181 4471
rect 5215 4468 5227 4471
rect 8018 4468 8024 4480
rect 5215 4440 8024 4468
rect 5215 4437 5227 4440
rect 5169 4431 5227 4437
rect 8018 4428 8024 4440
rect 8076 4428 8082 4480
rect 9490 4428 9496 4480
rect 9548 4428 9554 4480
rect 10597 4471 10655 4477
rect 10597 4437 10609 4471
rect 10643 4468 10655 4471
rect 11146 4468 11152 4480
rect 10643 4440 11152 4468
rect 10643 4437 10655 4440
rect 10597 4431 10655 4437
rect 11146 4428 11152 4440
rect 11204 4428 11210 4480
rect 11514 4428 11520 4480
rect 11572 4468 11578 4480
rect 12802 4468 12808 4480
rect 11572 4440 12808 4468
rect 11572 4428 11578 4440
rect 12802 4428 12808 4440
rect 12860 4428 12866 4480
rect 12897 4471 12955 4477
rect 12897 4437 12909 4471
rect 12943 4468 12955 4471
rect 15764 4468 15792 4576
rect 16301 4573 16313 4576
rect 16347 4573 16359 4607
rect 16301 4567 16359 4573
rect 16316 4536 16344 4567
rect 16482 4564 16488 4616
rect 16540 4564 16546 4616
rect 18141 4607 18199 4613
rect 18141 4573 18153 4607
rect 18187 4573 18199 4607
rect 18141 4567 18199 4573
rect 18156 4536 18184 4567
rect 20070 4564 20076 4616
rect 20128 4564 20134 4616
rect 20254 4564 20260 4616
rect 20312 4564 20318 4616
rect 21726 4564 21732 4616
rect 21784 4604 21790 4616
rect 21913 4607 21971 4613
rect 21913 4604 21925 4607
rect 21784 4576 21925 4604
rect 21784 4564 21790 4576
rect 21913 4573 21925 4576
rect 21959 4573 21971 4607
rect 22281 4607 22339 4613
rect 22281 4604 22293 4607
rect 21913 4567 21971 4573
rect 22066 4576 22293 4604
rect 16316 4508 18184 4536
rect 20088 4536 20116 4564
rect 22066 4536 22094 4576
rect 22281 4573 22293 4576
rect 22327 4573 22339 4607
rect 22281 4567 22339 4573
rect 24394 4564 24400 4616
rect 24452 4564 24458 4616
rect 24670 4564 24676 4616
rect 24728 4604 24734 4616
rect 24949 4607 25007 4613
rect 24949 4604 24961 4607
rect 24728 4576 24961 4604
rect 24728 4564 24734 4576
rect 24949 4573 24961 4576
rect 24995 4573 25007 4607
rect 24949 4567 25007 4573
rect 20088 4508 22094 4536
rect 12943 4440 15792 4468
rect 15841 4471 15899 4477
rect 12943 4437 12955 4440
rect 12897 4431 12955 4437
rect 15841 4437 15853 4471
rect 15887 4468 15899 4471
rect 16206 4468 16212 4480
rect 15887 4440 16212 4468
rect 15887 4437 15899 4440
rect 15841 4431 15899 4437
rect 16206 4428 16212 4440
rect 16264 4428 16270 4480
rect 20073 4471 20131 4477
rect 20073 4437 20085 4471
rect 20119 4468 20131 4471
rect 20622 4468 20628 4480
rect 20119 4440 20628 4468
rect 20119 4437 20131 4440
rect 20073 4431 20131 4437
rect 20622 4428 20628 4440
rect 20680 4428 20686 4480
rect 21634 4428 21640 4480
rect 21692 4468 21698 4480
rect 21818 4468 21824 4480
rect 21692 4440 21824 4468
rect 21692 4428 21698 4440
rect 21818 4428 21824 4440
rect 21876 4468 21882 4480
rect 22373 4471 22431 4477
rect 22373 4468 22385 4471
rect 21876 4440 22385 4468
rect 21876 4428 21882 4440
rect 22373 4437 22385 4440
rect 22419 4437 22431 4471
rect 22373 4431 22431 4437
rect 1104 4378 27876 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 27876 4378
rect 1104 4304 27876 4326
rect 6546 4224 6552 4276
rect 6604 4264 6610 4276
rect 6604 4236 9812 4264
rect 6604 4224 6610 4236
rect 8018 4156 8024 4208
rect 8076 4196 8082 4208
rect 9784 4196 9812 4236
rect 9950 4224 9956 4276
rect 10008 4264 10014 4276
rect 11517 4267 11575 4273
rect 10008 4236 11100 4264
rect 10008 4224 10014 4236
rect 10226 4196 10232 4208
rect 8076 4168 9720 4196
rect 8076 4156 8082 4168
rect 9692 4060 9720 4168
rect 9784 4168 10232 4196
rect 9784 4137 9812 4168
rect 10226 4156 10232 4168
rect 10284 4196 10290 4208
rect 10284 4168 11008 4196
rect 10284 4156 10290 4168
rect 9769 4131 9827 4137
rect 9769 4097 9781 4131
rect 9815 4097 9827 4131
rect 9769 4091 9827 4097
rect 9950 4088 9956 4140
rect 10008 4088 10014 4140
rect 10045 4131 10103 4137
rect 10045 4097 10057 4131
rect 10091 4097 10103 4131
rect 10045 4091 10103 4097
rect 10413 4131 10471 4137
rect 10413 4097 10425 4131
rect 10459 4128 10471 4131
rect 10778 4128 10784 4140
rect 10459 4100 10784 4128
rect 10459 4097 10471 4100
rect 10413 4091 10471 4097
rect 10060 4060 10088 4091
rect 10778 4088 10784 4100
rect 10836 4088 10842 4140
rect 10870 4088 10876 4140
rect 10928 4088 10934 4140
rect 10980 4137 11008 4168
rect 11072 4137 11100 4236
rect 11517 4233 11529 4267
rect 11563 4264 11575 4267
rect 11698 4264 11704 4276
rect 11563 4236 11704 4264
rect 11563 4233 11575 4236
rect 11517 4227 11575 4233
rect 11698 4224 11704 4236
rect 11756 4224 11762 4276
rect 12802 4224 12808 4276
rect 12860 4264 12866 4276
rect 13446 4264 13452 4276
rect 12860 4236 13452 4264
rect 12860 4224 12866 4236
rect 13446 4224 13452 4236
rect 13504 4264 13510 4276
rect 14550 4264 14556 4276
rect 13504 4236 14556 4264
rect 13504 4224 13510 4236
rect 14550 4224 14556 4236
rect 14608 4224 14614 4276
rect 19794 4224 19800 4276
rect 19852 4264 19858 4276
rect 20070 4264 20076 4276
rect 19852 4236 20076 4264
rect 19852 4224 19858 4236
rect 20070 4224 20076 4236
rect 20128 4224 20134 4276
rect 20346 4224 20352 4276
rect 20404 4264 20410 4276
rect 20530 4264 20536 4276
rect 20404 4236 20536 4264
rect 20404 4224 20410 4236
rect 20530 4224 20536 4236
rect 20588 4264 20594 4276
rect 24949 4267 25007 4273
rect 20588 4236 20944 4264
rect 20588 4224 20594 4236
rect 11606 4156 11612 4208
rect 11664 4196 11670 4208
rect 12161 4199 12219 4205
rect 12161 4196 12173 4199
rect 11664 4168 12173 4196
rect 11664 4156 11670 4168
rect 12161 4165 12173 4168
rect 12207 4165 12219 4199
rect 12161 4159 12219 4165
rect 15749 4199 15807 4205
rect 15749 4165 15761 4199
rect 15795 4196 15807 4199
rect 15933 4199 15991 4205
rect 15933 4196 15945 4199
rect 15795 4168 15945 4196
rect 15795 4165 15807 4168
rect 15749 4159 15807 4165
rect 15933 4165 15945 4168
rect 15979 4196 15991 4199
rect 17770 4196 17776 4208
rect 15979 4168 17776 4196
rect 15979 4165 15991 4168
rect 15933 4159 15991 4165
rect 17770 4156 17776 4168
rect 17828 4156 17834 4208
rect 20438 4156 20444 4208
rect 20496 4196 20502 4208
rect 20916 4196 20944 4236
rect 24504 4236 24808 4264
rect 24504 4205 24532 4236
rect 24489 4199 24547 4205
rect 20496 4168 20668 4196
rect 20916 4168 21128 4196
rect 20496 4156 20502 4168
rect 10965 4131 11023 4137
rect 10965 4097 10977 4131
rect 11011 4097 11023 4131
rect 10965 4091 11023 4097
rect 11057 4131 11115 4137
rect 11057 4097 11069 4131
rect 11103 4097 11115 4131
rect 11057 4091 11115 4097
rect 11146 4088 11152 4140
rect 11204 4088 11210 4140
rect 11701 4131 11759 4137
rect 11701 4097 11713 4131
rect 11747 4097 11759 4131
rect 13262 4128 13268 4140
rect 11701 4091 11759 4097
rect 12406 4100 13268 4128
rect 10597 4063 10655 4069
rect 9692 4032 10548 4060
rect 10410 3952 10416 4004
rect 10468 3952 10474 4004
rect 10520 3992 10548 4032
rect 10597 4029 10609 4063
rect 10643 4060 10655 4063
rect 10689 4063 10747 4069
rect 10689 4060 10701 4063
rect 10643 4032 10701 4060
rect 10643 4029 10655 4032
rect 10597 4023 10655 4029
rect 10689 4029 10701 4032
rect 10735 4029 10747 4063
rect 11422 4060 11428 4072
rect 10689 4023 10747 4029
rect 10980 4032 11428 4060
rect 10980 3992 11008 4032
rect 11422 4020 11428 4032
rect 11480 4060 11486 4072
rect 11716 4060 11744 4091
rect 11480 4032 11744 4060
rect 11793 4063 11851 4069
rect 11480 4020 11486 4032
rect 11793 4029 11805 4063
rect 11839 4060 11851 4063
rect 12406 4060 12434 4100
rect 13262 4088 13268 4100
rect 13320 4088 13326 4140
rect 14829 4131 14887 4137
rect 14829 4097 14841 4131
rect 14875 4097 14887 4131
rect 14829 4091 14887 4097
rect 11839 4032 12434 4060
rect 14844 4060 14872 4091
rect 15194 4088 15200 4140
rect 15252 4088 15258 4140
rect 15286 4088 15292 4140
rect 15344 4088 15350 4140
rect 15470 4088 15476 4140
rect 15528 4088 15534 4140
rect 15565 4131 15623 4137
rect 15565 4097 15577 4131
rect 15611 4128 15623 4131
rect 15654 4128 15660 4140
rect 15611 4100 15660 4128
rect 15611 4097 15623 4100
rect 15565 4091 15623 4097
rect 15654 4088 15660 4100
rect 15712 4088 15718 4140
rect 16301 4131 16359 4137
rect 16301 4097 16313 4131
rect 16347 4128 16359 4131
rect 17129 4131 17187 4137
rect 17129 4128 17141 4131
rect 16347 4100 17141 4128
rect 16347 4097 16359 4100
rect 16301 4091 16359 4097
rect 17129 4097 17141 4100
rect 17175 4128 17187 4131
rect 17218 4128 17224 4140
rect 17175 4100 17224 4128
rect 17175 4097 17187 4100
rect 17129 4091 17187 4097
rect 17218 4088 17224 4100
rect 17276 4088 17282 4140
rect 17313 4131 17371 4137
rect 17313 4097 17325 4131
rect 17359 4128 17371 4131
rect 17586 4128 17592 4140
rect 17359 4100 17592 4128
rect 17359 4097 17371 4100
rect 17313 4091 17371 4097
rect 15378 4060 15384 4072
rect 14844 4032 15384 4060
rect 11839 4029 11851 4032
rect 11793 4023 11851 4029
rect 11808 3992 11836 4023
rect 15378 4020 15384 4032
rect 15436 4020 15442 4072
rect 16574 4020 16580 4072
rect 16632 4060 16638 4072
rect 17328 4060 17356 4091
rect 17586 4088 17592 4100
rect 17644 4088 17650 4140
rect 19702 4088 19708 4140
rect 19760 4128 19766 4140
rect 19797 4131 19855 4137
rect 19797 4128 19809 4131
rect 19760 4100 19809 4128
rect 19760 4088 19766 4100
rect 19797 4097 19809 4100
rect 19843 4097 19855 4131
rect 19797 4091 19855 4097
rect 20070 4088 20076 4140
rect 20128 4088 20134 4140
rect 20254 4088 20260 4140
rect 20312 4088 20318 4140
rect 20530 4088 20536 4140
rect 20588 4088 20594 4140
rect 20640 4128 20668 4168
rect 20993 4131 21051 4137
rect 20993 4128 21005 4131
rect 20640 4100 21005 4128
rect 20993 4097 21005 4100
rect 21039 4097 21051 4131
rect 21100 4128 21128 4168
rect 24489 4165 24501 4199
rect 24535 4165 24547 4199
rect 24489 4159 24547 4165
rect 21361 4131 21419 4137
rect 21361 4128 21373 4131
rect 21100 4100 21373 4128
rect 20993 4091 21051 4097
rect 21361 4097 21373 4100
rect 21407 4097 21419 4131
rect 21361 4091 21419 4097
rect 22278 4088 22284 4140
rect 22336 4088 22342 4140
rect 22370 4088 22376 4140
rect 22428 4128 22434 4140
rect 22741 4131 22799 4137
rect 22741 4128 22753 4131
rect 22428 4100 22753 4128
rect 22428 4088 22434 4100
rect 22741 4097 22753 4100
rect 22787 4097 22799 4131
rect 22741 4091 22799 4097
rect 23198 4088 23204 4140
rect 23256 4088 23262 4140
rect 23385 4131 23443 4137
rect 23385 4097 23397 4131
rect 23431 4097 23443 4131
rect 23385 4091 23443 4097
rect 16632 4032 17356 4060
rect 16632 4020 16638 4032
rect 21818 4020 21824 4072
rect 21876 4020 21882 4072
rect 22189 4063 22247 4069
rect 22189 4060 22201 4063
rect 22066 4032 22201 4060
rect 10520 3964 11008 3992
rect 11716 3964 11836 3992
rect 15396 3992 15424 4020
rect 17678 3992 17684 4004
rect 15396 3964 17684 3992
rect 9953 3927 10011 3933
rect 9953 3893 9965 3927
rect 9999 3924 10011 3927
rect 10502 3924 10508 3936
rect 9999 3896 10508 3924
rect 9999 3893 10011 3896
rect 9953 3887 10011 3893
rect 10502 3884 10508 3896
rect 10560 3884 10566 3936
rect 10686 3884 10692 3936
rect 10744 3924 10750 3936
rect 11716 3924 11744 3964
rect 17678 3952 17684 3964
rect 17736 3952 17742 4004
rect 20622 3952 20628 4004
rect 20680 3992 20686 4004
rect 21450 3992 21456 4004
rect 20680 3964 21456 3992
rect 20680 3952 20686 3964
rect 21450 3952 21456 3964
rect 21508 3992 21514 4004
rect 22066 3992 22094 4032
rect 22189 4029 22201 4032
rect 22235 4029 22247 4063
rect 22189 4023 22247 4029
rect 22465 4063 22523 4069
rect 22465 4029 22477 4063
rect 22511 4060 22523 4063
rect 22557 4063 22615 4069
rect 22557 4060 22569 4063
rect 22511 4032 22569 4060
rect 22511 4029 22523 4032
rect 22465 4023 22523 4029
rect 22557 4029 22569 4032
rect 22603 4029 22615 4063
rect 23400 4060 23428 4091
rect 23474 4088 23480 4140
rect 23532 4128 23538 4140
rect 23845 4131 23903 4137
rect 23845 4128 23857 4131
rect 23532 4100 23857 4128
rect 23532 4088 23538 4100
rect 23845 4097 23857 4100
rect 23891 4097 23903 4131
rect 23845 4091 23903 4097
rect 24302 4088 24308 4140
rect 24360 4088 24366 4140
rect 24581 4131 24639 4137
rect 24581 4097 24593 4131
rect 24627 4097 24639 4131
rect 24581 4091 24639 4097
rect 23658 4060 23664 4072
rect 23400 4032 23664 4060
rect 22557 4023 22615 4029
rect 23658 4020 23664 4032
rect 23716 4020 23722 4072
rect 24029 4063 24087 4069
rect 24029 4029 24041 4063
rect 24075 4060 24087 4063
rect 24596 4060 24624 4091
rect 24670 4088 24676 4140
rect 24728 4088 24734 4140
rect 24780 4128 24808 4236
rect 24949 4233 24961 4267
rect 24995 4264 25007 4267
rect 25130 4264 25136 4276
rect 24995 4236 25136 4264
rect 24995 4233 25007 4236
rect 24949 4227 25007 4233
rect 25130 4224 25136 4236
rect 25188 4224 25194 4276
rect 24946 4128 24952 4140
rect 24780 4100 24952 4128
rect 24946 4088 24952 4100
rect 25004 4128 25010 4140
rect 25409 4131 25467 4137
rect 25409 4128 25421 4131
rect 25004 4100 25421 4128
rect 25004 4088 25010 4100
rect 25409 4097 25421 4100
rect 25455 4097 25467 4131
rect 25409 4091 25467 4097
rect 24075 4032 25084 4060
rect 24075 4029 24087 4032
rect 24029 4023 24087 4029
rect 21508 3964 22094 3992
rect 22925 3995 22983 4001
rect 21508 3952 21514 3964
rect 22925 3961 22937 3995
rect 22971 3992 22983 3995
rect 23474 3992 23480 4004
rect 22971 3964 23480 3992
rect 22971 3961 22983 3964
rect 22925 3955 22983 3961
rect 23474 3952 23480 3964
rect 23532 3952 23538 4004
rect 25056 4001 25084 4032
rect 25041 3995 25099 4001
rect 25041 3961 25053 3995
rect 25087 3961 25099 3995
rect 25424 3992 25452 4091
rect 25498 4088 25504 4140
rect 25556 4088 25562 4140
rect 25685 3995 25743 4001
rect 25685 3992 25697 3995
rect 25424 3964 25697 3992
rect 25041 3955 25099 3961
rect 25685 3961 25697 3964
rect 25731 3961 25743 3995
rect 25685 3955 25743 3961
rect 10744 3896 11744 3924
rect 10744 3884 10750 3896
rect 11790 3884 11796 3936
rect 11848 3884 11854 3936
rect 15013 3927 15071 3933
rect 15013 3893 15025 3927
rect 15059 3924 15071 3927
rect 16574 3924 16580 3936
rect 15059 3896 16580 3924
rect 15059 3893 15071 3896
rect 15013 3887 15071 3893
rect 16574 3884 16580 3896
rect 16632 3884 16638 3936
rect 16942 3884 16948 3936
rect 17000 3884 17006 3936
rect 23017 3927 23075 3933
rect 23017 3893 23029 3927
rect 23063 3924 23075 3927
rect 24394 3924 24400 3936
rect 23063 3896 24400 3924
rect 23063 3893 23075 3896
rect 23017 3887 23075 3893
rect 24394 3884 24400 3896
rect 24452 3884 24458 3936
rect 24854 3884 24860 3936
rect 24912 3884 24918 3936
rect 1104 3834 27876 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 27876 3834
rect 1104 3760 27876 3782
rect 10134 3680 10140 3732
rect 10192 3720 10198 3732
rect 10192 3692 16160 3720
rect 10192 3680 10198 3692
rect 13909 3655 13967 3661
rect 13909 3621 13921 3655
rect 13955 3652 13967 3655
rect 15194 3652 15200 3664
rect 13955 3624 15200 3652
rect 13955 3621 13967 3624
rect 13909 3615 13967 3621
rect 15194 3612 15200 3624
rect 15252 3612 15258 3664
rect 15378 3612 15384 3664
rect 15436 3652 15442 3664
rect 15657 3655 15715 3661
rect 15657 3652 15669 3655
rect 15436 3624 15669 3652
rect 15436 3612 15442 3624
rect 15657 3621 15669 3624
rect 15703 3621 15715 3655
rect 15657 3615 15715 3621
rect 10410 3544 10416 3596
rect 10468 3584 10474 3596
rect 10468 3556 14136 3584
rect 10468 3544 10474 3556
rect 9030 3476 9036 3528
rect 9088 3476 9094 3528
rect 9490 3476 9496 3528
rect 9548 3476 9554 3528
rect 11238 3476 11244 3528
rect 11296 3476 11302 3528
rect 11422 3476 11428 3528
rect 11480 3476 11486 3528
rect 11882 3476 11888 3528
rect 11940 3476 11946 3528
rect 13446 3516 13452 3528
rect 12406 3488 13452 3516
rect 10045 3451 10103 3457
rect 10045 3417 10057 3451
rect 10091 3448 10103 3451
rect 11146 3448 11152 3460
rect 10091 3420 11152 3448
rect 10091 3417 10103 3420
rect 10045 3411 10103 3417
rect 11146 3408 11152 3420
rect 11204 3408 11210 3460
rect 11609 3451 11667 3457
rect 11609 3417 11621 3451
rect 11655 3448 11667 3451
rect 12406 3448 12434 3488
rect 13446 3476 13452 3488
rect 13504 3476 13510 3528
rect 13538 3476 13544 3528
rect 13596 3476 13602 3528
rect 14108 3525 14136 3556
rect 16022 3544 16028 3596
rect 16080 3584 16086 3596
rect 16132 3584 16160 3692
rect 16298 3680 16304 3732
rect 16356 3720 16362 3732
rect 18874 3720 18880 3732
rect 16356 3692 18880 3720
rect 16356 3680 16362 3692
rect 18874 3680 18880 3692
rect 18932 3680 18938 3732
rect 19794 3680 19800 3732
rect 19852 3680 19858 3732
rect 20438 3680 20444 3732
rect 20496 3680 20502 3732
rect 21910 3680 21916 3732
rect 21968 3680 21974 3732
rect 23198 3680 23204 3732
rect 23256 3720 23262 3732
rect 23477 3723 23535 3729
rect 23477 3720 23489 3723
rect 23256 3692 23489 3720
rect 23256 3680 23262 3692
rect 23477 3689 23489 3692
rect 23523 3689 23535 3723
rect 23477 3683 23535 3689
rect 23845 3723 23903 3729
rect 23845 3689 23857 3723
rect 23891 3720 23903 3723
rect 25498 3720 25504 3732
rect 23891 3692 25504 3720
rect 23891 3689 23903 3692
rect 23845 3683 23903 3689
rect 25498 3680 25504 3692
rect 25556 3680 25562 3732
rect 16206 3612 16212 3664
rect 16264 3652 16270 3664
rect 17681 3655 17739 3661
rect 16264 3624 17080 3652
rect 16264 3612 16270 3624
rect 16669 3587 16727 3593
rect 16080 3556 16528 3584
rect 16080 3544 16086 3556
rect 13634 3519 13692 3525
rect 13634 3485 13646 3519
rect 13680 3485 13692 3519
rect 13634 3479 13692 3485
rect 14093 3519 14151 3525
rect 14093 3485 14105 3519
rect 14139 3485 14151 3519
rect 14093 3479 14151 3485
rect 11655 3420 12434 3448
rect 11655 3417 11667 3420
rect 11609 3411 11667 3417
rect 13262 3408 13268 3460
rect 13320 3448 13326 3460
rect 13648 3448 13676 3479
rect 14550 3476 14556 3528
rect 14608 3476 14614 3528
rect 15013 3519 15071 3525
rect 15013 3485 15025 3519
rect 15059 3485 15071 3519
rect 15013 3479 15071 3485
rect 15381 3519 15439 3525
rect 15381 3485 15393 3519
rect 15427 3485 15439 3519
rect 15381 3479 15439 3485
rect 13320 3420 13676 3448
rect 13320 3408 13326 3420
rect 13722 3408 13728 3460
rect 13780 3448 13786 3460
rect 15028 3448 15056 3479
rect 13780 3420 15056 3448
rect 13780 3408 13786 3420
rect 10870 3340 10876 3392
rect 10928 3380 10934 3392
rect 11793 3383 11851 3389
rect 11793 3380 11805 3383
rect 10928 3352 11805 3380
rect 10928 3340 10934 3352
rect 11793 3349 11805 3352
rect 11839 3349 11851 3383
rect 11793 3343 11851 3349
rect 13538 3340 13544 3392
rect 13596 3380 13602 3392
rect 15396 3380 15424 3479
rect 15654 3476 15660 3528
rect 15712 3516 15718 3528
rect 15749 3519 15807 3525
rect 15749 3516 15761 3519
rect 15712 3488 15761 3516
rect 15712 3476 15718 3488
rect 15749 3485 15761 3488
rect 15795 3516 15807 3519
rect 16298 3516 16304 3528
rect 15795 3488 16304 3516
rect 15795 3485 15807 3488
rect 15749 3479 15807 3485
rect 16298 3476 16304 3488
rect 16356 3476 16362 3528
rect 16390 3476 16396 3528
rect 16448 3476 16454 3528
rect 16500 3525 16528 3556
rect 16669 3553 16681 3587
rect 16715 3584 16727 3587
rect 16942 3584 16948 3596
rect 16715 3556 16948 3584
rect 16715 3553 16727 3556
rect 16669 3547 16727 3553
rect 16942 3544 16948 3556
rect 17000 3544 17006 3596
rect 16485 3519 16543 3525
rect 16485 3485 16497 3519
rect 16531 3485 16543 3519
rect 16485 3479 16543 3485
rect 16574 3476 16580 3528
rect 16632 3516 16638 3528
rect 17052 3525 17080 3624
rect 17681 3621 17693 3655
rect 17727 3621 17739 3655
rect 17681 3615 17739 3621
rect 18509 3655 18567 3661
rect 18509 3621 18521 3655
rect 18555 3652 18567 3655
rect 21266 3652 21272 3664
rect 18555 3624 21272 3652
rect 18555 3621 18567 3624
rect 18509 3615 18567 3621
rect 17696 3584 17724 3615
rect 21266 3612 21272 3624
rect 21324 3652 21330 3664
rect 22097 3655 22155 3661
rect 21324 3624 22048 3652
rect 21324 3612 21330 3624
rect 17144 3556 17724 3584
rect 17865 3587 17923 3593
rect 16761 3519 16819 3525
rect 16761 3516 16773 3519
rect 16632 3488 16773 3516
rect 16632 3476 16638 3488
rect 16761 3485 16773 3488
rect 16807 3516 16819 3519
rect 17037 3519 17095 3525
rect 16807 3488 16988 3516
rect 16807 3485 16819 3488
rect 16761 3479 16819 3485
rect 15562 3408 15568 3460
rect 15620 3448 15626 3460
rect 16853 3451 16911 3457
rect 16853 3448 16865 3451
rect 15620 3420 16865 3448
rect 15620 3408 15626 3420
rect 16853 3417 16865 3420
rect 16899 3417 16911 3451
rect 16960 3448 16988 3488
rect 17037 3485 17049 3519
rect 17083 3485 17095 3519
rect 17037 3479 17095 3485
rect 17144 3448 17172 3556
rect 17865 3553 17877 3587
rect 17911 3584 17923 3587
rect 18049 3587 18107 3593
rect 18049 3584 18061 3587
rect 17911 3556 18061 3584
rect 17911 3553 17923 3556
rect 17865 3547 17923 3553
rect 18049 3553 18061 3556
rect 18095 3584 18107 3587
rect 18414 3584 18420 3596
rect 18095 3556 18420 3584
rect 18095 3553 18107 3556
rect 18049 3547 18107 3553
rect 18414 3544 18420 3556
rect 18472 3544 18478 3596
rect 20622 3544 20628 3596
rect 20680 3544 20686 3596
rect 21818 3584 21824 3596
rect 20732 3556 21824 3584
rect 17310 3476 17316 3528
rect 17368 3476 17374 3528
rect 17405 3519 17463 3525
rect 17405 3485 17417 3519
rect 17451 3516 17463 3519
rect 17586 3516 17592 3528
rect 17451 3488 17592 3516
rect 17451 3485 17463 3488
rect 17405 3479 17463 3485
rect 16960 3420 17172 3448
rect 17221 3451 17279 3457
rect 16853 3411 16911 3417
rect 17221 3417 17233 3451
rect 17267 3448 17279 3451
rect 17420 3448 17448 3479
rect 17586 3476 17592 3488
rect 17644 3476 17650 3528
rect 18141 3519 18199 3525
rect 18141 3485 18153 3519
rect 18187 3516 18199 3519
rect 18230 3516 18236 3528
rect 18187 3488 18236 3516
rect 18187 3485 18199 3488
rect 18141 3479 18199 3485
rect 18230 3476 18236 3488
rect 18288 3476 18294 3528
rect 20070 3476 20076 3528
rect 20128 3476 20134 3528
rect 20165 3519 20223 3525
rect 20165 3485 20177 3519
rect 20211 3516 20223 3519
rect 20254 3516 20260 3528
rect 20211 3488 20260 3516
rect 20211 3485 20223 3488
rect 20165 3479 20223 3485
rect 20254 3476 20260 3488
rect 20312 3476 20318 3528
rect 20346 3476 20352 3528
rect 20404 3516 20410 3528
rect 20533 3519 20591 3525
rect 20533 3516 20545 3519
rect 20404 3488 20545 3516
rect 20404 3476 20410 3488
rect 20533 3485 20545 3488
rect 20579 3485 20591 3519
rect 20533 3479 20591 3485
rect 20732 3448 20760 3556
rect 20809 3519 20867 3525
rect 20809 3485 20821 3519
rect 20855 3518 20867 3519
rect 20855 3490 20944 3518
rect 20855 3485 20867 3490
rect 20809 3479 20867 3485
rect 17267 3420 17448 3448
rect 19306 3420 20760 3448
rect 17267 3417 17279 3420
rect 17221 3411 17279 3417
rect 13596 3352 15424 3380
rect 16209 3383 16267 3389
rect 13596 3340 13602 3352
rect 16209 3349 16221 3383
rect 16255 3380 16267 3383
rect 19306 3380 19334 3420
rect 16255 3352 19334 3380
rect 20257 3383 20315 3389
rect 16255 3349 16267 3352
rect 16209 3343 16267 3349
rect 20257 3349 20269 3383
rect 20303 3380 20315 3383
rect 20530 3380 20536 3392
rect 20303 3352 20536 3380
rect 20303 3349 20315 3352
rect 20257 3343 20315 3349
rect 20530 3340 20536 3352
rect 20588 3380 20594 3392
rect 20916 3380 20944 3490
rect 21008 3516 21036 3556
rect 21818 3544 21824 3556
rect 21876 3584 21882 3596
rect 22020 3584 22048 3624
rect 22097 3621 22109 3655
rect 22143 3652 22155 3655
rect 22370 3652 22376 3664
rect 22143 3624 22376 3652
rect 22143 3621 22155 3624
rect 22097 3615 22155 3621
rect 22370 3612 22376 3624
rect 22428 3612 22434 3664
rect 22741 3655 22799 3661
rect 22741 3621 22753 3655
rect 22787 3652 22799 3655
rect 23109 3655 23167 3661
rect 23109 3652 23121 3655
rect 22787 3624 23121 3652
rect 22787 3621 22799 3624
rect 22741 3615 22799 3621
rect 23109 3621 23121 3624
rect 23155 3652 23167 3655
rect 23155 3624 23980 3652
rect 23155 3621 23167 3624
rect 23109 3615 23167 3621
rect 23293 3587 23351 3593
rect 21876 3556 21956 3584
rect 21876 3544 21882 3556
rect 21073 3519 21131 3525
rect 21073 3516 21085 3519
rect 21008 3488 21085 3516
rect 21073 3485 21085 3488
rect 21119 3485 21131 3519
rect 21073 3479 21131 3485
rect 21266 3476 21272 3528
rect 21324 3476 21330 3528
rect 21634 3476 21640 3528
rect 21692 3516 21698 3528
rect 21928 3525 21956 3556
rect 22020 3556 22692 3584
rect 21729 3519 21787 3525
rect 21729 3516 21741 3519
rect 21692 3488 21741 3516
rect 21692 3476 21698 3488
rect 21729 3485 21741 3488
rect 21775 3485 21787 3519
rect 21729 3479 21787 3485
rect 21913 3519 21971 3525
rect 21913 3485 21925 3519
rect 21959 3485 21971 3519
rect 22020 3516 22048 3556
rect 22189 3519 22247 3525
rect 22189 3516 22201 3519
rect 22020 3488 22201 3516
rect 21913 3479 21971 3485
rect 22189 3485 22201 3488
rect 22235 3485 22247 3519
rect 22189 3479 22247 3485
rect 22370 3476 22376 3528
rect 22428 3476 22434 3528
rect 22557 3519 22615 3525
rect 22557 3485 22569 3519
rect 22603 3485 22615 3519
rect 22664 3516 22692 3556
rect 23293 3553 23305 3587
rect 23339 3584 23351 3587
rect 23339 3556 23888 3584
rect 23339 3553 23351 3556
rect 23293 3547 23351 3553
rect 23385 3519 23443 3525
rect 23385 3516 23397 3519
rect 22664 3488 23397 3516
rect 22557 3479 22615 3485
rect 23385 3485 23397 3488
rect 23431 3485 23443 3519
rect 23385 3479 23443 3485
rect 23569 3519 23627 3525
rect 23569 3485 23581 3519
rect 23615 3485 23627 3519
rect 23569 3479 23627 3485
rect 20993 3451 21051 3457
rect 20993 3417 21005 3451
rect 21039 3448 21051 3451
rect 21039 3420 21404 3448
rect 21039 3417 21051 3420
rect 20993 3411 21051 3417
rect 21177 3383 21235 3389
rect 21177 3380 21189 3383
rect 20588 3352 21189 3380
rect 20588 3340 20594 3352
rect 21177 3349 21189 3352
rect 21223 3349 21235 3383
rect 21376 3380 21404 3420
rect 21450 3408 21456 3460
rect 21508 3408 21514 3460
rect 22462 3408 22468 3460
rect 22520 3408 22526 3460
rect 21910 3380 21916 3392
rect 21376 3352 21916 3380
rect 21177 3343 21235 3349
rect 21910 3340 21916 3352
rect 21968 3380 21974 3392
rect 22572 3380 22600 3479
rect 22833 3451 22891 3457
rect 22833 3417 22845 3451
rect 22879 3448 22891 3451
rect 23474 3448 23480 3460
rect 22879 3420 23480 3448
rect 22879 3417 22891 3420
rect 22833 3411 22891 3417
rect 23474 3408 23480 3420
rect 23532 3448 23538 3460
rect 23584 3448 23612 3479
rect 23658 3476 23664 3528
rect 23716 3476 23722 3528
rect 23860 3525 23888 3556
rect 23845 3519 23903 3525
rect 23845 3485 23857 3519
rect 23891 3485 23903 3519
rect 23952 3516 23980 3624
rect 24854 3612 24860 3664
rect 24912 3612 24918 3664
rect 25225 3655 25283 3661
rect 25225 3621 25237 3655
rect 25271 3652 25283 3655
rect 25682 3652 25688 3664
rect 25271 3624 25688 3652
rect 25271 3621 25283 3624
rect 25225 3615 25283 3621
rect 25682 3612 25688 3624
rect 25740 3612 25746 3664
rect 24872 3584 24900 3612
rect 24949 3587 25007 3593
rect 24949 3584 24961 3587
rect 24872 3556 24961 3584
rect 24949 3553 24961 3556
rect 24995 3553 25007 3587
rect 24949 3547 25007 3553
rect 24857 3519 24915 3525
rect 24857 3516 24869 3519
rect 23952 3488 24869 3516
rect 23845 3479 23903 3485
rect 24857 3485 24869 3488
rect 24903 3485 24915 3519
rect 24857 3479 24915 3485
rect 24670 3448 24676 3460
rect 23532 3420 24676 3448
rect 23532 3408 23538 3420
rect 24670 3408 24676 3420
rect 24728 3408 24734 3460
rect 21968 3352 22600 3380
rect 21968 3340 21974 3352
rect 1104 3290 27876 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 27876 3290
rect 1104 3216 27876 3238
rect 10134 3136 10140 3188
rect 10192 3136 10198 3188
rect 10873 3179 10931 3185
rect 10873 3176 10885 3179
rect 10428 3148 10885 3176
rect 10428 3117 10456 3148
rect 10873 3145 10885 3148
rect 10919 3145 10931 3179
rect 10873 3139 10931 3145
rect 11146 3136 11152 3188
rect 11204 3176 11210 3188
rect 15654 3176 15660 3188
rect 11204 3148 13768 3176
rect 11204 3136 11210 3148
rect 10413 3111 10471 3117
rect 10413 3077 10425 3111
rect 10459 3077 10471 3111
rect 10413 3071 10471 3077
rect 10502 3068 10508 3120
rect 10560 3108 10566 3120
rect 11606 3108 11612 3120
rect 10560 3080 11612 3108
rect 10560 3068 10566 3080
rect 11606 3068 11612 3080
rect 11664 3068 11670 3120
rect 12529 3111 12587 3117
rect 12529 3077 12541 3111
rect 12575 3108 12587 3111
rect 12575 3080 13492 3108
rect 12575 3077 12587 3080
rect 12529 3071 12587 3077
rect 9769 3043 9827 3049
rect 9769 3009 9781 3043
rect 9815 3040 9827 3043
rect 9950 3040 9956 3052
rect 9815 3012 9956 3040
rect 9815 3009 9827 3012
rect 9769 3003 9827 3009
rect 9950 3000 9956 3012
rect 10008 3000 10014 3052
rect 10226 3000 10232 3052
rect 10284 3000 10290 3052
rect 10597 3043 10655 3049
rect 10597 3009 10609 3043
rect 10643 3009 10655 3043
rect 10597 3003 10655 3009
rect 842 2932 848 2984
rect 900 2972 906 2984
rect 1397 2975 1455 2981
rect 1397 2972 1409 2975
rect 900 2944 1409 2972
rect 900 2932 906 2944
rect 1397 2941 1409 2944
rect 1443 2941 1455 2975
rect 1397 2935 1455 2941
rect 9861 2975 9919 2981
rect 9861 2941 9873 2975
rect 9907 2972 9919 2975
rect 10410 2972 10416 2984
rect 9907 2944 10416 2972
rect 9907 2941 9919 2944
rect 9861 2935 9919 2941
rect 10410 2932 10416 2944
rect 10468 2972 10474 2984
rect 10612 2972 10640 3003
rect 10870 3000 10876 3052
rect 10928 3040 10934 3052
rect 11057 3043 11115 3049
rect 11057 3040 11069 3043
rect 10928 3012 11069 3040
rect 10928 3000 10934 3012
rect 11057 3009 11069 3012
rect 11103 3009 11115 3043
rect 11057 3003 11115 3009
rect 11146 3000 11152 3052
rect 11204 3040 11210 3052
rect 11241 3043 11299 3049
rect 11241 3040 11253 3043
rect 11204 3012 11253 3040
rect 11204 3000 11210 3012
rect 11241 3009 11253 3012
rect 11287 3009 11299 3043
rect 11241 3003 11299 3009
rect 11790 3000 11796 3052
rect 11848 3040 11854 3052
rect 11977 3043 12035 3049
rect 11977 3040 11989 3043
rect 11848 3012 11989 3040
rect 11848 3000 11854 3012
rect 11977 3009 11989 3012
rect 12023 3040 12035 3043
rect 12437 3043 12495 3049
rect 12437 3040 12449 3043
rect 12023 3012 12449 3040
rect 12023 3009 12035 3012
rect 11977 3003 12035 3009
rect 12437 3009 12449 3012
rect 12483 3009 12495 3043
rect 12437 3003 12495 3009
rect 12621 3043 12679 3049
rect 12621 3009 12633 3043
rect 12667 3009 12679 3043
rect 12621 3003 12679 3009
rect 10468 2944 10640 2972
rect 10468 2932 10474 2944
rect 12066 2932 12072 2984
rect 12124 2972 12130 2984
rect 12636 2972 12664 3003
rect 13262 3000 13268 3052
rect 13320 3000 13326 3052
rect 13464 3049 13492 3080
rect 13449 3043 13507 3049
rect 13449 3009 13461 3043
rect 13495 3009 13507 3043
rect 13449 3003 13507 3009
rect 13740 3030 13768 3148
rect 15212 3148 15660 3176
rect 15212 3108 15240 3148
rect 15654 3136 15660 3148
rect 15712 3136 15718 3188
rect 15930 3136 15936 3188
rect 15988 3136 15994 3188
rect 16393 3179 16451 3185
rect 16393 3145 16405 3179
rect 16439 3176 16451 3179
rect 16574 3176 16580 3188
rect 16439 3148 16580 3176
rect 16439 3145 16451 3148
rect 16393 3139 16451 3145
rect 16574 3136 16580 3148
rect 16632 3176 16638 3188
rect 16961 3179 17019 3185
rect 16961 3176 16973 3179
rect 16632 3148 16973 3176
rect 16632 3136 16638 3148
rect 16961 3145 16973 3148
rect 17007 3145 17019 3179
rect 16961 3139 17019 3145
rect 17221 3179 17279 3185
rect 17221 3145 17233 3179
rect 17267 3176 17279 3179
rect 19705 3179 19763 3185
rect 17267 3148 19656 3176
rect 17267 3145 17279 3148
rect 17221 3139 17279 3145
rect 14398 3080 15240 3108
rect 15286 3068 15292 3120
rect 15344 3108 15350 3120
rect 15746 3108 15752 3120
rect 15344 3080 15752 3108
rect 15344 3068 15350 3080
rect 15746 3068 15752 3080
rect 15804 3108 15810 3120
rect 16025 3111 16083 3117
rect 16025 3108 16037 3111
rect 15804 3080 16037 3108
rect 15804 3068 15810 3080
rect 16025 3077 16037 3080
rect 16071 3077 16083 3111
rect 16025 3071 16083 3077
rect 16206 3068 16212 3120
rect 16264 3068 16270 3120
rect 16761 3111 16819 3117
rect 16761 3077 16773 3111
rect 16807 3108 16819 3111
rect 19628 3108 19656 3148
rect 19705 3145 19717 3179
rect 19751 3176 19763 3179
rect 20070 3176 20076 3188
rect 19751 3148 20076 3176
rect 19751 3145 19763 3148
rect 19705 3139 19763 3145
rect 20070 3136 20076 3148
rect 20128 3136 20134 3188
rect 20162 3136 20168 3188
rect 20220 3176 20226 3188
rect 20441 3179 20499 3185
rect 20441 3176 20453 3179
rect 20220 3148 20453 3176
rect 20220 3136 20226 3148
rect 20441 3145 20453 3148
rect 20487 3145 20499 3179
rect 20441 3139 20499 3145
rect 21361 3179 21419 3185
rect 21361 3145 21373 3179
rect 21407 3176 21419 3179
rect 21726 3176 21732 3188
rect 21407 3148 21732 3176
rect 21407 3145 21419 3148
rect 21361 3139 21419 3145
rect 21726 3136 21732 3148
rect 21784 3136 21790 3188
rect 22189 3179 22247 3185
rect 22189 3176 22201 3179
rect 22066 3148 22201 3176
rect 20625 3111 20683 3117
rect 16807 3080 18184 3108
rect 19628 3080 20300 3108
rect 16807 3077 16819 3080
rect 16761 3071 16819 3077
rect 15194 3040 15200 3052
rect 13924 3030 15200 3040
rect 13740 3012 15200 3030
rect 13740 3002 13952 3012
rect 15194 3000 15200 3012
rect 15252 3000 15258 3052
rect 15562 3000 15568 3052
rect 15620 3000 15626 3052
rect 15654 3000 15660 3052
rect 15712 3040 15718 3052
rect 16776 3040 16804 3071
rect 15712 3012 16804 3040
rect 15712 3000 15718 3012
rect 17126 3000 17132 3052
rect 17184 3040 17190 3052
rect 17405 3043 17463 3049
rect 17405 3040 17417 3043
rect 17184 3012 17417 3040
rect 17184 3000 17190 3012
rect 17405 3009 17417 3012
rect 17451 3040 17463 3043
rect 17770 3040 17776 3052
rect 17451 3012 17776 3040
rect 17451 3009 17463 3012
rect 17405 3003 17463 3009
rect 17770 3000 17776 3012
rect 17828 3000 17834 3052
rect 18156 3049 18184 3080
rect 18141 3043 18199 3049
rect 18141 3009 18153 3043
rect 18187 3009 18199 3043
rect 18141 3003 18199 3009
rect 18230 3000 18236 3052
rect 18288 3040 18294 3052
rect 18325 3043 18383 3049
rect 18325 3040 18337 3043
rect 18288 3012 18337 3040
rect 18288 3000 18294 3012
rect 18325 3009 18337 3012
rect 18371 3009 18383 3043
rect 18325 3003 18383 3009
rect 18414 3000 18420 3052
rect 18472 3000 18478 3052
rect 18690 3000 18696 3052
rect 18748 3000 18754 3052
rect 18874 3000 18880 3052
rect 18932 3040 18938 3052
rect 19981 3043 20039 3049
rect 19981 3040 19993 3043
rect 18932 3012 19993 3040
rect 18932 3000 18938 3012
rect 19981 3009 19993 3012
rect 20027 3009 20039 3043
rect 19981 3003 20039 3009
rect 12124 2944 12664 2972
rect 16868 2944 17448 2972
rect 12124 2932 12130 2944
rect 10781 2907 10839 2913
rect 10781 2873 10793 2907
rect 10827 2904 10839 2907
rect 12345 2907 12403 2913
rect 10827 2876 11652 2904
rect 10827 2873 10839 2876
rect 10781 2867 10839 2873
rect 9950 2796 9956 2848
rect 10008 2836 10014 2848
rect 11057 2839 11115 2845
rect 11057 2836 11069 2839
rect 10008 2808 11069 2836
rect 10008 2796 10014 2808
rect 11057 2805 11069 2808
rect 11103 2805 11115 2839
rect 11624 2836 11652 2876
rect 12345 2873 12357 2907
rect 12391 2904 12403 2907
rect 13630 2904 13636 2916
rect 12391 2876 13636 2904
rect 12391 2873 12403 2876
rect 12345 2867 12403 2873
rect 13630 2864 13636 2876
rect 13688 2864 13694 2916
rect 15212 2876 15884 2904
rect 13446 2836 13452 2848
rect 11624 2808 13452 2836
rect 11057 2799 11115 2805
rect 13446 2796 13452 2808
rect 13504 2836 13510 2848
rect 15212 2836 15240 2876
rect 13504 2808 15240 2836
rect 15856 2836 15884 2876
rect 16868 2836 16896 2944
rect 17126 2864 17132 2916
rect 17184 2864 17190 2916
rect 17420 2904 17448 2944
rect 17494 2932 17500 2984
rect 17552 2932 17558 2984
rect 17865 2975 17923 2981
rect 17865 2941 17877 2975
rect 17911 2972 17923 2975
rect 17957 2975 18015 2981
rect 17957 2972 17969 2975
rect 17911 2944 17969 2972
rect 17911 2941 17923 2944
rect 17865 2935 17923 2941
rect 17957 2941 17969 2944
rect 18003 2941 18015 2975
rect 17957 2935 18015 2941
rect 18248 2904 18276 3000
rect 19889 2975 19947 2981
rect 19889 2941 19901 2975
rect 19935 2941 19947 2975
rect 19889 2935 19947 2941
rect 17420 2876 18276 2904
rect 18690 2864 18696 2916
rect 18748 2904 18754 2916
rect 19904 2904 19932 2935
rect 18748 2876 19932 2904
rect 20272 2904 20300 3080
rect 20625 3077 20637 3111
rect 20671 3108 20683 3111
rect 22066 3108 22094 3148
rect 22189 3145 22201 3148
rect 22235 3176 22247 3179
rect 22462 3176 22468 3188
rect 22235 3148 22468 3176
rect 22235 3145 22247 3148
rect 22189 3139 22247 3145
rect 22462 3136 22468 3148
rect 22520 3136 22526 3188
rect 22557 3179 22615 3185
rect 22557 3145 22569 3179
rect 22603 3176 22615 3179
rect 23658 3176 23664 3188
rect 22603 3148 23664 3176
rect 22603 3145 22615 3148
rect 22557 3139 22615 3145
rect 23658 3136 23664 3148
rect 23716 3136 23722 3188
rect 20671 3080 22094 3108
rect 20671 3077 20683 3080
rect 20625 3071 20683 3077
rect 20349 2975 20407 2981
rect 20349 2941 20361 2975
rect 20395 2972 20407 2975
rect 20640 2972 20668 3071
rect 21284 3049 21312 3080
rect 20809 3043 20867 3049
rect 20809 3009 20821 3043
rect 20855 3009 20867 3043
rect 20809 3003 20867 3009
rect 21269 3043 21327 3049
rect 21269 3009 21281 3043
rect 21315 3009 21327 3043
rect 21269 3003 21327 3009
rect 21453 3043 21511 3049
rect 21453 3009 21465 3043
rect 21499 3040 21511 3043
rect 22097 3043 22155 3049
rect 22097 3040 22109 3043
rect 21499 3012 22109 3040
rect 21499 3009 21511 3012
rect 21453 3003 21511 3009
rect 22097 3009 22109 3012
rect 22143 3009 22155 3043
rect 22097 3003 22155 3009
rect 20395 2944 20668 2972
rect 20824 2972 20852 3003
rect 21468 2972 21496 3003
rect 20824 2944 21496 2972
rect 20395 2941 20407 2944
rect 20349 2935 20407 2941
rect 20824 2904 20852 2944
rect 21910 2932 21916 2984
rect 21968 2932 21974 2984
rect 27522 2932 27528 2984
rect 27580 2932 27586 2984
rect 20272 2876 20852 2904
rect 18748 2864 18754 2876
rect 16945 2839 17003 2845
rect 16945 2836 16957 2839
rect 15856 2808 16957 2836
rect 13504 2796 13510 2808
rect 16945 2805 16957 2808
rect 16991 2805 17003 2839
rect 16945 2799 17003 2805
rect 1104 2746 27876 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 27876 2746
rect 1104 2672 27876 2694
rect 10410 2592 10416 2644
rect 10468 2592 10474 2644
rect 12066 2592 12072 2644
rect 12124 2592 12130 2644
rect 13538 2592 13544 2644
rect 13596 2592 13602 2644
rect 15565 2635 15623 2641
rect 15565 2601 15577 2635
rect 15611 2632 15623 2635
rect 16390 2632 16396 2644
rect 15611 2604 16396 2632
rect 15611 2601 15623 2604
rect 15565 2595 15623 2601
rect 16390 2592 16396 2604
rect 16448 2592 16454 2644
rect 17865 2635 17923 2641
rect 17865 2601 17877 2635
rect 17911 2632 17923 2635
rect 18690 2632 18696 2644
rect 17911 2604 18696 2632
rect 17911 2601 17923 2604
rect 17865 2595 17923 2601
rect 18690 2592 18696 2604
rect 18748 2592 18754 2644
rect 15194 2524 15200 2576
rect 15252 2564 15258 2576
rect 15381 2567 15439 2573
rect 15381 2564 15393 2567
rect 15252 2536 15393 2564
rect 15252 2524 15258 2536
rect 15381 2533 15393 2536
rect 15427 2533 15439 2567
rect 15381 2527 15439 2533
rect 10962 2496 10968 2508
rect 10244 2468 10968 2496
rect 10244 2437 10272 2468
rect 10962 2456 10968 2468
rect 11020 2456 11026 2508
rect 15396 2496 15424 2527
rect 15746 2524 15752 2576
rect 15804 2524 15810 2576
rect 15396 2468 15700 2496
rect 10229 2431 10287 2437
rect 10229 2397 10241 2431
rect 10275 2397 10287 2431
rect 10229 2391 10287 2397
rect 10413 2431 10471 2437
rect 10413 2397 10425 2431
rect 10459 2428 10471 2431
rect 11238 2428 11244 2440
rect 10459 2400 11244 2428
rect 10459 2397 10471 2400
rect 10413 2391 10471 2397
rect 11238 2388 11244 2400
rect 11296 2388 11302 2440
rect 11606 2388 11612 2440
rect 11664 2388 11670 2440
rect 11885 2431 11943 2437
rect 11885 2397 11897 2431
rect 11931 2397 11943 2431
rect 11885 2391 11943 2397
rect 11256 2360 11284 2388
rect 11900 2360 11928 2391
rect 13446 2388 13452 2440
rect 13504 2388 13510 2440
rect 13630 2388 13636 2440
rect 13688 2388 13694 2440
rect 15105 2431 15163 2437
rect 15105 2397 15117 2431
rect 15151 2428 15163 2431
rect 15378 2428 15384 2440
rect 15151 2400 15384 2428
rect 15151 2397 15163 2400
rect 15105 2391 15163 2397
rect 15378 2388 15384 2400
rect 15436 2388 15442 2440
rect 15672 2437 15700 2468
rect 15657 2431 15715 2437
rect 15657 2397 15669 2431
rect 15703 2397 15715 2431
rect 15657 2391 15715 2397
rect 15838 2388 15844 2440
rect 15896 2388 15902 2440
rect 16942 2388 16948 2440
rect 17000 2428 17006 2440
rect 17681 2431 17739 2437
rect 17681 2428 17693 2431
rect 17000 2400 17693 2428
rect 17000 2388 17006 2400
rect 17681 2397 17693 2400
rect 17727 2397 17739 2431
rect 17681 2391 17739 2397
rect 17770 2388 17776 2440
rect 17828 2428 17834 2440
rect 17865 2431 17923 2437
rect 17865 2428 17877 2431
rect 17828 2400 17877 2428
rect 17828 2388 17834 2400
rect 17865 2397 17877 2400
rect 17911 2397 17923 2431
rect 17865 2391 17923 2397
rect 11256 2332 11928 2360
rect 13648 2360 13676 2388
rect 15562 2360 15568 2372
rect 13648 2332 15568 2360
rect 15562 2320 15568 2332
rect 15620 2320 15626 2372
rect 11701 2295 11759 2301
rect 11701 2261 11713 2295
rect 11747 2292 11759 2295
rect 11882 2292 11888 2304
rect 11747 2264 11888 2292
rect 11747 2261 11759 2264
rect 11701 2255 11759 2261
rect 11882 2252 11888 2264
rect 11940 2252 11946 2304
rect 1104 2202 27876 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 27876 2202
rect 1104 2128 27876 2150
<< via1 >>
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 5816 28704 5868 28756
rect 6460 28704 6512 28756
rect 9036 28704 9088 28756
rect 3240 28568 3292 28620
rect 4620 28500 4672 28552
rect 5540 28500 5592 28552
rect 6184 28500 6236 28552
rect 8392 28500 8444 28552
rect 9128 28500 9180 28552
rect 9680 28543 9732 28552
rect 9680 28509 9689 28543
rect 9689 28509 9723 28543
rect 9723 28509 9732 28543
rect 9680 28500 9732 28509
rect 4712 28475 4764 28484
rect 4712 28441 4721 28475
rect 4721 28441 4755 28475
rect 4755 28441 4764 28475
rect 4712 28432 4764 28441
rect 7748 28432 7800 28484
rect 12532 28543 12584 28552
rect 12532 28509 12541 28543
rect 12541 28509 12575 28543
rect 12575 28509 12584 28543
rect 12532 28500 12584 28509
rect 17040 28543 17092 28552
rect 17040 28509 17049 28543
rect 17049 28509 17083 28543
rect 17083 28509 17092 28543
rect 17040 28500 17092 28509
rect 13176 28432 13228 28484
rect 16856 28432 16908 28484
rect 6552 28364 6604 28416
rect 7288 28364 7340 28416
rect 8484 28407 8536 28416
rect 8484 28373 8493 28407
rect 8493 28373 8527 28407
rect 8527 28373 8536 28407
rect 8484 28364 8536 28373
rect 12716 28364 12768 28416
rect 17132 28407 17184 28416
rect 17132 28373 17141 28407
rect 17141 28373 17175 28407
rect 17175 28373 17184 28407
rect 17132 28364 17184 28373
rect 4874 28262 4926 28314
rect 4938 28262 4990 28314
rect 5002 28262 5054 28314
rect 5066 28262 5118 28314
rect 5130 28262 5182 28314
rect 4712 28160 4764 28212
rect 6184 28203 6236 28212
rect 6184 28169 6193 28203
rect 6193 28169 6227 28203
rect 6227 28169 6236 28203
rect 6184 28160 6236 28169
rect 2964 28092 3016 28144
rect 4804 28092 4856 28144
rect 1768 28024 1820 28076
rect 1860 28067 1912 28076
rect 1860 28033 1869 28067
rect 1869 28033 1903 28067
rect 1903 28033 1912 28067
rect 1860 28024 1912 28033
rect 3332 28024 3384 28076
rect 1400 27956 1452 28008
rect 4896 28024 4948 28076
rect 5632 28024 5684 28076
rect 5816 28067 5868 28076
rect 5816 28033 5825 28067
rect 5825 28033 5859 28067
rect 5859 28033 5868 28067
rect 5816 28024 5868 28033
rect 5908 28067 5960 28076
rect 5908 28033 5917 28067
rect 5917 28033 5951 28067
rect 5951 28033 5960 28067
rect 5908 28024 5960 28033
rect 6552 28135 6604 28144
rect 6552 28101 6561 28135
rect 6561 28101 6595 28135
rect 6595 28101 6604 28135
rect 6552 28092 6604 28101
rect 6644 28067 6696 28076
rect 6276 27956 6328 28008
rect 6644 28033 6653 28067
rect 6653 28033 6687 28067
rect 6687 28033 6696 28067
rect 6644 28024 6696 28033
rect 6736 28067 6788 28076
rect 6736 28033 6745 28067
rect 6745 28033 6779 28067
rect 6779 28033 6788 28067
rect 6736 28024 6788 28033
rect 7104 28160 7156 28212
rect 9128 28203 9180 28212
rect 9128 28169 9137 28203
rect 9137 28169 9171 28203
rect 9171 28169 9180 28203
rect 9128 28160 9180 28169
rect 8484 28092 8536 28144
rect 9680 28160 9732 28212
rect 16580 28160 16632 28212
rect 17040 28160 17092 28212
rect 10416 28067 10468 28076
rect 14096 28092 14148 28144
rect 10416 28033 10434 28067
rect 10434 28033 10468 28067
rect 10416 28024 10468 28033
rect 12716 28024 12768 28076
rect 14740 28067 14792 28076
rect 14740 28033 14774 28067
rect 14774 28033 14792 28067
rect 14740 28024 14792 28033
rect 18604 28092 18656 28144
rect 7748 27999 7800 28008
rect 7748 27965 7757 27999
rect 7757 27965 7791 27999
rect 7791 27965 7800 27999
rect 7748 27956 7800 27965
rect 10876 27956 10928 28008
rect 10968 27888 11020 27940
rect 12624 27888 12676 27940
rect 1676 27863 1728 27872
rect 1676 27829 1685 27863
rect 1685 27829 1719 27863
rect 1719 27829 1728 27863
rect 1676 27820 1728 27829
rect 3884 27863 3936 27872
rect 3884 27829 3893 27863
rect 3893 27829 3927 27863
rect 3927 27829 3936 27863
rect 3884 27820 3936 27829
rect 4804 27863 4856 27872
rect 4804 27829 4813 27863
rect 4813 27829 4847 27863
rect 4847 27829 4856 27863
rect 4804 27820 4856 27829
rect 5816 27820 5868 27872
rect 6276 27820 6328 27872
rect 11336 27863 11388 27872
rect 11336 27829 11345 27863
rect 11345 27829 11379 27863
rect 11379 27829 11388 27863
rect 11336 27820 11388 27829
rect 14004 27863 14056 27872
rect 14004 27829 14013 27863
rect 14013 27829 14047 27863
rect 14047 27829 14056 27863
rect 14004 27820 14056 27829
rect 15752 27820 15804 27872
rect 16120 27863 16172 27872
rect 16120 27829 16129 27863
rect 16129 27829 16163 27863
rect 16163 27829 16172 27863
rect 16120 27820 16172 27829
rect 16764 28024 16816 28076
rect 16856 27820 16908 27872
rect 18144 27863 18196 27872
rect 18144 27829 18153 27863
rect 18153 27829 18187 27863
rect 18187 27829 18196 27863
rect 18144 27820 18196 27829
rect 18236 27820 18288 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 3148 27659 3200 27668
rect 3148 27625 3157 27659
rect 3157 27625 3191 27659
rect 3191 27625 3200 27659
rect 3148 27616 3200 27625
rect 4712 27616 4764 27668
rect 6644 27616 6696 27668
rect 12532 27616 12584 27668
rect 17132 27616 17184 27668
rect 4620 27548 4672 27600
rect 5908 27548 5960 27600
rect 6276 27591 6328 27600
rect 6276 27557 6285 27591
rect 6285 27557 6319 27591
rect 6319 27557 6328 27591
rect 6276 27548 6328 27557
rect 10416 27591 10468 27600
rect 10416 27557 10425 27591
rect 10425 27557 10459 27591
rect 10459 27557 10468 27591
rect 10416 27548 10468 27557
rect 1400 27523 1452 27532
rect 1400 27489 1409 27523
rect 1409 27489 1443 27523
rect 1443 27489 1452 27523
rect 1400 27480 1452 27489
rect 2412 27480 2464 27532
rect 9680 27523 9732 27532
rect 9680 27489 9689 27523
rect 9689 27489 9723 27523
rect 9723 27489 9732 27523
rect 9680 27480 9732 27489
rect 1676 27455 1728 27464
rect 1676 27421 1710 27455
rect 1710 27421 1728 27455
rect 1676 27412 1728 27421
rect 3332 27412 3384 27464
rect 3424 27455 3476 27464
rect 3424 27421 3433 27455
rect 3433 27421 3467 27455
rect 3467 27421 3476 27455
rect 3424 27412 3476 27421
rect 3700 27412 3752 27464
rect 2596 27344 2648 27396
rect 3884 27344 3936 27396
rect 4804 27455 4856 27464
rect 4804 27421 4813 27455
rect 4813 27421 4847 27455
rect 4847 27421 4856 27455
rect 4804 27412 4856 27421
rect 6184 27455 6236 27464
rect 6184 27421 6193 27455
rect 6193 27421 6227 27455
rect 6227 27421 6236 27455
rect 6184 27412 6236 27421
rect 8852 27412 8904 27464
rect 6828 27344 6880 27396
rect 7472 27344 7524 27396
rect 7656 27387 7708 27396
rect 7656 27353 7690 27387
rect 7690 27353 7708 27387
rect 7656 27344 7708 27353
rect 7748 27344 7800 27396
rect 10876 27480 10928 27532
rect 16764 27548 16816 27600
rect 18236 27548 18288 27600
rect 14004 27480 14056 27532
rect 17132 27480 17184 27532
rect 18144 27480 18196 27532
rect 11336 27412 11388 27464
rect 13636 27455 13688 27464
rect 13636 27421 13645 27455
rect 13645 27421 13679 27455
rect 13679 27421 13688 27455
rect 13636 27412 13688 27421
rect 15752 27455 15804 27464
rect 3424 27276 3476 27328
rect 3792 27319 3844 27328
rect 3792 27285 3801 27319
rect 3801 27285 3835 27319
rect 3835 27285 3844 27319
rect 3792 27276 3844 27285
rect 6368 27276 6420 27328
rect 8760 27319 8812 27328
rect 8760 27285 8769 27319
rect 8769 27285 8803 27319
rect 8803 27285 8812 27319
rect 8760 27276 8812 27285
rect 13360 27344 13412 27396
rect 13544 27344 13596 27396
rect 15752 27421 15761 27455
rect 15761 27421 15795 27455
rect 15795 27421 15804 27455
rect 15752 27412 15804 27421
rect 12624 27319 12676 27328
rect 12624 27285 12633 27319
rect 12633 27285 12667 27319
rect 12667 27285 12676 27319
rect 12624 27276 12676 27285
rect 15660 27344 15712 27396
rect 16120 27344 16172 27396
rect 14280 27276 14332 27328
rect 4874 27174 4926 27226
rect 4938 27174 4990 27226
rect 5002 27174 5054 27226
rect 5066 27174 5118 27226
rect 5130 27174 5182 27226
rect 1768 27072 1820 27124
rect 1860 27072 1912 27124
rect 3792 27072 3844 27124
rect 7656 27072 7708 27124
rect 2044 26936 2096 26988
rect 2412 26979 2464 26988
rect 2412 26945 2421 26979
rect 2421 26945 2455 26979
rect 2455 26945 2464 26979
rect 2412 26936 2464 26945
rect 2596 26979 2648 26988
rect 2596 26945 2605 26979
rect 2605 26945 2639 26979
rect 2639 26945 2648 26979
rect 2596 26936 2648 26945
rect 4160 27004 4212 27056
rect 4804 27004 4856 27056
rect 8116 27047 8168 27056
rect 8116 27013 8143 27047
rect 8143 27013 8168 27047
rect 8116 27004 8168 27013
rect 8300 27047 8352 27056
rect 8300 27013 8309 27047
rect 8309 27013 8343 27047
rect 8343 27013 8352 27047
rect 8300 27004 8352 27013
rect 2872 26911 2924 26920
rect 2872 26877 2881 26911
rect 2881 26877 2915 26911
rect 2915 26877 2924 26911
rect 2872 26868 2924 26877
rect 4620 26936 4672 26988
rect 5816 26936 5868 26988
rect 6644 26936 6696 26988
rect 9312 26979 9364 26988
rect 9312 26945 9321 26979
rect 9321 26945 9355 26979
rect 9355 26945 9364 26979
rect 9312 26936 9364 26945
rect 9496 26979 9548 26988
rect 9496 26945 9505 26979
rect 9505 26945 9539 26979
rect 9539 26945 9548 26979
rect 9496 26936 9548 26945
rect 12440 26979 12492 26988
rect 12440 26945 12449 26979
rect 12449 26945 12483 26979
rect 12483 26945 12492 26979
rect 12440 26936 12492 26945
rect 13912 27072 13964 27124
rect 13544 27047 13596 27056
rect 13544 27013 13553 27047
rect 13553 27013 13587 27047
rect 13587 27013 13596 27047
rect 13544 27004 13596 27013
rect 13820 27047 13872 27056
rect 13820 27013 13847 27047
rect 13847 27013 13872 27047
rect 13820 27004 13872 27013
rect 14188 27072 14240 27124
rect 15660 27072 15712 27124
rect 13636 26936 13688 26988
rect 9404 26868 9456 26920
rect 12992 26868 13044 26920
rect 14280 26979 14332 26988
rect 14280 26945 14289 26979
rect 14289 26945 14323 26979
rect 14323 26945 14332 26979
rect 14280 26936 14332 26945
rect 14372 26936 14424 26988
rect 15476 26979 15528 26988
rect 15476 26945 15485 26979
rect 15485 26945 15519 26979
rect 15519 26945 15528 26979
rect 15476 26936 15528 26945
rect 16028 26936 16080 26988
rect 16488 26936 16540 26988
rect 16856 26936 16908 26988
rect 17316 26936 17368 26988
rect 18512 26979 18564 26988
rect 18512 26945 18521 26979
rect 18521 26945 18555 26979
rect 18555 26945 18564 26979
rect 18512 26936 18564 26945
rect 18604 26979 18656 26988
rect 18604 26945 18613 26979
rect 18613 26945 18647 26979
rect 18647 26945 18656 26979
rect 18604 26936 18656 26945
rect 20996 26979 21048 26988
rect 20996 26945 21005 26979
rect 21005 26945 21039 26979
rect 21039 26945 21048 26979
rect 20996 26936 21048 26945
rect 1952 26732 2004 26784
rect 2964 26775 3016 26784
rect 2964 26741 2973 26775
rect 2973 26741 3007 26775
rect 3007 26741 3016 26775
rect 2964 26732 3016 26741
rect 4804 26732 4856 26784
rect 5172 26775 5224 26784
rect 5172 26741 5181 26775
rect 5181 26741 5215 26775
rect 5215 26741 5224 26775
rect 5172 26732 5224 26741
rect 7196 26732 7248 26784
rect 7380 26732 7432 26784
rect 7840 26732 7892 26784
rect 10600 26775 10652 26784
rect 10600 26741 10609 26775
rect 10609 26741 10643 26775
rect 10643 26741 10652 26775
rect 10600 26732 10652 26741
rect 12624 26775 12676 26784
rect 12624 26741 12633 26775
rect 12633 26741 12667 26775
rect 12667 26741 12676 26775
rect 12624 26732 12676 26741
rect 13176 26775 13228 26784
rect 13176 26741 13185 26775
rect 13185 26741 13219 26775
rect 13219 26741 13228 26775
rect 13176 26732 13228 26741
rect 14004 26800 14056 26852
rect 14740 26868 14792 26920
rect 16120 26911 16172 26920
rect 16120 26877 16129 26911
rect 16129 26877 16163 26911
rect 16163 26877 16172 26911
rect 16120 26868 16172 26877
rect 17132 26911 17184 26920
rect 17132 26877 17141 26911
rect 17141 26877 17175 26911
rect 17175 26877 17184 26911
rect 17132 26868 17184 26877
rect 13636 26775 13688 26784
rect 13636 26741 13645 26775
rect 13645 26741 13679 26775
rect 13679 26741 13688 26775
rect 13636 26732 13688 26741
rect 14280 26732 14332 26784
rect 14372 26732 14424 26784
rect 17500 26843 17552 26852
rect 17500 26809 17509 26843
rect 17509 26809 17543 26843
rect 17543 26809 17552 26843
rect 17500 26800 17552 26809
rect 17592 26775 17644 26784
rect 17592 26741 17601 26775
rect 17601 26741 17635 26775
rect 17635 26741 17644 26775
rect 17592 26732 17644 26741
rect 20076 26775 20128 26784
rect 20076 26741 20085 26775
rect 20085 26741 20119 26775
rect 20119 26741 20128 26775
rect 20076 26732 20128 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 1216 26528 1268 26580
rect 3792 26528 3844 26580
rect 4620 26528 4672 26580
rect 1860 26324 1912 26376
rect 3884 26392 3936 26444
rect 2964 26324 3016 26376
rect 3148 26324 3200 26376
rect 3332 26324 3384 26376
rect 3700 26324 3752 26376
rect 4436 26324 4488 26376
rect 4804 26367 4856 26376
rect 4804 26333 4821 26367
rect 4821 26333 4856 26367
rect 4804 26324 4856 26333
rect 5172 26460 5224 26512
rect 5356 26460 5408 26512
rect 5264 26435 5316 26444
rect 5264 26401 5273 26435
rect 5273 26401 5307 26435
rect 5307 26401 5316 26435
rect 5264 26392 5316 26401
rect 4988 26367 5040 26376
rect 4988 26333 4997 26367
rect 4997 26333 5031 26367
rect 5031 26333 5040 26367
rect 4988 26324 5040 26333
rect 5632 26528 5684 26580
rect 6460 26571 6512 26580
rect 6460 26537 6469 26571
rect 6469 26537 6503 26571
rect 6503 26537 6512 26571
rect 6460 26528 6512 26537
rect 6736 26528 6788 26580
rect 7380 26571 7432 26580
rect 7380 26537 7389 26571
rect 7389 26537 7423 26571
rect 7423 26537 7432 26571
rect 7380 26528 7432 26537
rect 7472 26528 7524 26580
rect 8116 26528 8168 26580
rect 14004 26528 14056 26580
rect 15476 26571 15528 26580
rect 15476 26537 15485 26571
rect 15485 26537 15519 26571
rect 15519 26537 15528 26571
rect 15476 26528 15528 26537
rect 6368 26392 6420 26444
rect 7012 26460 7064 26512
rect 7104 26460 7156 26512
rect 12716 26460 12768 26512
rect 6920 26435 6972 26444
rect 6920 26401 6930 26435
rect 6930 26401 6964 26435
rect 6964 26401 6972 26435
rect 6920 26392 6972 26401
rect 8392 26435 8444 26444
rect 5724 26367 5776 26376
rect 5724 26333 5733 26367
rect 5733 26333 5767 26367
rect 5767 26333 5776 26367
rect 5724 26324 5776 26333
rect 4068 26256 4120 26308
rect 5908 26299 5960 26308
rect 5908 26265 5917 26299
rect 5917 26265 5951 26299
rect 5951 26265 5960 26299
rect 5908 26256 5960 26265
rect 1492 26231 1544 26240
rect 1492 26197 1501 26231
rect 1501 26197 1535 26231
rect 1535 26197 1544 26231
rect 1492 26188 1544 26197
rect 2780 26188 2832 26240
rect 6000 26231 6052 26240
rect 6000 26197 6009 26231
rect 6009 26197 6043 26231
rect 6043 26197 6052 26231
rect 6000 26188 6052 26197
rect 6276 26367 6328 26376
rect 6276 26333 6285 26367
rect 6285 26333 6319 26367
rect 6319 26333 6328 26367
rect 6276 26324 6328 26333
rect 6552 26324 6604 26376
rect 6368 26256 6420 26308
rect 7472 26367 7524 26376
rect 7472 26333 7481 26367
rect 7481 26333 7515 26367
rect 7515 26333 7524 26367
rect 7472 26324 7524 26333
rect 8392 26401 8401 26435
rect 8401 26401 8435 26435
rect 8435 26401 8444 26435
rect 8392 26392 8444 26401
rect 9404 26392 9456 26444
rect 14096 26435 14148 26444
rect 7196 26256 7248 26308
rect 8576 26367 8628 26376
rect 8576 26333 8585 26367
rect 8585 26333 8619 26367
rect 8619 26333 8628 26367
rect 8576 26324 8628 26333
rect 6644 26188 6696 26240
rect 8208 26256 8260 26308
rect 10600 26324 10652 26376
rect 10876 26324 10928 26376
rect 11612 26324 11664 26376
rect 14096 26401 14105 26435
rect 14105 26401 14139 26435
rect 14139 26401 14148 26435
rect 14096 26392 14148 26401
rect 16488 26571 16540 26580
rect 16488 26537 16497 26571
rect 16497 26537 16531 26571
rect 16531 26537 16540 26571
rect 16488 26528 16540 26537
rect 16672 26571 16724 26580
rect 16672 26537 16681 26571
rect 16681 26537 16715 26571
rect 16715 26537 16724 26571
rect 16672 26528 16724 26537
rect 17132 26528 17184 26580
rect 18512 26528 18564 26580
rect 16580 26460 16632 26512
rect 11244 26256 11296 26308
rect 13268 26324 13320 26376
rect 14188 26324 14240 26376
rect 15108 26324 15160 26376
rect 15936 26367 15988 26376
rect 15936 26333 15945 26367
rect 15945 26333 15979 26367
rect 15979 26333 15988 26367
rect 15936 26324 15988 26333
rect 17592 26324 17644 26376
rect 18604 26324 18656 26376
rect 20996 26392 21048 26444
rect 20076 26324 20128 26376
rect 9404 26188 9456 26240
rect 12992 26256 13044 26308
rect 13544 26299 13596 26308
rect 13544 26265 13553 26299
rect 13553 26265 13587 26299
rect 13587 26265 13596 26299
rect 13544 26256 13596 26265
rect 12440 26188 12492 26240
rect 13268 26188 13320 26240
rect 13728 26231 13780 26240
rect 16856 26299 16908 26308
rect 16856 26265 16865 26299
rect 16865 26265 16899 26299
rect 16899 26265 16908 26299
rect 16856 26256 16908 26265
rect 16948 26299 17000 26308
rect 16948 26265 16957 26299
rect 16957 26265 16991 26299
rect 16991 26265 17000 26299
rect 16948 26256 17000 26265
rect 13728 26197 13753 26231
rect 13753 26197 13780 26231
rect 13728 26188 13780 26197
rect 16580 26188 16632 26240
rect 17040 26231 17092 26240
rect 17040 26197 17049 26231
rect 17049 26197 17083 26231
rect 17083 26197 17092 26231
rect 17040 26188 17092 26197
rect 17224 26299 17276 26308
rect 17224 26265 17233 26299
rect 17233 26265 17267 26299
rect 17267 26265 17276 26299
rect 17224 26256 17276 26265
rect 18144 26256 18196 26308
rect 4874 26086 4926 26138
rect 4938 26086 4990 26138
rect 5002 26086 5054 26138
rect 5066 26086 5118 26138
rect 5130 26086 5182 26138
rect 2596 25984 2648 26036
rect 1860 25891 1912 25900
rect 1860 25857 1869 25891
rect 1869 25857 1903 25891
rect 1903 25857 1912 25891
rect 1860 25848 1912 25857
rect 2780 25916 2832 25968
rect 3608 25916 3660 25968
rect 2504 25848 2556 25900
rect 2964 25848 3016 25900
rect 3240 25780 3292 25832
rect 3424 25891 3476 25900
rect 3424 25857 3433 25891
rect 3433 25857 3467 25891
rect 3467 25857 3476 25891
rect 3424 25848 3476 25857
rect 3884 25984 3936 26036
rect 4068 26027 4120 26036
rect 4068 25993 4077 26027
rect 4077 25993 4111 26027
rect 4111 25993 4120 26027
rect 4068 25984 4120 25993
rect 3976 25916 4028 25968
rect 4988 25984 5040 26036
rect 5540 26027 5592 26036
rect 5540 25993 5549 26027
rect 5549 25993 5583 26027
rect 5583 25993 5592 26027
rect 5540 25984 5592 25993
rect 5908 25984 5960 26036
rect 6736 26027 6788 26036
rect 6736 25993 6745 26027
rect 6745 25993 6779 26027
rect 6779 25993 6788 26027
rect 6736 25984 6788 25993
rect 7196 26027 7248 26036
rect 7196 25993 7205 26027
rect 7205 25993 7239 26027
rect 7239 25993 7248 26027
rect 7196 25984 7248 25993
rect 4068 25848 4120 25900
rect 4436 25916 4488 25968
rect 4712 25916 4764 25968
rect 4620 25848 4672 25900
rect 5356 25916 5408 25968
rect 6460 25916 6512 25968
rect 6276 25848 6328 25900
rect 6552 25891 6604 25900
rect 6552 25857 6561 25891
rect 6561 25857 6595 25891
rect 6595 25857 6604 25891
rect 6552 25848 6604 25857
rect 7012 25916 7064 25968
rect 9496 25984 9548 26036
rect 11244 26027 11296 26036
rect 11244 25993 11253 26027
rect 11253 25993 11287 26027
rect 11287 25993 11296 26027
rect 11244 25984 11296 25993
rect 13084 25984 13136 26036
rect 13452 25984 13504 26036
rect 13728 26027 13780 26036
rect 13728 25993 13737 26027
rect 13737 25993 13771 26027
rect 13771 25993 13780 26027
rect 13728 25984 13780 25993
rect 14096 26027 14148 26036
rect 14096 25993 14105 26027
rect 14105 25993 14139 26027
rect 14139 25993 14148 26027
rect 14096 25984 14148 25993
rect 14188 25984 14240 26036
rect 16120 26027 16172 26036
rect 16120 25993 16129 26027
rect 16129 25993 16163 26027
rect 16163 25993 16172 26027
rect 16120 25984 16172 25993
rect 17500 26027 17552 26036
rect 17500 25993 17509 26027
rect 17509 25993 17543 26027
rect 17543 25993 17552 26027
rect 17500 25984 17552 25993
rect 21088 26027 21140 26036
rect 21088 25993 21097 26027
rect 21097 25993 21131 26027
rect 21131 25993 21140 26027
rect 21088 25984 21140 25993
rect 13268 25916 13320 25968
rect 13820 25916 13872 25968
rect 15476 25959 15528 25968
rect 15476 25925 15485 25959
rect 15485 25925 15519 25959
rect 15519 25925 15528 25959
rect 15476 25916 15528 25925
rect 16028 25916 16080 25968
rect 17224 25916 17276 25968
rect 20536 25916 20588 25968
rect 20904 25959 20956 25968
rect 20904 25925 20929 25959
rect 20929 25925 20956 25959
rect 20904 25916 20956 25925
rect 3884 25712 3936 25764
rect 4620 25712 4672 25764
rect 4804 25780 4856 25832
rect 6000 25780 6052 25832
rect 7196 25848 7248 25900
rect 8208 25891 8260 25900
rect 8208 25857 8217 25891
rect 8217 25857 8251 25891
rect 8251 25857 8260 25891
rect 8208 25848 8260 25857
rect 8392 25848 8444 25900
rect 8576 25848 8628 25900
rect 8760 25891 8812 25900
rect 8760 25857 8769 25891
rect 8769 25857 8803 25891
rect 8803 25857 8812 25891
rect 8760 25848 8812 25857
rect 9404 25848 9456 25900
rect 9588 25891 9640 25900
rect 9588 25857 9597 25891
rect 9597 25857 9631 25891
rect 9631 25857 9640 25891
rect 9588 25848 9640 25857
rect 10968 25848 11020 25900
rect 12716 25891 12768 25900
rect 12716 25857 12725 25891
rect 12725 25857 12759 25891
rect 12759 25857 12768 25891
rect 12716 25848 12768 25857
rect 13544 25891 13596 25900
rect 13544 25857 13553 25891
rect 13553 25857 13587 25891
rect 13587 25857 13596 25891
rect 13544 25848 13596 25857
rect 13636 25891 13688 25900
rect 13636 25857 13645 25891
rect 13645 25857 13679 25891
rect 13679 25857 13688 25891
rect 13636 25848 13688 25857
rect 14372 25848 14424 25900
rect 14556 25891 14608 25900
rect 14556 25857 14565 25891
rect 14565 25857 14599 25891
rect 14599 25857 14608 25891
rect 14556 25848 14608 25857
rect 15752 25891 15804 25900
rect 15752 25857 15761 25891
rect 15761 25857 15795 25891
rect 15795 25857 15804 25891
rect 15752 25848 15804 25857
rect 5264 25712 5316 25764
rect 6184 25712 6236 25764
rect 6552 25712 6604 25764
rect 7472 25712 7524 25764
rect 8300 25712 8352 25764
rect 13084 25780 13136 25832
rect 13360 25780 13412 25832
rect 16856 25848 16908 25900
rect 17316 25891 17368 25900
rect 17316 25857 17325 25891
rect 17325 25857 17359 25891
rect 17359 25857 17368 25891
rect 17316 25848 17368 25857
rect 16488 25780 16540 25832
rect 17224 25823 17276 25832
rect 17224 25789 17233 25823
rect 17233 25789 17267 25823
rect 17267 25789 17276 25823
rect 17224 25780 17276 25789
rect 1768 25644 1820 25696
rect 3700 25687 3752 25696
rect 3700 25653 3709 25687
rect 3709 25653 3743 25687
rect 3743 25653 3752 25687
rect 3700 25644 3752 25653
rect 4896 25644 4948 25696
rect 7380 25687 7432 25696
rect 7380 25653 7389 25687
rect 7389 25653 7423 25687
rect 7423 25653 7432 25687
rect 7380 25644 7432 25653
rect 8024 25644 8076 25696
rect 12992 25687 13044 25696
rect 12992 25653 13001 25687
rect 13001 25653 13035 25687
rect 13035 25653 13044 25687
rect 12992 25644 13044 25653
rect 13176 25644 13228 25696
rect 13452 25687 13504 25696
rect 13452 25653 13461 25687
rect 13461 25653 13495 25687
rect 13495 25653 13504 25687
rect 13452 25644 13504 25653
rect 16948 25644 17000 25696
rect 19984 25823 20036 25832
rect 19984 25789 19993 25823
rect 19993 25789 20027 25823
rect 20027 25789 20036 25823
rect 19984 25780 20036 25789
rect 19340 25644 19392 25696
rect 20812 25644 20864 25696
rect 20996 25644 21048 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 3976 25440 4028 25492
rect 4712 25440 4764 25492
rect 5356 25440 5408 25492
rect 848 25372 900 25424
rect 4344 25372 4396 25424
rect 1768 25279 1820 25288
rect 1768 25245 1777 25279
rect 1777 25245 1811 25279
rect 1811 25245 1820 25279
rect 1768 25236 1820 25245
rect 3700 25236 3752 25288
rect 3792 25168 3844 25220
rect 4068 25236 4120 25288
rect 4896 25279 4948 25288
rect 4896 25245 4905 25279
rect 4905 25245 4939 25279
rect 4939 25245 4948 25279
rect 4896 25236 4948 25245
rect 4988 25279 5040 25288
rect 4988 25245 4997 25279
rect 4997 25245 5031 25279
rect 5031 25245 5040 25279
rect 4988 25236 5040 25245
rect 5448 25236 5500 25288
rect 5632 25279 5684 25288
rect 5632 25245 5641 25279
rect 5641 25245 5675 25279
rect 5675 25245 5684 25279
rect 5632 25236 5684 25245
rect 5908 25440 5960 25492
rect 6184 25440 6236 25492
rect 7380 25372 7432 25424
rect 7564 25372 7616 25424
rect 8760 25372 8812 25424
rect 6736 25347 6788 25356
rect 5816 25236 5868 25288
rect 6736 25313 6745 25347
rect 6745 25313 6779 25347
rect 6779 25313 6788 25347
rect 6736 25304 6788 25313
rect 6828 25347 6880 25356
rect 6828 25313 6837 25347
rect 6837 25313 6871 25347
rect 6871 25313 6880 25347
rect 6828 25304 6880 25313
rect 7288 25347 7340 25356
rect 7288 25313 7297 25347
rect 7297 25313 7331 25347
rect 7331 25313 7340 25347
rect 7288 25304 7340 25313
rect 7472 25304 7524 25356
rect 7748 25304 7800 25356
rect 8300 25304 8352 25356
rect 9588 25304 9640 25356
rect 11612 25304 11664 25356
rect 13268 25440 13320 25492
rect 15936 25440 15988 25492
rect 19984 25440 20036 25492
rect 20904 25440 20956 25492
rect 18604 25304 18656 25356
rect 6184 25236 6236 25288
rect 6920 25236 6972 25288
rect 8208 25236 8260 25288
rect 10048 25236 10100 25288
rect 14556 25236 14608 25288
rect 14924 25236 14976 25288
rect 4712 25100 4764 25152
rect 5356 25100 5408 25152
rect 10968 25168 11020 25220
rect 12440 25168 12492 25220
rect 6736 25100 6788 25152
rect 7932 25143 7984 25152
rect 7932 25109 7941 25143
rect 7941 25109 7975 25143
rect 7975 25109 7984 25143
rect 7932 25100 7984 25109
rect 8300 25100 8352 25152
rect 8484 25100 8536 25152
rect 9312 25100 9364 25152
rect 10508 25100 10560 25152
rect 12624 25100 12676 25152
rect 13544 25100 13596 25152
rect 15476 25143 15528 25152
rect 15476 25109 15485 25143
rect 15485 25109 15519 25143
rect 15519 25109 15528 25143
rect 15476 25100 15528 25109
rect 19340 25279 19392 25288
rect 19340 25245 19349 25279
rect 19349 25245 19383 25279
rect 19383 25245 19392 25279
rect 19340 25236 19392 25245
rect 16488 25211 16540 25220
rect 16488 25177 16497 25211
rect 16497 25177 16531 25211
rect 16531 25177 16540 25211
rect 16488 25168 16540 25177
rect 20996 25168 21048 25220
rect 16672 25100 16724 25152
rect 20536 25100 20588 25152
rect 4874 24998 4926 25050
rect 4938 24998 4990 25050
rect 5002 24998 5054 25050
rect 5066 24998 5118 25050
rect 5130 24998 5182 25050
rect 1952 24828 2004 24880
rect 6460 24896 6512 24948
rect 6828 24896 6880 24948
rect 2872 24871 2924 24880
rect 2872 24837 2899 24871
rect 2899 24837 2924 24871
rect 2872 24828 2924 24837
rect 3148 24828 3200 24880
rect 3700 24828 3752 24880
rect 2964 24760 3016 24812
rect 8116 24828 8168 24880
rect 4528 24760 4580 24812
rect 848 24624 900 24676
rect 2044 24599 2096 24608
rect 2044 24565 2053 24599
rect 2053 24565 2087 24599
rect 2087 24565 2096 24599
rect 2044 24556 2096 24565
rect 2228 24556 2280 24608
rect 4344 24735 4396 24744
rect 4344 24701 4353 24735
rect 4353 24701 4387 24735
rect 4387 24701 4396 24735
rect 4344 24692 4396 24701
rect 5356 24803 5408 24812
rect 5356 24769 5365 24803
rect 5365 24769 5399 24803
rect 5399 24769 5408 24803
rect 5356 24760 5408 24769
rect 4712 24692 4764 24744
rect 5448 24692 5500 24744
rect 5816 24803 5868 24812
rect 5816 24769 5825 24803
rect 5825 24769 5859 24803
rect 5859 24769 5868 24803
rect 5816 24760 5868 24769
rect 6276 24760 6328 24812
rect 6368 24803 6420 24812
rect 6368 24769 6377 24803
rect 6377 24769 6411 24803
rect 6411 24769 6420 24803
rect 6368 24760 6420 24769
rect 6552 24803 6604 24812
rect 6552 24769 6561 24803
rect 6561 24769 6595 24803
rect 6595 24769 6604 24803
rect 6552 24760 6604 24769
rect 6736 24803 6788 24812
rect 6736 24769 6745 24803
rect 6745 24769 6779 24803
rect 6779 24769 6788 24803
rect 6736 24760 6788 24769
rect 6828 24803 6880 24812
rect 6828 24769 6837 24803
rect 6837 24769 6871 24803
rect 6871 24769 6880 24803
rect 6828 24760 6880 24769
rect 6920 24803 6972 24812
rect 6920 24769 6929 24803
rect 6929 24769 6963 24803
rect 6963 24769 6972 24803
rect 6920 24760 6972 24769
rect 7380 24760 7432 24812
rect 7564 24803 7616 24812
rect 7564 24769 7573 24803
rect 7573 24769 7607 24803
rect 7607 24769 7616 24803
rect 7564 24760 7616 24769
rect 7748 24760 7800 24812
rect 8024 24803 8076 24812
rect 8024 24769 8033 24803
rect 8033 24769 8067 24803
rect 8067 24769 8076 24803
rect 8024 24760 8076 24769
rect 4804 24624 4856 24676
rect 5264 24624 5316 24676
rect 5816 24624 5868 24676
rect 6552 24624 6604 24676
rect 6828 24624 6880 24676
rect 15936 24896 15988 24948
rect 20536 24896 20588 24948
rect 8392 24803 8444 24812
rect 8392 24769 8401 24803
rect 8401 24769 8435 24803
rect 8435 24769 8444 24803
rect 8392 24760 8444 24769
rect 9956 24760 10008 24812
rect 10324 24760 10376 24812
rect 10508 24760 10560 24812
rect 10048 24735 10100 24744
rect 10048 24701 10057 24735
rect 10057 24701 10091 24735
rect 10091 24701 10100 24735
rect 10048 24692 10100 24701
rect 10784 24692 10836 24744
rect 11612 24692 11664 24744
rect 12348 24692 12400 24744
rect 15016 24760 15068 24812
rect 15384 24803 15436 24812
rect 15384 24769 15418 24803
rect 15418 24769 15436 24803
rect 15384 24760 15436 24769
rect 16856 24760 16908 24812
rect 18604 24803 18656 24812
rect 18604 24769 18613 24803
rect 18613 24769 18647 24803
rect 18647 24769 18656 24803
rect 18604 24760 18656 24769
rect 18696 24760 18748 24812
rect 20536 24760 20588 24812
rect 16488 24624 16540 24676
rect 3424 24556 3476 24608
rect 3976 24556 4028 24608
rect 7104 24599 7156 24608
rect 7104 24565 7113 24599
rect 7113 24565 7147 24599
rect 7147 24565 7156 24599
rect 7104 24556 7156 24565
rect 8392 24556 8444 24608
rect 10416 24556 10468 24608
rect 12072 24556 12124 24608
rect 20076 24599 20128 24608
rect 20076 24565 20085 24599
rect 20085 24565 20119 24599
rect 20119 24565 20128 24599
rect 20076 24556 20128 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 2964 24395 3016 24404
rect 2964 24361 2973 24395
rect 2973 24361 3007 24395
rect 3007 24361 3016 24395
rect 2964 24352 3016 24361
rect 3424 24395 3476 24404
rect 3424 24361 3433 24395
rect 3433 24361 3467 24395
rect 3467 24361 3476 24395
rect 3424 24352 3476 24361
rect 7840 24352 7892 24404
rect 3148 24284 3200 24336
rect 5448 24284 5500 24336
rect 1400 24259 1452 24268
rect 1400 24225 1409 24259
rect 1409 24225 1443 24259
rect 1443 24225 1452 24259
rect 1400 24216 1452 24225
rect 2044 24148 2096 24200
rect 2780 24148 2832 24200
rect 6368 24259 6420 24268
rect 6368 24225 6377 24259
rect 6377 24225 6411 24259
rect 6411 24225 6420 24259
rect 6368 24216 6420 24225
rect 6460 24259 6512 24268
rect 6460 24225 6469 24259
rect 6469 24225 6503 24259
rect 6503 24225 6512 24259
rect 6460 24216 6512 24225
rect 3240 24148 3292 24200
rect 6736 24148 6788 24200
rect 6828 24191 6880 24200
rect 6828 24157 6837 24191
rect 6837 24157 6871 24191
rect 6871 24157 6880 24191
rect 6828 24148 6880 24157
rect 6920 24148 6972 24200
rect 8300 24395 8352 24404
rect 8300 24361 8309 24395
rect 8309 24361 8343 24395
rect 8343 24361 8352 24395
rect 8300 24352 8352 24361
rect 12440 24395 12492 24404
rect 12440 24361 12449 24395
rect 12449 24361 12483 24395
rect 12483 24361 12492 24395
rect 12440 24352 12492 24361
rect 16856 24395 16908 24404
rect 16856 24361 16865 24395
rect 16865 24361 16899 24395
rect 16899 24361 16908 24395
rect 16856 24352 16908 24361
rect 18696 24395 18748 24404
rect 18696 24361 18705 24395
rect 18705 24361 18739 24395
rect 18739 24361 18748 24395
rect 18696 24352 18748 24361
rect 20812 24352 20864 24404
rect 16488 24284 16540 24336
rect 8116 24216 8168 24268
rect 8300 24191 8352 24200
rect 8300 24157 8309 24191
rect 8309 24157 8343 24191
rect 8343 24157 8352 24191
rect 8300 24148 8352 24157
rect 12348 24259 12400 24268
rect 12348 24225 12357 24259
rect 12357 24225 12391 24259
rect 12391 24225 12400 24259
rect 12348 24216 12400 24225
rect 8852 24148 8904 24200
rect 3056 24012 3108 24064
rect 3976 24012 4028 24064
rect 7104 24080 7156 24132
rect 8944 24123 8996 24132
rect 8944 24089 8953 24123
rect 8953 24089 8987 24123
rect 8987 24089 8996 24123
rect 8944 24080 8996 24089
rect 12072 24191 12124 24200
rect 12072 24157 12090 24191
rect 12090 24157 12124 24191
rect 12072 24148 12124 24157
rect 12624 24191 12676 24200
rect 12624 24157 12633 24191
rect 12633 24157 12667 24191
rect 12667 24157 12676 24191
rect 12624 24148 12676 24157
rect 13452 24216 13504 24268
rect 16672 24216 16724 24268
rect 18604 24216 18656 24268
rect 19248 24216 19300 24268
rect 12808 24191 12860 24200
rect 12808 24157 12817 24191
rect 12817 24157 12851 24191
rect 12851 24157 12860 24191
rect 12808 24148 12860 24157
rect 12992 24191 13044 24200
rect 12992 24157 13001 24191
rect 13001 24157 13035 24191
rect 13035 24157 13044 24191
rect 12992 24148 13044 24157
rect 13084 24191 13136 24200
rect 13084 24157 13093 24191
rect 13093 24157 13127 24191
rect 13127 24157 13136 24191
rect 13084 24148 13136 24157
rect 13820 24148 13872 24200
rect 15200 24148 15252 24200
rect 13176 24080 13228 24132
rect 14648 24080 14700 24132
rect 6184 24055 6236 24064
rect 6184 24021 6193 24055
rect 6193 24021 6227 24055
rect 6227 24021 6236 24055
rect 6184 24012 6236 24021
rect 7196 24012 7248 24064
rect 9404 24012 9456 24064
rect 10048 24012 10100 24064
rect 12072 24012 12124 24064
rect 12900 24055 12952 24064
rect 12900 24021 12909 24055
rect 12909 24021 12943 24055
rect 12943 24021 12952 24055
rect 12900 24012 12952 24021
rect 13360 24055 13412 24064
rect 13360 24021 13369 24055
rect 13369 24021 13403 24055
rect 13403 24021 13412 24055
rect 13360 24012 13412 24021
rect 15108 24012 15160 24064
rect 19800 24080 19852 24132
rect 20076 24080 20128 24132
rect 15568 24055 15620 24064
rect 15568 24021 15577 24055
rect 15577 24021 15611 24055
rect 15611 24021 15620 24055
rect 15568 24012 15620 24021
rect 21180 24055 21232 24064
rect 21180 24021 21189 24055
rect 21189 24021 21223 24055
rect 21223 24021 21232 24055
rect 21180 24012 21232 24021
rect 4874 23910 4926 23962
rect 4938 23910 4990 23962
rect 5002 23910 5054 23962
rect 5066 23910 5118 23962
rect 5130 23910 5182 23962
rect 1216 23808 1268 23860
rect 2780 23851 2832 23860
rect 2228 23740 2280 23792
rect 1952 23715 2004 23724
rect 1952 23681 1961 23715
rect 1961 23681 1995 23715
rect 1995 23681 2004 23715
rect 1952 23672 2004 23681
rect 2780 23817 2789 23851
rect 2789 23817 2823 23851
rect 2823 23817 2832 23851
rect 2780 23808 2832 23817
rect 3240 23808 3292 23860
rect 5816 23808 5868 23860
rect 7196 23851 7248 23860
rect 7196 23817 7205 23851
rect 7205 23817 7239 23851
rect 7239 23817 7248 23851
rect 7196 23808 7248 23817
rect 10416 23808 10468 23860
rect 9956 23740 10008 23792
rect 2872 23672 2924 23724
rect 2964 23715 3016 23724
rect 2964 23681 2973 23715
rect 2973 23681 3007 23715
rect 3007 23681 3016 23715
rect 2964 23672 3016 23681
rect 3976 23672 4028 23724
rect 6920 23672 6972 23724
rect 10324 23672 10376 23724
rect 3424 23604 3476 23656
rect 4804 23604 4856 23656
rect 7380 23604 7432 23656
rect 10416 23647 10468 23656
rect 10416 23613 10425 23647
rect 10425 23613 10459 23647
rect 10459 23613 10468 23647
rect 10416 23604 10468 23613
rect 7104 23536 7156 23588
rect 8392 23579 8444 23588
rect 8392 23545 8401 23579
rect 8401 23545 8435 23579
rect 8435 23545 8444 23579
rect 8392 23536 8444 23545
rect 10968 23715 11020 23724
rect 10968 23681 10977 23715
rect 10977 23681 11011 23715
rect 11011 23681 11020 23715
rect 10968 23672 11020 23681
rect 14648 23851 14700 23860
rect 14648 23817 14657 23851
rect 14657 23817 14691 23851
rect 14691 23817 14700 23851
rect 14648 23808 14700 23817
rect 15292 23851 15344 23860
rect 15292 23817 15301 23851
rect 15301 23817 15335 23851
rect 15335 23817 15344 23851
rect 15292 23808 15344 23817
rect 15476 23851 15528 23860
rect 15476 23817 15503 23851
rect 15503 23817 15528 23851
rect 15476 23808 15528 23817
rect 16488 23808 16540 23860
rect 12900 23740 12952 23792
rect 13360 23740 13412 23792
rect 12072 23715 12124 23724
rect 12072 23681 12081 23715
rect 12081 23681 12115 23715
rect 12115 23681 12124 23715
rect 12072 23672 12124 23681
rect 13084 23672 13136 23724
rect 12440 23647 12492 23656
rect 12440 23613 12449 23647
rect 12449 23613 12483 23647
rect 12483 23613 12492 23647
rect 12440 23604 12492 23613
rect 14924 23672 14976 23724
rect 15568 23672 15620 23724
rect 15936 23715 15988 23724
rect 15936 23681 15945 23715
rect 15945 23681 15979 23715
rect 15979 23681 15988 23715
rect 15936 23672 15988 23681
rect 16672 23672 16724 23724
rect 20076 23740 20128 23792
rect 21180 23672 21232 23724
rect 19800 23647 19852 23656
rect 19800 23613 19809 23647
rect 19809 23613 19843 23647
rect 19843 23613 19852 23647
rect 19800 23604 19852 23613
rect 13820 23579 13872 23588
rect 13820 23545 13829 23579
rect 13829 23545 13863 23579
rect 13863 23545 13872 23579
rect 13820 23536 13872 23545
rect 1676 23468 1728 23520
rect 6184 23468 6236 23520
rect 7748 23468 7800 23520
rect 10784 23511 10836 23520
rect 10784 23477 10793 23511
rect 10793 23477 10827 23511
rect 10827 23477 10836 23511
rect 10784 23468 10836 23477
rect 14004 23468 14056 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 2872 23264 2924 23316
rect 3976 23307 4028 23316
rect 3976 23273 3985 23307
rect 3985 23273 4019 23307
rect 4019 23273 4028 23307
rect 3976 23264 4028 23273
rect 12808 23307 12860 23316
rect 12808 23273 12817 23307
rect 12817 23273 12851 23307
rect 12851 23273 12860 23307
rect 12808 23264 12860 23273
rect 12992 23264 13044 23316
rect 20904 23264 20956 23316
rect 20260 23196 20312 23248
rect 3056 23128 3108 23180
rect 10140 23128 10192 23180
rect 3240 23103 3292 23112
rect 3240 23069 3249 23103
rect 3249 23069 3283 23103
rect 3283 23069 3292 23103
rect 3240 23060 3292 23069
rect 3424 23060 3476 23112
rect 4804 23060 4856 23112
rect 6828 23060 6880 23112
rect 7288 22992 7340 23044
rect 8392 23060 8444 23112
rect 8668 23060 8720 23112
rect 9312 23060 9364 23112
rect 9772 23103 9824 23112
rect 9772 23069 9781 23103
rect 9781 23069 9815 23103
rect 9815 23069 9824 23103
rect 9772 23060 9824 23069
rect 10784 23060 10836 23112
rect 12624 23060 12676 23112
rect 2688 22967 2740 22976
rect 2688 22933 2697 22967
rect 2697 22933 2731 22967
rect 2731 22933 2740 22967
rect 2688 22924 2740 22933
rect 9036 22967 9088 22976
rect 9036 22933 9045 22967
rect 9045 22933 9079 22967
rect 9079 22933 9088 22967
rect 9036 22924 9088 22933
rect 9220 22924 9272 22976
rect 12716 22924 12768 22976
rect 13176 23128 13228 23180
rect 13912 23171 13964 23180
rect 13912 23137 13921 23171
rect 13921 23137 13955 23171
rect 13955 23137 13964 23171
rect 13912 23128 13964 23137
rect 19248 23171 19300 23180
rect 19248 23137 19257 23171
rect 19257 23137 19291 23171
rect 19291 23137 19300 23171
rect 19248 23128 19300 23137
rect 20812 23171 20864 23180
rect 20812 23137 20821 23171
rect 20821 23137 20855 23171
rect 20855 23137 20864 23171
rect 20812 23128 20864 23137
rect 14648 23103 14700 23112
rect 14648 23069 14657 23103
rect 14657 23069 14691 23103
rect 14691 23069 14700 23103
rect 14648 23060 14700 23069
rect 15016 23060 15068 23112
rect 16672 23060 16724 23112
rect 20720 23060 20772 23112
rect 13820 22992 13872 23044
rect 17316 22992 17368 23044
rect 18972 22992 19024 23044
rect 14004 22924 14056 22976
rect 18788 22967 18840 22976
rect 18788 22933 18797 22967
rect 18797 22933 18831 22967
rect 18831 22933 18840 22967
rect 18788 22924 18840 22933
rect 21272 22967 21324 22976
rect 21272 22933 21281 22967
rect 21281 22933 21315 22967
rect 21315 22933 21324 22967
rect 21272 22924 21324 22933
rect 4874 22822 4926 22874
rect 4938 22822 4990 22874
rect 5002 22822 5054 22874
rect 5066 22822 5118 22874
rect 5130 22822 5182 22874
rect 6920 22720 6972 22772
rect 8576 22720 8628 22772
rect 2688 22652 2740 22704
rect 10784 22763 10836 22772
rect 10784 22729 10793 22763
rect 10793 22729 10827 22763
rect 10827 22729 10836 22763
rect 10784 22720 10836 22729
rect 10324 22652 10376 22704
rect 10968 22652 11020 22704
rect 12072 22720 12124 22772
rect 14648 22720 14700 22772
rect 1400 22584 1452 22636
rect 2320 22584 2372 22636
rect 5448 22584 5500 22636
rect 6828 22584 6880 22636
rect 7656 22627 7708 22636
rect 7656 22593 7690 22627
rect 7690 22593 7708 22627
rect 7656 22584 7708 22593
rect 9404 22627 9456 22636
rect 9404 22593 9413 22627
rect 9413 22593 9447 22627
rect 9447 22593 9456 22627
rect 9404 22584 9456 22593
rect 4804 22559 4856 22568
rect 4804 22525 4813 22559
rect 4813 22525 4847 22559
rect 4847 22525 4856 22559
rect 4804 22516 4856 22525
rect 4712 22448 4764 22500
rect 6736 22516 6788 22568
rect 7288 22516 7340 22568
rect 7380 22559 7432 22568
rect 7380 22525 7389 22559
rect 7389 22525 7423 22559
rect 7423 22525 7432 22559
rect 7380 22516 7432 22525
rect 9956 22584 10008 22636
rect 10968 22516 11020 22568
rect 11244 22584 11296 22636
rect 13912 22652 13964 22704
rect 16212 22720 16264 22772
rect 18972 22763 19024 22772
rect 18972 22729 18981 22763
rect 18981 22729 19015 22763
rect 19015 22729 19024 22763
rect 18972 22720 19024 22729
rect 21272 22763 21324 22772
rect 21272 22729 21281 22763
rect 21281 22729 21315 22763
rect 21315 22729 21324 22763
rect 21272 22720 21324 22729
rect 17040 22652 17092 22704
rect 9220 22491 9272 22500
rect 9220 22457 9229 22491
rect 9229 22457 9263 22491
rect 9263 22457 9272 22491
rect 9220 22448 9272 22457
rect 10416 22448 10468 22500
rect 15844 22627 15896 22636
rect 15844 22593 15853 22627
rect 15853 22593 15887 22627
rect 15887 22593 15896 22627
rect 15844 22584 15896 22593
rect 16120 22627 16172 22636
rect 16120 22593 16129 22627
rect 16129 22593 16163 22627
rect 16163 22593 16172 22627
rect 16120 22584 16172 22593
rect 16304 22584 16356 22636
rect 16672 22627 16724 22636
rect 13636 22559 13688 22568
rect 13636 22525 13645 22559
rect 13645 22525 13679 22559
rect 13679 22525 13688 22559
rect 13636 22516 13688 22525
rect 16672 22593 16681 22627
rect 16681 22593 16715 22627
rect 16715 22593 16724 22627
rect 16672 22584 16724 22593
rect 18696 22584 18748 22636
rect 19340 22627 19392 22636
rect 19340 22593 19349 22627
rect 19349 22593 19383 22627
rect 19383 22593 19392 22627
rect 19340 22584 19392 22593
rect 18144 22516 18196 22568
rect 18788 22559 18840 22568
rect 18788 22525 18797 22559
rect 18797 22525 18831 22559
rect 18831 22525 18840 22559
rect 18788 22516 18840 22525
rect 20260 22559 20312 22568
rect 20260 22525 20269 22559
rect 20269 22525 20303 22559
rect 20303 22525 20312 22559
rect 20260 22516 20312 22525
rect 3884 22423 3936 22432
rect 3884 22389 3893 22423
rect 3893 22389 3927 22423
rect 3927 22389 3936 22423
rect 3884 22380 3936 22389
rect 8300 22380 8352 22432
rect 9036 22380 9088 22432
rect 10784 22380 10836 22432
rect 12072 22423 12124 22432
rect 12072 22389 12081 22423
rect 12081 22389 12115 22423
rect 12115 22389 12124 22423
rect 12072 22380 12124 22389
rect 12164 22380 12216 22432
rect 14372 22448 14424 22500
rect 21364 22559 21416 22568
rect 21364 22525 21373 22559
rect 21373 22525 21407 22559
rect 21407 22525 21416 22559
rect 21364 22516 21416 22525
rect 22192 22627 22244 22636
rect 22192 22593 22201 22627
rect 22201 22593 22235 22627
rect 22235 22593 22244 22627
rect 22192 22584 22244 22593
rect 22100 22559 22152 22568
rect 22100 22525 22109 22559
rect 22109 22525 22143 22559
rect 22143 22525 22152 22559
rect 22100 22516 22152 22525
rect 12900 22380 12952 22432
rect 13084 22423 13136 22432
rect 13084 22389 13093 22423
rect 13093 22389 13127 22423
rect 13127 22389 13136 22423
rect 13084 22380 13136 22389
rect 16028 22380 16080 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 3240 22176 3292 22228
rect 1400 22083 1452 22092
rect 1400 22049 1409 22083
rect 1409 22049 1443 22083
rect 1443 22049 1452 22083
rect 1400 22040 1452 22049
rect 2412 22040 2464 22092
rect 4804 22176 4856 22228
rect 6920 22176 6972 22228
rect 7656 22176 7708 22228
rect 7012 22040 7064 22092
rect 1676 22015 1728 22024
rect 1676 21981 1710 22015
rect 1710 21981 1728 22015
rect 1676 21972 1728 21981
rect 3884 21972 3936 22024
rect 7196 21972 7248 22024
rect 9772 22108 9824 22160
rect 10968 22108 11020 22160
rect 8208 21972 8260 22024
rect 8392 22015 8444 22024
rect 8392 21981 8401 22015
rect 8401 21981 8435 22015
rect 8435 21981 8444 22015
rect 8392 21972 8444 21981
rect 8484 22015 8536 22024
rect 8484 21981 8493 22015
rect 8493 21981 8527 22015
rect 8527 21981 8536 22015
rect 8484 21972 8536 21981
rect 9956 21972 10008 22024
rect 10784 21972 10836 22024
rect 12072 22108 12124 22160
rect 12532 22176 12584 22228
rect 13636 22219 13688 22228
rect 13636 22185 13645 22219
rect 13645 22185 13679 22219
rect 13679 22185 13688 22219
rect 13636 22176 13688 22185
rect 13728 22176 13780 22228
rect 16304 22176 16356 22228
rect 17316 22219 17368 22228
rect 17316 22185 17325 22219
rect 17325 22185 17359 22219
rect 17359 22185 17368 22219
rect 17316 22176 17368 22185
rect 7012 21947 7064 21956
rect 7012 21913 7021 21947
rect 7021 21913 7055 21947
rect 7055 21913 7064 21947
rect 7012 21904 7064 21913
rect 5264 21836 5316 21888
rect 6736 21836 6788 21888
rect 7748 21947 7800 21956
rect 7748 21913 7757 21947
rect 7757 21913 7791 21947
rect 7791 21913 7800 21947
rect 7748 21904 7800 21913
rect 9772 21904 9824 21956
rect 10416 21904 10468 21956
rect 8944 21836 8996 21888
rect 10140 21879 10192 21888
rect 10140 21845 10149 21879
rect 10149 21845 10183 21879
rect 10183 21845 10192 21879
rect 10140 21836 10192 21845
rect 11520 21879 11572 21888
rect 11520 21845 11529 21879
rect 11529 21845 11563 21879
rect 11563 21845 11572 21879
rect 11520 21836 11572 21845
rect 11704 21947 11756 21956
rect 11704 21913 11713 21947
rect 11713 21913 11747 21947
rect 11747 21913 11756 21947
rect 11704 21904 11756 21913
rect 12164 21972 12216 22024
rect 12072 21904 12124 21956
rect 12532 22040 12584 22092
rect 12348 21904 12400 21956
rect 12900 22108 12952 22160
rect 12992 22083 13044 22092
rect 12992 22049 13001 22083
rect 13001 22049 13035 22083
rect 13035 22049 13044 22083
rect 12992 22040 13044 22049
rect 13728 22040 13780 22092
rect 13360 22015 13412 22024
rect 13360 21981 13369 22015
rect 13369 21981 13403 22015
rect 13403 21981 13412 22015
rect 13360 21972 13412 21981
rect 13820 22015 13872 22024
rect 13820 21981 13829 22015
rect 13829 21981 13863 22015
rect 13863 21981 13872 22015
rect 16948 22108 17000 22160
rect 15476 22040 15528 22092
rect 18144 22040 18196 22092
rect 13820 21972 13872 21981
rect 14648 21972 14700 22024
rect 15568 22015 15620 22024
rect 15568 21981 15577 22015
rect 15577 21981 15611 22015
rect 15611 21981 15620 22015
rect 15568 21972 15620 21981
rect 16120 21972 16172 22024
rect 16672 21972 16724 22024
rect 17040 22015 17092 22024
rect 17040 21981 17049 22015
rect 17049 21981 17083 22015
rect 17083 21981 17092 22015
rect 17040 21972 17092 21981
rect 12624 21879 12676 21888
rect 12624 21845 12633 21879
rect 12633 21845 12667 21879
rect 12667 21845 12676 21879
rect 12624 21836 12676 21845
rect 12808 21947 12860 21956
rect 12808 21913 12817 21947
rect 12817 21913 12851 21947
rect 12851 21913 12860 21947
rect 12808 21904 12860 21913
rect 16212 21904 16264 21956
rect 16948 21947 17000 21956
rect 16948 21913 16957 21947
rect 16957 21913 16991 21947
rect 16991 21913 17000 21947
rect 16948 21904 17000 21913
rect 17592 22015 17644 22024
rect 17592 21981 17601 22015
rect 17601 21981 17635 22015
rect 17635 21981 17644 22015
rect 17592 21972 17644 21981
rect 17868 22015 17920 22024
rect 17868 21981 17877 22015
rect 17877 21981 17911 22015
rect 17911 21981 17920 22015
rect 17868 21972 17920 21981
rect 18420 21972 18472 22024
rect 18696 22015 18748 22024
rect 18696 21981 18705 22015
rect 18705 21981 18739 22015
rect 18739 21981 18748 22015
rect 18696 21972 18748 21981
rect 19248 22083 19300 22092
rect 19248 22049 19257 22083
rect 19257 22049 19291 22083
rect 19291 22049 19300 22083
rect 19248 22040 19300 22049
rect 19340 21972 19392 22024
rect 20996 22040 21048 22092
rect 22284 22040 22336 22092
rect 13176 21836 13228 21888
rect 13636 21836 13688 21888
rect 14924 21836 14976 21888
rect 15660 21879 15712 21888
rect 15660 21845 15669 21879
rect 15669 21845 15703 21879
rect 15703 21845 15712 21879
rect 15660 21836 15712 21845
rect 16304 21836 16356 21888
rect 16764 21836 16816 21888
rect 17316 21836 17368 21888
rect 17776 21879 17828 21888
rect 17776 21845 17785 21879
rect 17785 21845 17819 21879
rect 17819 21845 17828 21879
rect 17776 21836 17828 21845
rect 18052 21879 18104 21888
rect 18052 21845 18061 21879
rect 18061 21845 18095 21879
rect 18095 21845 18104 21879
rect 18052 21836 18104 21845
rect 18604 21947 18656 21956
rect 18604 21913 18613 21947
rect 18613 21913 18647 21947
rect 18647 21913 18656 21947
rect 18604 21904 18656 21913
rect 20168 21836 20220 21888
rect 20720 21836 20772 21888
rect 4874 21734 4926 21786
rect 4938 21734 4990 21786
rect 5002 21734 5054 21786
rect 5066 21734 5118 21786
rect 5130 21734 5182 21786
rect 5448 21675 5500 21684
rect 5448 21641 5457 21675
rect 5457 21641 5491 21675
rect 5491 21641 5500 21675
rect 5448 21632 5500 21641
rect 848 21496 900 21548
rect 2320 21539 2372 21548
rect 2320 21505 2329 21539
rect 2329 21505 2363 21539
rect 2363 21505 2372 21539
rect 2320 21496 2372 21505
rect 2872 21496 2924 21548
rect 5264 21564 5316 21616
rect 7104 21632 7156 21684
rect 7196 21675 7248 21684
rect 7196 21641 7205 21675
rect 7205 21641 7239 21675
rect 7239 21641 7248 21675
rect 7196 21632 7248 21641
rect 6920 21564 6972 21616
rect 4804 21428 4856 21480
rect 7104 21539 7156 21548
rect 7104 21505 7113 21539
rect 7113 21505 7147 21539
rect 7147 21505 7156 21539
rect 7104 21496 7156 21505
rect 7196 21496 7248 21548
rect 5264 21428 5316 21480
rect 5448 21360 5500 21412
rect 5724 21471 5776 21480
rect 5724 21437 5733 21471
rect 5733 21437 5767 21471
rect 5767 21437 5776 21471
rect 5724 21428 5776 21437
rect 6644 21360 6696 21412
rect 1584 21335 1636 21344
rect 1584 21301 1593 21335
rect 1593 21301 1627 21335
rect 1627 21301 1636 21335
rect 1584 21292 1636 21301
rect 4620 21292 4672 21344
rect 6920 21471 6972 21480
rect 6920 21437 6929 21471
rect 6929 21437 6963 21471
rect 6963 21437 6972 21471
rect 6920 21428 6972 21437
rect 7104 21360 7156 21412
rect 7472 21632 7524 21684
rect 7840 21632 7892 21684
rect 7932 21564 7984 21616
rect 7472 21539 7524 21548
rect 7472 21505 7481 21539
rect 7481 21505 7515 21539
rect 7515 21505 7524 21539
rect 7472 21496 7524 21505
rect 8024 21496 8076 21548
rect 13636 21632 13688 21684
rect 14648 21632 14700 21684
rect 15568 21632 15620 21684
rect 12164 21607 12216 21616
rect 12164 21573 12173 21607
rect 12173 21573 12207 21607
rect 12207 21573 12216 21607
rect 12164 21564 12216 21573
rect 11520 21496 11572 21548
rect 12256 21539 12308 21548
rect 12256 21505 12265 21539
rect 12265 21505 12299 21539
rect 12299 21505 12308 21539
rect 12256 21496 12308 21505
rect 8944 21360 8996 21412
rect 11888 21360 11940 21412
rect 7840 21292 7892 21344
rect 13360 21564 13412 21616
rect 12532 21539 12584 21548
rect 12532 21505 12541 21539
rect 12541 21505 12575 21539
rect 12575 21505 12584 21539
rect 12532 21496 12584 21505
rect 15292 21607 15344 21616
rect 15292 21573 15301 21607
rect 15301 21573 15335 21607
rect 15335 21573 15344 21607
rect 15292 21564 15344 21573
rect 15844 21675 15896 21684
rect 15844 21641 15853 21675
rect 15853 21641 15887 21675
rect 15887 21641 15896 21675
rect 15844 21632 15896 21641
rect 16672 21675 16724 21684
rect 16672 21641 16681 21675
rect 16681 21641 16715 21675
rect 16715 21641 16724 21675
rect 16672 21632 16724 21641
rect 16028 21564 16080 21616
rect 16396 21564 16448 21616
rect 14924 21496 14976 21548
rect 15384 21539 15436 21548
rect 15384 21505 15393 21539
rect 15393 21505 15427 21539
rect 15427 21505 15436 21539
rect 15384 21496 15436 21505
rect 15660 21496 15712 21548
rect 15844 21539 15896 21548
rect 15844 21505 15853 21539
rect 15853 21505 15887 21539
rect 15887 21505 15896 21539
rect 15844 21496 15896 21505
rect 16120 21539 16172 21548
rect 16120 21505 16129 21539
rect 16129 21505 16163 21539
rect 16163 21505 16172 21539
rect 17316 21564 17368 21616
rect 16120 21496 16172 21505
rect 16028 21428 16080 21480
rect 16396 21428 16448 21480
rect 12716 21292 12768 21344
rect 14556 21360 14608 21412
rect 17040 21539 17092 21548
rect 17040 21505 17049 21539
rect 17049 21505 17083 21539
rect 17083 21505 17092 21539
rect 17040 21496 17092 21505
rect 17224 21496 17276 21548
rect 18420 21675 18472 21684
rect 18420 21641 18429 21675
rect 18429 21641 18463 21675
rect 18463 21641 18472 21675
rect 18420 21632 18472 21641
rect 18604 21632 18656 21684
rect 17500 21564 17552 21616
rect 22560 21632 22612 21684
rect 17592 21428 17644 21480
rect 13912 21292 13964 21344
rect 14648 21292 14700 21344
rect 15108 21292 15160 21344
rect 15660 21335 15712 21344
rect 15660 21301 15669 21335
rect 15669 21301 15703 21335
rect 15703 21301 15712 21335
rect 15660 21292 15712 21301
rect 18052 21471 18104 21480
rect 18052 21437 18061 21471
rect 18061 21437 18095 21471
rect 18095 21437 18104 21471
rect 18052 21428 18104 21437
rect 17868 21292 17920 21344
rect 18696 21539 18748 21548
rect 18696 21505 18705 21539
rect 18705 21505 18739 21539
rect 18739 21505 18748 21539
rect 18696 21496 18748 21505
rect 20168 21539 20220 21548
rect 20168 21505 20177 21539
rect 20177 21505 20211 21539
rect 20211 21505 20220 21539
rect 22192 21564 22244 21616
rect 22744 21632 22796 21684
rect 20168 21496 20220 21505
rect 22100 21539 22152 21548
rect 22100 21505 22109 21539
rect 22109 21505 22143 21539
rect 22143 21505 22152 21539
rect 22100 21496 22152 21505
rect 20812 21428 20864 21480
rect 23020 21564 23072 21616
rect 22652 21496 22704 21548
rect 22744 21539 22796 21548
rect 22744 21505 22753 21539
rect 22753 21505 22787 21539
rect 22787 21505 22796 21539
rect 22744 21496 22796 21505
rect 23388 21539 23440 21548
rect 23388 21505 23397 21539
rect 23397 21505 23431 21539
rect 23431 21505 23440 21539
rect 23388 21496 23440 21505
rect 22376 21471 22428 21480
rect 22376 21437 22385 21471
rect 22385 21437 22419 21471
rect 22419 21437 22428 21471
rect 22376 21428 22428 21437
rect 22468 21471 22520 21480
rect 22468 21437 22477 21471
rect 22477 21437 22511 21471
rect 22511 21437 22520 21471
rect 22468 21428 22520 21437
rect 23204 21428 23256 21480
rect 18512 21360 18564 21412
rect 20904 21360 20956 21412
rect 18604 21335 18656 21344
rect 18604 21301 18613 21335
rect 18613 21301 18647 21335
rect 18647 21301 18656 21335
rect 18604 21292 18656 21301
rect 20812 21292 20864 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 2872 21131 2924 21140
rect 2872 21097 2881 21131
rect 2881 21097 2915 21131
rect 2915 21097 2924 21131
rect 2872 21088 2924 21097
rect 5724 21088 5776 21140
rect 6828 21088 6880 21140
rect 8668 21088 8720 21140
rect 5448 20995 5500 21004
rect 5448 20961 5457 20995
rect 5457 20961 5491 20995
rect 5491 20961 5500 20995
rect 5448 20952 5500 20961
rect 1584 20816 1636 20868
rect 5264 20927 5316 20936
rect 5264 20893 5273 20927
rect 5273 20893 5307 20927
rect 5307 20893 5316 20927
rect 5264 20884 5316 20893
rect 5356 20927 5408 20936
rect 5356 20893 5365 20927
rect 5365 20893 5399 20927
rect 5399 20893 5408 20927
rect 5356 20884 5408 20893
rect 4620 20816 4672 20868
rect 6736 21063 6788 21072
rect 6736 21029 6745 21063
rect 6745 21029 6779 21063
rect 6779 21029 6788 21063
rect 6736 21020 6788 21029
rect 10600 21088 10652 21140
rect 10968 21088 11020 21140
rect 15476 21088 15528 21140
rect 15568 21088 15620 21140
rect 15936 21131 15988 21140
rect 15936 21097 15945 21131
rect 15945 21097 15979 21131
rect 15979 21097 15988 21131
rect 15936 21088 15988 21097
rect 16028 21088 16080 21140
rect 17500 21088 17552 21140
rect 17592 21131 17644 21140
rect 17592 21097 17601 21131
rect 17601 21097 17635 21131
rect 17635 21097 17644 21131
rect 17592 21088 17644 21097
rect 18604 21088 18656 21140
rect 18696 21088 18748 21140
rect 19800 21088 19852 21140
rect 20628 21088 20680 21140
rect 21364 21088 21416 21140
rect 22100 21088 22152 21140
rect 22652 21131 22704 21140
rect 22652 21097 22661 21131
rect 22661 21097 22695 21131
rect 22695 21097 22704 21131
rect 22652 21088 22704 21097
rect 22836 21088 22888 21140
rect 23296 21088 23348 21140
rect 12808 21020 12860 21072
rect 14096 21020 14148 21072
rect 16120 21020 16172 21072
rect 7196 20952 7248 21004
rect 8024 20952 8076 21004
rect 9404 20995 9456 21004
rect 9404 20961 9413 20995
rect 9413 20961 9447 20995
rect 9447 20961 9456 20995
rect 9404 20952 9456 20961
rect 13820 20952 13872 21004
rect 14924 20952 14976 21004
rect 15292 20952 15344 21004
rect 7564 20927 7616 20936
rect 7564 20893 7573 20927
rect 7573 20893 7607 20927
rect 7607 20893 7616 20927
rect 7564 20884 7616 20893
rect 7840 20927 7892 20936
rect 7840 20893 7849 20927
rect 7849 20893 7883 20927
rect 7883 20893 7892 20927
rect 7840 20884 7892 20893
rect 7104 20816 7156 20868
rect 9312 20884 9364 20936
rect 2780 20748 2832 20800
rect 5264 20748 5316 20800
rect 6276 20748 6328 20800
rect 7564 20748 7616 20800
rect 9036 20791 9088 20800
rect 9036 20757 9045 20791
rect 9045 20757 9079 20791
rect 9079 20757 9088 20791
rect 9036 20748 9088 20757
rect 9680 20859 9732 20868
rect 9680 20825 9714 20859
rect 9714 20825 9732 20859
rect 9680 20816 9732 20825
rect 14004 20816 14056 20868
rect 15752 20884 15804 20936
rect 15844 20884 15896 20936
rect 17500 20952 17552 21004
rect 15108 20816 15160 20868
rect 10140 20748 10192 20800
rect 10784 20748 10836 20800
rect 12348 20748 12400 20800
rect 14740 20748 14792 20800
rect 15568 20748 15620 20800
rect 16028 20816 16080 20868
rect 16304 20748 16356 20800
rect 16948 20791 17000 20800
rect 16948 20757 16957 20791
rect 16957 20757 16991 20791
rect 16991 20757 17000 20791
rect 16948 20748 17000 20757
rect 18052 20884 18104 20936
rect 18512 20884 18564 20936
rect 18604 20884 18656 20936
rect 18972 20927 19024 20936
rect 18972 20893 18981 20927
rect 18981 20893 19015 20927
rect 19015 20893 19024 20927
rect 18972 20884 19024 20893
rect 22468 21020 22520 21072
rect 19892 20884 19944 20936
rect 20260 20927 20312 20936
rect 20260 20893 20269 20927
rect 20269 20893 20303 20927
rect 20303 20893 20312 20927
rect 20260 20884 20312 20893
rect 20536 20927 20588 20936
rect 20536 20893 20545 20927
rect 20545 20893 20579 20927
rect 20579 20893 20588 20927
rect 20536 20884 20588 20893
rect 20628 20927 20680 20936
rect 20628 20893 20637 20927
rect 20637 20893 20671 20927
rect 20671 20893 20680 20927
rect 20628 20884 20680 20893
rect 20444 20816 20496 20868
rect 20812 20884 20864 20936
rect 20904 20927 20956 20936
rect 20904 20893 20913 20927
rect 20913 20893 20947 20927
rect 20947 20893 20956 20927
rect 20904 20884 20956 20893
rect 21088 20884 21140 20936
rect 22836 20927 22888 20936
rect 22836 20893 22845 20927
rect 22845 20893 22879 20927
rect 22879 20893 22888 20927
rect 22836 20884 22888 20893
rect 20996 20748 21048 20800
rect 22008 20816 22060 20868
rect 22376 20791 22428 20800
rect 22376 20757 22385 20791
rect 22385 20757 22419 20791
rect 22419 20757 22428 20791
rect 22376 20748 22428 20757
rect 23388 20884 23440 20936
rect 25320 20884 25372 20936
rect 23296 20859 23348 20868
rect 23296 20825 23305 20859
rect 23305 20825 23339 20859
rect 23339 20825 23348 20859
rect 23296 20816 23348 20825
rect 22744 20748 22796 20800
rect 4874 20646 4926 20698
rect 4938 20646 4990 20698
rect 5002 20646 5054 20698
rect 5066 20646 5118 20698
rect 5130 20646 5182 20698
rect 5356 20544 5408 20596
rect 6000 20544 6052 20596
rect 7012 20544 7064 20596
rect 9680 20544 9732 20596
rect 12808 20544 12860 20596
rect 13360 20544 13412 20596
rect 20260 20544 20312 20596
rect 5724 20476 5776 20528
rect 6828 20476 6880 20528
rect 8024 20476 8076 20528
rect 10784 20519 10836 20528
rect 10784 20485 10793 20519
rect 10793 20485 10827 20519
rect 10827 20485 10836 20519
rect 10784 20476 10836 20485
rect 3884 20408 3936 20460
rect 5264 20408 5316 20460
rect 6552 20408 6604 20460
rect 10600 20451 10652 20460
rect 10600 20417 10609 20451
rect 10609 20417 10643 20451
rect 10643 20417 10652 20451
rect 10600 20408 10652 20417
rect 3240 20383 3292 20392
rect 3240 20349 3249 20383
rect 3249 20349 3283 20383
rect 3283 20349 3292 20383
rect 3240 20340 3292 20349
rect 6368 20340 6420 20392
rect 9036 20383 9088 20392
rect 9036 20349 9045 20383
rect 9045 20349 9079 20383
rect 9079 20349 9088 20383
rect 9036 20340 9088 20349
rect 10324 20340 10376 20392
rect 11428 20408 11480 20460
rect 12624 20408 12676 20460
rect 13728 20451 13780 20460
rect 7196 20272 7248 20324
rect 8116 20272 8168 20324
rect 2688 20247 2740 20256
rect 2688 20213 2697 20247
rect 2697 20213 2731 20247
rect 2731 20213 2740 20247
rect 2688 20204 2740 20213
rect 4068 20204 4120 20256
rect 5632 20204 5684 20256
rect 6828 20204 6880 20256
rect 10784 20204 10836 20256
rect 13728 20417 13737 20451
rect 13737 20417 13771 20451
rect 13771 20417 13780 20451
rect 13728 20408 13780 20417
rect 16948 20476 17000 20528
rect 18788 20476 18840 20528
rect 20444 20476 20496 20528
rect 14188 20408 14240 20460
rect 14556 20451 14608 20460
rect 14556 20417 14565 20451
rect 14565 20417 14599 20451
rect 14599 20417 14608 20451
rect 14556 20408 14608 20417
rect 15384 20408 15436 20460
rect 17684 20408 17736 20460
rect 19892 20408 19944 20460
rect 15844 20340 15896 20392
rect 24216 20340 24268 20392
rect 15292 20272 15344 20324
rect 20536 20315 20588 20324
rect 20536 20281 20545 20315
rect 20545 20281 20579 20315
rect 20579 20281 20588 20315
rect 20536 20272 20588 20281
rect 24400 20272 24452 20324
rect 13452 20247 13504 20256
rect 13452 20213 13461 20247
rect 13461 20213 13495 20247
rect 13495 20213 13504 20247
rect 13452 20204 13504 20213
rect 14188 20204 14240 20256
rect 15752 20247 15804 20256
rect 15752 20213 15761 20247
rect 15761 20213 15795 20247
rect 15795 20213 15804 20247
rect 15752 20204 15804 20213
rect 21640 20204 21692 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 1308 20000 1360 20052
rect 6368 19975 6420 19984
rect 6368 19941 6377 19975
rect 6377 19941 6411 19975
rect 6411 19941 6420 19975
rect 6368 19932 6420 19941
rect 6552 19975 6604 19984
rect 6552 19941 6561 19975
rect 6561 19941 6595 19975
rect 6595 19941 6604 19975
rect 6552 19932 6604 19941
rect 8024 19975 8076 19984
rect 8024 19941 8033 19975
rect 8033 19941 8067 19975
rect 8067 19941 8076 19975
rect 8024 19932 8076 19941
rect 9312 19932 9364 19984
rect 6184 19864 6236 19916
rect 8116 19907 8168 19916
rect 8116 19873 8125 19907
rect 8125 19873 8159 19907
rect 8159 19873 8168 19907
rect 8116 19864 8168 19873
rect 848 19796 900 19848
rect 2780 19796 2832 19848
rect 2688 19728 2740 19780
rect 3884 19728 3936 19780
rect 8208 19796 8260 19848
rect 9772 19796 9824 19848
rect 10324 19796 10376 19848
rect 11888 20043 11940 20052
rect 11888 20009 11897 20043
rect 11897 20009 11931 20043
rect 11931 20009 11940 20043
rect 11888 20000 11940 20009
rect 15016 20000 15068 20052
rect 14648 19932 14700 19984
rect 15292 20000 15344 20052
rect 15752 20000 15804 20052
rect 16120 20000 16172 20052
rect 12624 19796 12676 19848
rect 13084 19796 13136 19848
rect 15476 19864 15528 19916
rect 15660 19864 15712 19916
rect 17684 20043 17736 20052
rect 17684 20009 17693 20043
rect 17693 20009 17727 20043
rect 17727 20009 17736 20043
rect 17684 20000 17736 20009
rect 18788 20043 18840 20052
rect 18788 20009 18797 20043
rect 18797 20009 18831 20043
rect 18831 20009 18840 20043
rect 18788 20000 18840 20009
rect 20444 20000 20496 20052
rect 20628 20000 20680 20052
rect 14096 19839 14148 19848
rect 14096 19805 14105 19839
rect 14105 19805 14139 19839
rect 14139 19805 14148 19839
rect 14096 19796 14148 19805
rect 6000 19771 6052 19780
rect 6000 19737 6009 19771
rect 6009 19737 6043 19771
rect 6043 19737 6052 19771
rect 6000 19728 6052 19737
rect 6092 19771 6144 19780
rect 6092 19737 6101 19771
rect 6101 19737 6135 19771
rect 6135 19737 6144 19771
rect 6092 19728 6144 19737
rect 7012 19728 7064 19780
rect 7564 19728 7616 19780
rect 1676 19660 1728 19712
rect 5908 19660 5960 19712
rect 6460 19660 6512 19712
rect 13820 19728 13872 19780
rect 14556 19771 14608 19780
rect 9680 19660 9732 19712
rect 10140 19660 10192 19712
rect 14556 19737 14565 19771
rect 14565 19737 14599 19771
rect 14599 19737 14608 19771
rect 14556 19728 14608 19737
rect 15384 19771 15436 19780
rect 15384 19737 15393 19771
rect 15393 19737 15427 19771
rect 15427 19737 15436 19771
rect 15384 19728 15436 19737
rect 15568 19728 15620 19780
rect 15936 19839 15988 19848
rect 15936 19805 15945 19839
rect 15945 19805 15979 19839
rect 15979 19805 15988 19839
rect 15936 19796 15988 19805
rect 16304 19839 16356 19848
rect 16304 19805 16313 19839
rect 16313 19805 16347 19839
rect 16347 19805 16356 19839
rect 16304 19796 16356 19805
rect 18696 19864 18748 19916
rect 22468 20000 22520 20052
rect 24032 20043 24084 20052
rect 24032 20009 24041 20043
rect 24041 20009 24075 20043
rect 24075 20009 24084 20043
rect 24032 20000 24084 20009
rect 24216 20043 24268 20052
rect 24216 20009 24225 20043
rect 24225 20009 24259 20043
rect 24259 20009 24268 20043
rect 24216 20000 24268 20009
rect 17040 19796 17092 19848
rect 18604 19796 18656 19848
rect 14280 19703 14332 19712
rect 14280 19669 14289 19703
rect 14289 19669 14323 19703
rect 14323 19669 14332 19703
rect 14280 19660 14332 19669
rect 14648 19703 14700 19712
rect 14648 19669 14657 19703
rect 14657 19669 14691 19703
rect 14691 19669 14700 19703
rect 14648 19660 14700 19669
rect 14924 19660 14976 19712
rect 15476 19703 15528 19712
rect 15476 19669 15485 19703
rect 15485 19669 15519 19703
rect 15519 19669 15528 19703
rect 16396 19728 16448 19780
rect 16672 19728 16724 19780
rect 18328 19728 18380 19780
rect 18972 19728 19024 19780
rect 19616 19839 19668 19848
rect 19616 19805 19625 19839
rect 19625 19805 19659 19839
rect 19659 19805 19668 19839
rect 19616 19796 19668 19805
rect 19892 19839 19944 19848
rect 19892 19805 19901 19839
rect 19901 19805 19935 19839
rect 19935 19805 19944 19839
rect 19892 19796 19944 19805
rect 20076 19839 20128 19848
rect 20076 19805 20085 19839
rect 20085 19805 20119 19839
rect 20119 19805 20128 19839
rect 20076 19796 20128 19805
rect 19984 19728 20036 19780
rect 22468 19864 22520 19916
rect 21732 19796 21784 19848
rect 21916 19839 21968 19848
rect 21916 19805 21925 19839
rect 21925 19805 21959 19839
rect 21959 19805 21968 19839
rect 21916 19796 21968 19805
rect 20904 19728 20956 19780
rect 15476 19660 15528 19669
rect 16856 19660 16908 19712
rect 17776 19703 17828 19712
rect 17776 19669 17785 19703
rect 17785 19669 17819 19703
rect 17819 19669 17828 19703
rect 17776 19660 17828 19669
rect 21088 19660 21140 19712
rect 21548 19660 21600 19712
rect 23204 19839 23256 19848
rect 23204 19805 23213 19839
rect 23213 19805 23247 19839
rect 23247 19805 23256 19839
rect 23204 19796 23256 19805
rect 22376 19728 22428 19780
rect 23480 19839 23532 19848
rect 23480 19805 23489 19839
rect 23489 19805 23523 19839
rect 23523 19805 23532 19839
rect 23480 19796 23532 19805
rect 24400 19839 24452 19848
rect 24400 19805 24409 19839
rect 24409 19805 24443 19839
rect 24443 19805 24452 19839
rect 24400 19796 24452 19805
rect 25228 19796 25280 19848
rect 23848 19771 23900 19780
rect 23848 19737 23857 19771
rect 23857 19737 23891 19771
rect 23891 19737 23900 19771
rect 23848 19728 23900 19737
rect 23664 19703 23716 19712
rect 23664 19669 23673 19703
rect 23673 19669 23707 19703
rect 23707 19669 23716 19703
rect 23664 19660 23716 19669
rect 23756 19660 23808 19712
rect 4874 19558 4926 19610
rect 4938 19558 4990 19610
rect 5002 19558 5054 19610
rect 5066 19558 5118 19610
rect 5130 19558 5182 19610
rect 6092 19456 6144 19508
rect 6184 19456 6236 19508
rect 6736 19456 6788 19508
rect 7012 19499 7064 19508
rect 7012 19465 7021 19499
rect 7021 19465 7055 19499
rect 7055 19465 7064 19499
rect 7012 19456 7064 19465
rect 7656 19456 7708 19508
rect 2780 19388 2832 19440
rect 1676 19363 1728 19372
rect 1676 19329 1710 19363
rect 1710 19329 1728 19363
rect 1676 19320 1728 19329
rect 3240 19320 3292 19372
rect 6920 19388 6972 19440
rect 9312 19456 9364 19508
rect 10784 19499 10836 19508
rect 10784 19465 10793 19499
rect 10793 19465 10827 19499
rect 10827 19465 10836 19499
rect 10784 19456 10836 19465
rect 11428 19456 11480 19508
rect 13820 19499 13872 19508
rect 13820 19465 13829 19499
rect 13829 19465 13863 19499
rect 13863 19465 13872 19499
rect 13820 19456 13872 19465
rect 3884 19320 3936 19372
rect 4068 19363 4120 19372
rect 4068 19329 4102 19363
rect 4102 19329 4120 19363
rect 4068 19320 4120 19329
rect 5632 19363 5684 19372
rect 5632 19329 5641 19363
rect 5641 19329 5675 19363
rect 5675 19329 5684 19363
rect 5632 19320 5684 19329
rect 5908 19363 5960 19372
rect 5908 19329 5917 19363
rect 5917 19329 5951 19363
rect 5951 19329 5960 19363
rect 5908 19320 5960 19329
rect 6184 19320 6236 19372
rect 6276 19320 6328 19372
rect 6460 19363 6512 19372
rect 6460 19329 6470 19363
rect 6470 19329 6504 19363
rect 6504 19329 6512 19363
rect 6460 19320 6512 19329
rect 6736 19363 6788 19372
rect 6736 19329 6745 19363
rect 6745 19329 6779 19363
rect 6779 19329 6788 19363
rect 6736 19320 6788 19329
rect 6828 19363 6880 19372
rect 6828 19329 6842 19363
rect 6842 19329 6876 19363
rect 6876 19329 6880 19363
rect 6828 19320 6880 19329
rect 10232 19431 10284 19440
rect 10232 19397 10241 19431
rect 10241 19397 10275 19431
rect 10275 19397 10284 19431
rect 10232 19388 10284 19397
rect 10324 19388 10376 19440
rect 14004 19456 14056 19508
rect 7564 19320 7616 19372
rect 7748 19363 7800 19372
rect 7748 19329 7757 19363
rect 7757 19329 7791 19363
rect 7791 19329 7800 19363
rect 7748 19320 7800 19329
rect 9772 19320 9824 19372
rect 11796 19363 11848 19372
rect 11796 19329 11805 19363
rect 11805 19329 11839 19363
rect 11839 19329 11848 19363
rect 11796 19320 11848 19329
rect 14280 19431 14332 19440
rect 14280 19397 14315 19431
rect 14315 19397 14332 19431
rect 14280 19388 14332 19397
rect 12808 19320 12860 19372
rect 12900 19363 12952 19372
rect 12900 19329 12909 19363
rect 12909 19329 12943 19363
rect 12943 19329 12952 19363
rect 12900 19320 12952 19329
rect 13084 19363 13136 19372
rect 13084 19329 13093 19363
rect 13093 19329 13127 19363
rect 13127 19329 13136 19363
rect 13084 19320 13136 19329
rect 13176 19363 13228 19372
rect 13176 19329 13185 19363
rect 13185 19329 13219 19363
rect 13219 19329 13228 19363
rect 13176 19320 13228 19329
rect 13360 19320 13412 19372
rect 13912 19320 13964 19372
rect 7104 19252 7156 19304
rect 7012 19184 7064 19236
rect 10048 19252 10100 19304
rect 11704 19295 11756 19304
rect 11704 19261 11722 19295
rect 11722 19261 11756 19295
rect 11704 19252 11756 19261
rect 10416 19184 10468 19236
rect 11244 19184 11296 19236
rect 12440 19252 12492 19304
rect 13452 19252 13504 19304
rect 14188 19363 14240 19372
rect 14188 19329 14197 19363
rect 14197 19329 14231 19363
rect 14231 19329 14240 19363
rect 14188 19320 14240 19329
rect 14924 19320 14976 19372
rect 15936 19456 15988 19508
rect 16672 19499 16724 19508
rect 16672 19465 16681 19499
rect 16681 19465 16715 19499
rect 16715 19465 16724 19499
rect 16672 19456 16724 19465
rect 19524 19456 19576 19508
rect 19616 19456 19668 19508
rect 12348 19184 12400 19236
rect 14648 19252 14700 19304
rect 14740 19252 14792 19304
rect 15384 19363 15436 19372
rect 15384 19329 15393 19363
rect 15393 19329 15427 19363
rect 15427 19329 15436 19363
rect 15384 19320 15436 19329
rect 15292 19252 15344 19304
rect 15660 19363 15712 19372
rect 15660 19329 15669 19363
rect 15669 19329 15703 19363
rect 15703 19329 15712 19363
rect 15660 19320 15712 19329
rect 15752 19320 15804 19372
rect 16764 19320 16816 19372
rect 16856 19363 16908 19372
rect 16856 19329 16865 19363
rect 16865 19329 16899 19363
rect 16899 19329 16908 19363
rect 16856 19320 16908 19329
rect 17040 19363 17092 19372
rect 17040 19329 17049 19363
rect 17049 19329 17083 19363
rect 17083 19329 17092 19363
rect 17040 19320 17092 19329
rect 17776 19320 17828 19372
rect 18052 19320 18104 19372
rect 8944 19116 8996 19168
rect 9496 19116 9548 19168
rect 11152 19116 11204 19168
rect 13544 19159 13596 19168
rect 13544 19125 13553 19159
rect 13553 19125 13587 19159
rect 13587 19125 13596 19159
rect 13544 19116 13596 19125
rect 14832 19116 14884 19168
rect 18696 19363 18748 19372
rect 18696 19329 18705 19363
rect 18705 19329 18739 19363
rect 18739 19329 18748 19363
rect 18696 19320 18748 19329
rect 18972 19363 19024 19372
rect 18972 19329 18981 19363
rect 18981 19329 19015 19363
rect 19015 19329 19024 19363
rect 18972 19320 19024 19329
rect 19984 19320 20036 19372
rect 20076 19363 20128 19372
rect 20076 19329 20085 19363
rect 20085 19329 20119 19363
rect 20119 19329 20128 19363
rect 20076 19320 20128 19329
rect 20628 19363 20680 19372
rect 20628 19329 20637 19363
rect 20637 19329 20671 19363
rect 20671 19329 20680 19363
rect 20628 19320 20680 19329
rect 21088 19456 21140 19508
rect 23848 19499 23900 19508
rect 23848 19465 23857 19499
rect 23857 19465 23891 19499
rect 23891 19465 23900 19499
rect 23848 19456 23900 19465
rect 20904 19363 20956 19372
rect 20904 19329 20913 19363
rect 20913 19329 20947 19363
rect 20947 19329 20956 19363
rect 20904 19320 20956 19329
rect 23388 19388 23440 19440
rect 23572 19388 23624 19440
rect 23664 19320 23716 19372
rect 23756 19363 23808 19372
rect 23756 19329 23765 19363
rect 23765 19329 23799 19363
rect 23799 19329 23808 19363
rect 23756 19320 23808 19329
rect 24032 19363 24084 19372
rect 24032 19329 24041 19363
rect 24041 19329 24075 19363
rect 24075 19329 24084 19363
rect 24032 19320 24084 19329
rect 25228 19320 25280 19372
rect 21640 19252 21692 19304
rect 24400 19252 24452 19304
rect 24952 19295 25004 19304
rect 24952 19261 24961 19295
rect 24961 19261 24995 19295
rect 24995 19261 25004 19295
rect 24952 19252 25004 19261
rect 18696 19184 18748 19236
rect 21456 19184 21508 19236
rect 18880 19159 18932 19168
rect 18880 19125 18889 19159
rect 18889 19125 18923 19159
rect 18923 19125 18932 19159
rect 18880 19116 18932 19125
rect 20260 19159 20312 19168
rect 20260 19125 20269 19159
rect 20269 19125 20303 19159
rect 20303 19125 20312 19159
rect 20260 19116 20312 19125
rect 21916 19116 21968 19168
rect 23112 19159 23164 19168
rect 23112 19125 23121 19159
rect 23121 19125 23155 19159
rect 23155 19125 23164 19159
rect 23112 19116 23164 19125
rect 23572 19116 23624 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 5264 18912 5316 18964
rect 8668 18912 8720 18964
rect 9864 18912 9916 18964
rect 10416 18955 10468 18964
rect 10416 18921 10425 18955
rect 10425 18921 10459 18955
rect 10459 18921 10468 18955
rect 10416 18912 10468 18921
rect 11244 18955 11296 18964
rect 10140 18844 10192 18896
rect 11244 18921 11253 18955
rect 11253 18921 11287 18955
rect 11287 18921 11296 18955
rect 11244 18912 11296 18921
rect 12348 18955 12400 18964
rect 12348 18921 12357 18955
rect 12357 18921 12391 18955
rect 12391 18921 12400 18955
rect 12348 18912 12400 18921
rect 13176 18955 13228 18964
rect 13176 18921 13185 18955
rect 13185 18921 13219 18955
rect 13219 18921 13228 18955
rect 13176 18912 13228 18921
rect 10692 18844 10744 18896
rect 3884 18819 3936 18828
rect 3884 18785 3893 18819
rect 3893 18785 3927 18819
rect 3927 18785 3936 18819
rect 3884 18776 3936 18785
rect 6000 18708 6052 18760
rect 9680 18708 9732 18760
rect 9956 18751 10008 18760
rect 9956 18717 9965 18751
rect 9965 18717 9999 18751
rect 9999 18717 10008 18751
rect 9956 18708 10008 18717
rect 10048 18751 10100 18760
rect 10048 18717 10057 18751
rect 10057 18717 10091 18751
rect 10091 18717 10100 18751
rect 10048 18708 10100 18717
rect 11152 18776 11204 18828
rect 21640 18955 21692 18964
rect 21640 18921 21649 18955
rect 21649 18921 21683 18955
rect 21683 18921 21692 18955
rect 21640 18912 21692 18921
rect 22836 18912 22888 18964
rect 23112 18912 23164 18964
rect 23756 18912 23808 18964
rect 15292 18844 15344 18896
rect 13360 18776 13412 18828
rect 14648 18776 14700 18828
rect 16120 18776 16172 18828
rect 4804 18640 4856 18692
rect 8300 18640 8352 18692
rect 10324 18640 10376 18692
rect 5724 18572 5776 18624
rect 6644 18572 6696 18624
rect 7012 18572 7064 18624
rect 7104 18572 7156 18624
rect 8944 18572 8996 18624
rect 9036 18615 9088 18624
rect 9036 18581 9045 18615
rect 9045 18581 9079 18615
rect 9079 18581 9088 18615
rect 9036 18572 9088 18581
rect 9680 18572 9732 18624
rect 10968 18572 11020 18624
rect 11612 18751 11664 18760
rect 11612 18717 11621 18751
rect 11621 18717 11655 18751
rect 11655 18717 11664 18751
rect 11612 18708 11664 18717
rect 11704 18708 11756 18760
rect 12164 18751 12216 18760
rect 12164 18717 12173 18751
rect 12173 18717 12207 18751
rect 12207 18717 12216 18751
rect 12164 18708 12216 18717
rect 13268 18751 13320 18760
rect 13268 18717 13277 18751
rect 13277 18717 13311 18751
rect 13311 18717 13320 18751
rect 13268 18708 13320 18717
rect 11980 18640 12032 18692
rect 12440 18640 12492 18692
rect 14740 18708 14792 18760
rect 15200 18708 15252 18760
rect 15476 18708 15528 18760
rect 14556 18640 14608 18692
rect 15384 18640 15436 18692
rect 12624 18572 12676 18624
rect 15752 18572 15804 18624
rect 17040 18572 17092 18624
rect 18328 18751 18380 18760
rect 18328 18717 18337 18751
rect 18337 18717 18371 18751
rect 18371 18717 18380 18751
rect 18328 18708 18380 18717
rect 18420 18751 18472 18760
rect 18420 18717 18429 18751
rect 18429 18717 18463 18751
rect 18463 18717 18472 18751
rect 18420 18708 18472 18717
rect 18696 18751 18748 18760
rect 18696 18717 18705 18751
rect 18705 18717 18739 18751
rect 18739 18717 18748 18751
rect 18696 18708 18748 18717
rect 18880 18751 18932 18760
rect 18880 18717 18889 18751
rect 18889 18717 18923 18751
rect 18923 18717 18932 18751
rect 18880 18708 18932 18717
rect 21456 18751 21508 18760
rect 21456 18717 21465 18751
rect 21465 18717 21499 18751
rect 21499 18717 21508 18751
rect 21456 18708 21508 18717
rect 21732 18751 21784 18760
rect 21732 18717 21741 18751
rect 21741 18717 21775 18751
rect 21775 18717 21784 18751
rect 21732 18708 21784 18717
rect 24676 18708 24728 18760
rect 19892 18640 19944 18692
rect 20628 18640 20680 18692
rect 22652 18683 22704 18692
rect 22652 18649 22661 18683
rect 22661 18649 22695 18683
rect 22695 18649 22704 18683
rect 22652 18640 22704 18649
rect 22836 18683 22888 18692
rect 22836 18649 22845 18683
rect 22845 18649 22879 18683
rect 22879 18649 22888 18683
rect 22836 18640 22888 18649
rect 23388 18640 23440 18692
rect 23848 18640 23900 18692
rect 19064 18572 19116 18624
rect 21456 18572 21508 18624
rect 23572 18572 23624 18624
rect 24032 18572 24084 18624
rect 4874 18470 4926 18522
rect 4938 18470 4990 18522
rect 5002 18470 5054 18522
rect 5066 18470 5118 18522
rect 5130 18470 5182 18522
rect 4804 18411 4856 18420
rect 4804 18377 4813 18411
rect 4813 18377 4847 18411
rect 4847 18377 4856 18411
rect 4804 18368 4856 18377
rect 4896 18368 4948 18420
rect 6000 18368 6052 18420
rect 6184 18368 6236 18420
rect 2320 18232 2372 18284
rect 2872 18232 2924 18284
rect 3056 18232 3108 18284
rect 3976 18232 4028 18284
rect 3884 18096 3936 18148
rect 4896 18232 4948 18284
rect 3608 18071 3660 18080
rect 3608 18037 3617 18071
rect 3617 18037 3651 18071
rect 3651 18037 3660 18071
rect 3608 18028 3660 18037
rect 4160 18028 4212 18080
rect 5172 18275 5224 18284
rect 5172 18241 5181 18275
rect 5181 18241 5215 18275
rect 5215 18241 5224 18275
rect 5172 18232 5224 18241
rect 5264 18275 5316 18284
rect 6644 18300 6696 18352
rect 9772 18368 9824 18420
rect 10324 18411 10376 18420
rect 10324 18377 10333 18411
rect 10333 18377 10367 18411
rect 10367 18377 10376 18411
rect 10324 18368 10376 18377
rect 11520 18368 11572 18420
rect 12348 18368 12400 18420
rect 19524 18411 19576 18420
rect 19524 18377 19533 18411
rect 19533 18377 19567 18411
rect 19567 18377 19576 18411
rect 19524 18368 19576 18377
rect 20260 18411 20312 18420
rect 20260 18377 20269 18411
rect 20269 18377 20303 18411
rect 20303 18377 20312 18411
rect 20260 18368 20312 18377
rect 5264 18241 5299 18275
rect 5299 18241 5316 18275
rect 5264 18232 5316 18241
rect 5724 18164 5776 18216
rect 7472 18275 7524 18284
rect 7472 18241 7506 18275
rect 7506 18241 7524 18275
rect 5540 18096 5592 18148
rect 6000 18096 6052 18148
rect 6644 18096 6696 18148
rect 7472 18232 7524 18241
rect 9312 18232 9364 18284
rect 10048 18275 10100 18284
rect 10048 18241 10057 18275
rect 10057 18241 10091 18275
rect 10091 18241 10100 18275
rect 10048 18232 10100 18241
rect 7012 18164 7064 18216
rect 6092 18028 6144 18080
rect 6552 18071 6604 18080
rect 6552 18037 6561 18071
rect 6561 18037 6595 18071
rect 6595 18037 6604 18071
rect 6552 18028 6604 18037
rect 6920 18028 6972 18080
rect 9496 18164 9548 18216
rect 11152 18232 11204 18284
rect 11980 18275 12032 18284
rect 11980 18241 11989 18275
rect 11989 18241 12023 18275
rect 12023 18241 12032 18275
rect 11980 18232 12032 18241
rect 12072 18232 12124 18284
rect 24676 18411 24728 18420
rect 24676 18377 24685 18411
rect 24685 18377 24719 18411
rect 24719 18377 24728 18411
rect 24676 18368 24728 18377
rect 15016 18300 15068 18352
rect 19064 18343 19116 18352
rect 19064 18309 19073 18343
rect 19073 18309 19107 18343
rect 19107 18309 19116 18343
rect 19064 18300 19116 18309
rect 20444 18343 20496 18352
rect 20444 18309 20453 18343
rect 20453 18309 20487 18343
rect 20487 18309 20496 18343
rect 20444 18300 20496 18309
rect 21916 18300 21968 18352
rect 23388 18343 23440 18352
rect 23388 18309 23397 18343
rect 23397 18309 23431 18343
rect 23431 18309 23440 18343
rect 23388 18300 23440 18309
rect 16764 18232 16816 18284
rect 18788 18232 18840 18284
rect 20076 18275 20128 18284
rect 12992 18164 13044 18216
rect 8668 18071 8720 18080
rect 8668 18037 8677 18071
rect 8677 18037 8711 18071
rect 8711 18037 8720 18071
rect 8668 18028 8720 18037
rect 10508 18028 10560 18080
rect 12716 18028 12768 18080
rect 15476 18028 15528 18080
rect 16304 18164 16356 18216
rect 18052 18164 18104 18216
rect 17684 18096 17736 18148
rect 20076 18241 20085 18275
rect 20085 18241 20119 18275
rect 20119 18241 20128 18275
rect 20076 18232 20128 18241
rect 19340 18164 19392 18216
rect 19800 18207 19852 18216
rect 19800 18173 19809 18207
rect 19809 18173 19843 18207
rect 19843 18173 19852 18207
rect 19800 18164 19852 18173
rect 19892 18164 19944 18216
rect 21824 18232 21876 18284
rect 22376 18275 22428 18284
rect 22376 18241 22385 18275
rect 22385 18241 22419 18275
rect 22419 18241 22428 18275
rect 22376 18232 22428 18241
rect 22836 18232 22888 18284
rect 23572 18275 23624 18284
rect 23572 18241 23581 18275
rect 23581 18241 23615 18275
rect 23615 18241 23624 18275
rect 23572 18232 23624 18241
rect 23756 18275 23808 18284
rect 23756 18241 23764 18275
rect 23764 18241 23798 18275
rect 23798 18241 23808 18275
rect 23756 18232 23808 18241
rect 23848 18275 23900 18284
rect 23848 18241 23857 18275
rect 23857 18241 23891 18275
rect 23891 18241 23900 18275
rect 23848 18232 23900 18241
rect 24400 18275 24452 18284
rect 24400 18241 24409 18275
rect 24409 18241 24443 18275
rect 24443 18241 24452 18275
rect 24400 18232 24452 18241
rect 20812 18207 20864 18216
rect 20812 18173 20821 18207
rect 20821 18173 20855 18207
rect 20855 18173 20864 18207
rect 20812 18164 20864 18173
rect 23664 18207 23716 18216
rect 23664 18173 23673 18207
rect 23673 18173 23707 18207
rect 23707 18173 23716 18207
rect 23664 18164 23716 18173
rect 24952 18232 25004 18284
rect 25596 18275 25648 18284
rect 25596 18241 25605 18275
rect 25605 18241 25639 18275
rect 25639 18241 25648 18275
rect 25596 18232 25648 18241
rect 25044 18207 25096 18216
rect 25044 18173 25053 18207
rect 25053 18173 25087 18207
rect 25087 18173 25096 18207
rect 25044 18164 25096 18173
rect 17960 18028 18012 18080
rect 19432 18071 19484 18080
rect 19432 18037 19441 18071
rect 19441 18037 19475 18071
rect 19475 18037 19484 18071
rect 19432 18028 19484 18037
rect 24584 18028 24636 18080
rect 25596 18028 25648 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 2872 17824 2924 17876
rect 4068 17688 4120 17740
rect 3056 17663 3108 17672
rect 3056 17629 3065 17663
rect 3065 17629 3099 17663
rect 3099 17629 3108 17663
rect 3056 17620 3108 17629
rect 3608 17620 3660 17672
rect 4160 17620 4212 17672
rect 2320 17552 2372 17604
rect 5264 17824 5316 17876
rect 5540 17867 5592 17876
rect 5540 17833 5549 17867
rect 5549 17833 5583 17867
rect 5583 17833 5592 17867
rect 5540 17824 5592 17833
rect 6092 17867 6144 17876
rect 6092 17833 6101 17867
rect 6101 17833 6135 17867
rect 6135 17833 6144 17867
rect 6092 17824 6144 17833
rect 6736 17824 6788 17876
rect 7104 17824 7156 17876
rect 7472 17824 7524 17876
rect 9956 17824 10008 17876
rect 10692 17824 10744 17876
rect 5172 17688 5224 17740
rect 4804 17620 4856 17672
rect 6184 17663 6236 17672
rect 6184 17629 6193 17663
rect 6193 17629 6227 17663
rect 6227 17629 6236 17663
rect 6184 17620 6236 17629
rect 5264 17552 5316 17604
rect 5724 17595 5776 17604
rect 5724 17561 5733 17595
rect 5733 17561 5767 17595
rect 5767 17561 5776 17595
rect 5724 17552 5776 17561
rect 6644 17663 6696 17672
rect 6644 17629 6653 17663
rect 6653 17629 6687 17663
rect 6687 17629 6696 17663
rect 6644 17620 6696 17629
rect 6920 17620 6972 17672
rect 8668 17688 8720 17740
rect 10048 17756 10100 17808
rect 10232 17756 10284 17808
rect 11612 17824 11664 17876
rect 12992 17867 13044 17876
rect 12992 17833 13001 17867
rect 13001 17833 13035 17867
rect 13035 17833 13044 17867
rect 12992 17824 13044 17833
rect 13544 17824 13596 17876
rect 12624 17756 12676 17808
rect 15292 17756 15344 17808
rect 16028 17824 16080 17876
rect 16764 17867 16816 17876
rect 16764 17833 16773 17867
rect 16773 17833 16807 17867
rect 16807 17833 16816 17867
rect 16764 17824 16816 17833
rect 18420 17824 18472 17876
rect 20076 17824 20128 17876
rect 22836 17867 22888 17876
rect 22836 17833 22845 17867
rect 22845 17833 22879 17867
rect 22879 17833 22888 17867
rect 22836 17824 22888 17833
rect 23664 17824 23716 17876
rect 24400 17867 24452 17876
rect 24400 17833 24409 17867
rect 24409 17833 24443 17867
rect 24443 17833 24452 17867
rect 24400 17824 24452 17833
rect 24584 17867 24636 17876
rect 24584 17833 24593 17867
rect 24593 17833 24627 17867
rect 24627 17833 24636 17867
rect 24584 17824 24636 17833
rect 25044 17824 25096 17876
rect 7656 17663 7708 17672
rect 7656 17629 7665 17663
rect 7665 17629 7699 17663
rect 7699 17629 7708 17663
rect 7656 17620 7708 17629
rect 8944 17620 8996 17672
rect 9312 17620 9364 17672
rect 9588 17731 9640 17740
rect 9588 17697 9597 17731
rect 9597 17697 9631 17731
rect 9631 17697 9640 17731
rect 9588 17688 9640 17697
rect 9680 17620 9732 17672
rect 11244 17688 11296 17740
rect 4712 17484 4764 17536
rect 7840 17595 7892 17604
rect 7840 17561 7875 17595
rect 7875 17561 7892 17595
rect 7840 17552 7892 17561
rect 9496 17552 9548 17604
rect 10508 17620 10560 17672
rect 12164 17620 12216 17672
rect 12900 17688 12952 17740
rect 14280 17688 14332 17740
rect 15844 17731 15896 17740
rect 15844 17697 15853 17731
rect 15853 17697 15887 17731
rect 15887 17697 15896 17731
rect 15844 17688 15896 17697
rect 12716 17663 12768 17672
rect 12716 17629 12725 17663
rect 12725 17629 12759 17663
rect 12759 17629 12768 17663
rect 12716 17620 12768 17629
rect 13176 17663 13228 17672
rect 13176 17629 13185 17663
rect 13185 17629 13219 17663
rect 13219 17629 13228 17663
rect 13176 17620 13228 17629
rect 9036 17484 9088 17536
rect 9404 17484 9456 17536
rect 11704 17595 11756 17604
rect 11704 17561 11713 17595
rect 11713 17561 11747 17595
rect 11747 17561 11756 17595
rect 11704 17552 11756 17561
rect 13084 17552 13136 17604
rect 10876 17484 10928 17536
rect 13268 17484 13320 17536
rect 13912 17620 13964 17672
rect 14740 17620 14792 17672
rect 15200 17620 15252 17672
rect 16212 17620 16264 17672
rect 18052 17688 18104 17740
rect 19248 17756 19300 17808
rect 16304 17552 16356 17604
rect 17040 17663 17092 17672
rect 17040 17629 17049 17663
rect 17049 17629 17083 17663
rect 17083 17629 17092 17663
rect 17040 17620 17092 17629
rect 17132 17663 17184 17672
rect 17132 17629 17141 17663
rect 17141 17629 17175 17663
rect 17175 17629 17184 17663
rect 17132 17620 17184 17629
rect 17592 17620 17644 17672
rect 17684 17620 17736 17672
rect 17868 17663 17920 17672
rect 17868 17629 17877 17663
rect 17877 17629 17911 17663
rect 17911 17629 17920 17663
rect 17868 17620 17920 17629
rect 18696 17688 18748 17740
rect 19892 17663 19944 17672
rect 17408 17552 17460 17604
rect 19892 17629 19901 17663
rect 19901 17629 19935 17663
rect 19935 17629 19944 17663
rect 19892 17620 19944 17629
rect 20444 17620 20496 17672
rect 22652 17663 22704 17672
rect 22652 17629 22661 17663
rect 22661 17629 22695 17663
rect 22695 17629 22704 17663
rect 22652 17620 22704 17629
rect 23020 17620 23072 17672
rect 24584 17620 24636 17672
rect 24860 17620 24912 17672
rect 20260 17552 20312 17604
rect 23204 17552 23256 17604
rect 23296 17552 23348 17604
rect 15568 17484 15620 17536
rect 16120 17484 16172 17536
rect 22192 17484 22244 17536
rect 23664 17484 23716 17536
rect 25780 17484 25832 17536
rect 4874 17382 4926 17434
rect 4938 17382 4990 17434
rect 5002 17382 5054 17434
rect 5066 17382 5118 17434
rect 5130 17382 5182 17434
rect 4160 17280 4212 17332
rect 4804 17280 4856 17332
rect 1952 17144 2004 17196
rect 3240 17076 3292 17128
rect 4068 17187 4120 17196
rect 4068 17153 4077 17187
rect 4077 17153 4111 17187
rect 4111 17153 4120 17187
rect 4068 17144 4120 17153
rect 4712 17187 4764 17196
rect 4712 17153 4721 17187
rect 4721 17153 4755 17187
rect 4755 17153 4764 17187
rect 4712 17144 4764 17153
rect 4804 17144 4856 17196
rect 4620 17076 4672 17128
rect 5264 17187 5316 17196
rect 5264 17153 5273 17187
rect 5273 17153 5307 17187
rect 5307 17153 5316 17187
rect 5264 17144 5316 17153
rect 5448 17144 5500 17196
rect 6184 17144 6236 17196
rect 6552 17144 6604 17196
rect 8116 17280 8168 17332
rect 9036 17280 9088 17332
rect 10140 17280 10192 17332
rect 10692 17280 10744 17332
rect 11796 17280 11848 17332
rect 14740 17323 14792 17332
rect 14740 17289 14749 17323
rect 14749 17289 14783 17323
rect 14783 17289 14792 17323
rect 14740 17280 14792 17289
rect 14924 17280 14976 17332
rect 9312 17212 9364 17264
rect 8116 17187 8168 17196
rect 8116 17153 8125 17187
rect 8125 17153 8159 17187
rect 8159 17153 8168 17187
rect 8116 17144 8168 17153
rect 8484 17187 8536 17196
rect 8484 17153 8493 17187
rect 8493 17153 8527 17187
rect 8527 17153 8536 17187
rect 8484 17144 8536 17153
rect 9404 17144 9456 17196
rect 10048 17187 10100 17196
rect 10048 17153 10057 17187
rect 10057 17153 10091 17187
rect 10091 17153 10100 17187
rect 10048 17144 10100 17153
rect 5724 17008 5776 17060
rect 9588 17076 9640 17128
rect 6552 17008 6604 17060
rect 10232 17119 10284 17128
rect 10232 17085 10241 17119
rect 10241 17085 10275 17119
rect 10275 17085 10284 17119
rect 10232 17076 10284 17085
rect 2412 16940 2464 16992
rect 2872 16983 2924 16992
rect 2872 16949 2881 16983
rect 2881 16949 2915 16983
rect 2915 16949 2924 16983
rect 2872 16940 2924 16949
rect 3608 16983 3660 16992
rect 3608 16949 3617 16983
rect 3617 16949 3651 16983
rect 3651 16949 3660 16983
rect 3608 16940 3660 16949
rect 3976 16940 4028 16992
rect 4068 16940 4120 16992
rect 5448 16983 5500 16992
rect 5448 16949 5457 16983
rect 5457 16949 5491 16983
rect 5491 16949 5500 16983
rect 5448 16940 5500 16949
rect 5816 16940 5868 16992
rect 6368 16983 6420 16992
rect 6368 16949 6377 16983
rect 6377 16949 6411 16983
rect 6411 16949 6420 16983
rect 6368 16940 6420 16949
rect 6460 16940 6512 16992
rect 7656 16983 7708 16992
rect 7656 16949 7665 16983
rect 7665 16949 7699 16983
rect 7699 16949 7708 16983
rect 7656 16940 7708 16949
rect 9956 16983 10008 16992
rect 9956 16949 9965 16983
rect 9965 16949 9999 16983
rect 9999 16949 10008 16983
rect 9956 16940 10008 16949
rect 10232 16983 10284 16992
rect 10232 16949 10241 16983
rect 10241 16949 10275 16983
rect 10275 16949 10284 16983
rect 10232 16940 10284 16949
rect 11336 17212 11388 17264
rect 11152 17144 11204 17196
rect 13820 17144 13872 17196
rect 17408 17280 17460 17332
rect 17592 17280 17644 17332
rect 11612 17008 11664 17060
rect 12072 17051 12124 17060
rect 12072 17017 12081 17051
rect 12081 17017 12115 17051
rect 12115 17017 12124 17051
rect 12072 17008 12124 17017
rect 12440 16940 12492 16992
rect 13912 17119 13964 17128
rect 13912 17085 13921 17119
rect 13921 17085 13955 17119
rect 13955 17085 13964 17119
rect 13912 17076 13964 17085
rect 15108 17187 15160 17196
rect 15108 17153 15117 17187
rect 15117 17153 15151 17187
rect 15151 17153 15160 17187
rect 15108 17144 15160 17153
rect 15660 17144 15712 17196
rect 15752 17187 15804 17196
rect 15752 17153 15761 17187
rect 15761 17153 15795 17187
rect 15795 17153 15804 17187
rect 15752 17144 15804 17153
rect 16672 17255 16724 17264
rect 16672 17221 16681 17255
rect 16681 17221 16715 17255
rect 16715 17221 16724 17255
rect 16672 17212 16724 17221
rect 17132 17212 17184 17264
rect 18052 17280 18104 17332
rect 20812 17280 20864 17332
rect 21824 17323 21876 17332
rect 21824 17289 21833 17323
rect 21833 17289 21867 17323
rect 21867 17289 21876 17323
rect 21824 17280 21876 17289
rect 22192 17280 22244 17332
rect 22284 17280 22336 17332
rect 16028 17187 16080 17196
rect 16028 17153 16037 17187
rect 16037 17153 16071 17187
rect 16071 17153 16080 17187
rect 16028 17144 16080 17153
rect 16304 17187 16356 17196
rect 16304 17153 16313 17187
rect 16313 17153 16347 17187
rect 16347 17153 16356 17187
rect 16304 17144 16356 17153
rect 17500 17187 17552 17196
rect 15384 17119 15436 17128
rect 15384 17085 15393 17119
rect 15393 17085 15427 17119
rect 15427 17085 15436 17119
rect 15384 17076 15436 17085
rect 15568 17076 15620 17128
rect 12808 16940 12860 16992
rect 16304 17008 16356 17060
rect 17500 17153 17509 17187
rect 17509 17153 17543 17187
rect 17543 17153 17552 17187
rect 17500 17144 17552 17153
rect 17868 17144 17920 17196
rect 17960 17187 18012 17196
rect 17960 17153 17969 17187
rect 17969 17153 18003 17187
rect 18003 17153 18012 17187
rect 17960 17144 18012 17153
rect 18052 17144 18104 17196
rect 20444 17187 20496 17196
rect 20444 17153 20453 17187
rect 20453 17153 20487 17187
rect 20487 17153 20496 17187
rect 20444 17144 20496 17153
rect 17960 17008 18012 17060
rect 19432 16940 19484 16992
rect 20720 17187 20772 17196
rect 20720 17153 20729 17187
rect 20729 17153 20763 17187
rect 20763 17153 20772 17187
rect 20720 17144 20772 17153
rect 20904 17187 20956 17196
rect 20904 17153 20913 17187
rect 20913 17153 20947 17187
rect 20947 17153 20956 17187
rect 20904 17144 20956 17153
rect 21180 17187 21232 17196
rect 21180 17153 21189 17187
rect 21189 17153 21223 17187
rect 21223 17153 21232 17187
rect 21180 17144 21232 17153
rect 22836 17280 22888 17332
rect 23204 17323 23256 17332
rect 23204 17289 23213 17323
rect 23213 17289 23247 17323
rect 23247 17289 23256 17323
rect 23204 17280 23256 17289
rect 24952 17280 25004 17332
rect 25320 17280 25372 17332
rect 26424 17280 26476 17332
rect 20996 17076 21048 17128
rect 21640 17187 21692 17196
rect 21640 17153 21649 17187
rect 21649 17153 21683 17187
rect 21683 17153 21692 17187
rect 21640 17144 21692 17153
rect 22376 17187 22428 17196
rect 22376 17153 22385 17187
rect 22385 17153 22419 17187
rect 22419 17153 22428 17187
rect 22376 17144 22428 17153
rect 23664 17144 23716 17196
rect 24584 17144 24636 17196
rect 24860 17144 24912 17196
rect 25504 17187 25556 17196
rect 25504 17153 25513 17187
rect 25513 17153 25547 17187
rect 25547 17153 25556 17187
rect 25504 17144 25556 17153
rect 21180 16940 21232 16992
rect 25780 17187 25832 17196
rect 25780 17153 25789 17187
rect 25789 17153 25823 17187
rect 25823 17153 25832 17187
rect 25780 17144 25832 17153
rect 25872 17144 25924 17196
rect 22836 16940 22888 16992
rect 23388 16983 23440 16992
rect 23388 16949 23397 16983
rect 23397 16949 23431 16983
rect 23431 16949 23440 16983
rect 23388 16940 23440 16949
rect 25596 16940 25648 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 1952 16779 2004 16788
rect 1952 16745 1961 16779
rect 1961 16745 1995 16779
rect 1995 16745 2004 16779
rect 1952 16736 2004 16745
rect 2596 16668 2648 16720
rect 2872 16668 2924 16720
rect 2964 16711 3016 16720
rect 2964 16677 2973 16711
rect 2973 16677 3007 16711
rect 3007 16677 3016 16711
rect 2964 16668 3016 16677
rect 2596 16575 2648 16584
rect 2596 16541 2605 16575
rect 2605 16541 2639 16575
rect 2639 16541 2648 16575
rect 2596 16532 2648 16541
rect 4804 16736 4856 16788
rect 6368 16736 6420 16788
rect 9588 16779 9640 16788
rect 9588 16745 9597 16779
rect 9597 16745 9631 16779
rect 9631 16745 9640 16779
rect 9588 16736 9640 16745
rect 10048 16736 10100 16788
rect 10600 16736 10652 16788
rect 11060 16779 11112 16788
rect 11060 16745 11069 16779
rect 11069 16745 11103 16779
rect 11103 16745 11112 16779
rect 11060 16736 11112 16745
rect 13084 16736 13136 16788
rect 13912 16736 13964 16788
rect 4436 16668 4488 16720
rect 5264 16668 5316 16720
rect 8576 16668 8628 16720
rect 9496 16668 9548 16720
rect 3884 16532 3936 16584
rect 3976 16575 4028 16584
rect 3976 16541 3985 16575
rect 3985 16541 4019 16575
rect 4019 16541 4028 16575
rect 3976 16532 4028 16541
rect 5448 16600 5500 16652
rect 9956 16600 10008 16652
rect 11520 16600 11572 16652
rect 11980 16643 12032 16652
rect 11980 16609 11989 16643
rect 11989 16609 12023 16643
rect 12023 16609 12032 16643
rect 11980 16600 12032 16609
rect 4436 16575 4488 16584
rect 4436 16541 4445 16575
rect 4445 16541 4479 16575
rect 4479 16541 4488 16575
rect 4436 16532 4488 16541
rect 4620 16575 4672 16584
rect 4620 16541 4629 16575
rect 4629 16541 4663 16575
rect 4663 16541 4672 16575
rect 4620 16532 4672 16541
rect 5816 16575 5868 16584
rect 5816 16541 5825 16575
rect 5825 16541 5859 16575
rect 5859 16541 5868 16575
rect 5816 16532 5868 16541
rect 6000 16532 6052 16584
rect 6460 16532 6512 16584
rect 6552 16575 6604 16584
rect 6552 16541 6561 16575
rect 6561 16541 6595 16575
rect 6595 16541 6604 16575
rect 6552 16532 6604 16541
rect 6828 16575 6880 16584
rect 6828 16541 6837 16575
rect 6837 16541 6871 16575
rect 6871 16541 6880 16575
rect 6828 16532 6880 16541
rect 7656 16532 7708 16584
rect 8852 16532 8904 16584
rect 2320 16507 2372 16516
rect 2320 16473 2329 16507
rect 2329 16473 2363 16507
rect 2363 16473 2372 16507
rect 2320 16464 2372 16473
rect 2504 16464 2556 16516
rect 3608 16464 3660 16516
rect 6184 16507 6236 16516
rect 6184 16473 6193 16507
rect 6193 16473 6227 16507
rect 6227 16473 6236 16507
rect 6184 16464 6236 16473
rect 9404 16532 9456 16584
rect 11888 16532 11940 16584
rect 12164 16575 12216 16584
rect 12164 16541 12173 16575
rect 12173 16541 12207 16575
rect 12207 16541 12216 16575
rect 12164 16532 12216 16541
rect 13452 16600 13504 16652
rect 14280 16600 14332 16652
rect 15476 16736 15528 16788
rect 17960 16736 18012 16788
rect 19984 16736 20036 16788
rect 20444 16736 20496 16788
rect 20996 16779 21048 16788
rect 20996 16745 21005 16779
rect 21005 16745 21039 16779
rect 21039 16745 21048 16779
rect 20996 16736 21048 16745
rect 21088 16736 21140 16788
rect 23572 16736 23624 16788
rect 17132 16668 17184 16720
rect 17224 16643 17276 16652
rect 17224 16609 17233 16643
rect 17233 16609 17267 16643
rect 17267 16609 17276 16643
rect 17224 16600 17276 16609
rect 19156 16600 19208 16652
rect 20720 16600 20772 16652
rect 20904 16668 20956 16720
rect 21640 16668 21692 16720
rect 21180 16600 21232 16652
rect 12808 16532 12860 16584
rect 14372 16532 14424 16584
rect 15568 16532 15620 16584
rect 18052 16532 18104 16584
rect 4252 16439 4304 16448
rect 4252 16405 4261 16439
rect 4261 16405 4295 16439
rect 4295 16405 4304 16439
rect 4252 16396 4304 16405
rect 4528 16439 4580 16448
rect 4528 16405 4537 16439
rect 4537 16405 4571 16439
rect 4571 16405 4580 16439
rect 4528 16396 4580 16405
rect 5632 16439 5684 16448
rect 5632 16405 5641 16439
rect 5641 16405 5675 16439
rect 5675 16405 5684 16439
rect 5632 16396 5684 16405
rect 9680 16464 9732 16516
rect 10692 16464 10744 16516
rect 8944 16396 8996 16448
rect 11704 16507 11756 16516
rect 11704 16473 11713 16507
rect 11713 16473 11747 16507
rect 11747 16473 11756 16507
rect 11704 16464 11756 16473
rect 14740 16507 14792 16516
rect 14740 16473 14774 16507
rect 14774 16473 14792 16507
rect 14740 16464 14792 16473
rect 19708 16464 19760 16516
rect 19984 16575 20036 16584
rect 19984 16541 19993 16575
rect 19993 16541 20027 16575
rect 20027 16541 20036 16575
rect 19984 16532 20036 16541
rect 20352 16575 20404 16584
rect 20352 16541 20361 16575
rect 20361 16541 20395 16575
rect 20395 16541 20404 16575
rect 20352 16532 20404 16541
rect 21364 16575 21416 16584
rect 21364 16541 21373 16575
rect 21373 16541 21407 16575
rect 21407 16541 21416 16575
rect 21364 16532 21416 16541
rect 20260 16464 20312 16516
rect 13268 16396 13320 16448
rect 14280 16439 14332 16448
rect 14280 16405 14289 16439
rect 14289 16405 14323 16439
rect 14323 16405 14332 16439
rect 14280 16396 14332 16405
rect 15660 16396 15712 16448
rect 19248 16396 19300 16448
rect 20352 16396 20404 16448
rect 20720 16396 20772 16448
rect 21916 16532 21968 16584
rect 23112 16575 23164 16584
rect 23112 16541 23121 16575
rect 23121 16541 23155 16575
rect 23155 16541 23164 16575
rect 23112 16532 23164 16541
rect 22836 16464 22888 16516
rect 24032 16575 24084 16584
rect 24032 16541 24041 16575
rect 24041 16541 24075 16575
rect 24075 16541 24084 16575
rect 24032 16532 24084 16541
rect 23388 16396 23440 16448
rect 25136 16396 25188 16448
rect 4874 16294 4926 16346
rect 4938 16294 4990 16346
rect 5002 16294 5054 16346
rect 5066 16294 5118 16346
rect 5130 16294 5182 16346
rect 2320 16192 2372 16244
rect 2504 16192 2556 16244
rect 7840 16192 7892 16244
rect 3976 16124 4028 16176
rect 4252 16099 4304 16108
rect 4252 16065 4261 16099
rect 4261 16065 4295 16099
rect 4295 16065 4304 16099
rect 4252 16056 4304 16065
rect 4804 16124 4856 16176
rect 11704 16192 11756 16244
rect 12532 16235 12584 16244
rect 12532 16201 12541 16235
rect 12541 16201 12575 16235
rect 12575 16201 12584 16235
rect 12532 16192 12584 16201
rect 10232 16167 10284 16176
rect 4528 16056 4580 16108
rect 4712 16056 4764 16108
rect 5724 16056 5776 16108
rect 5908 16056 5960 16108
rect 6828 16056 6880 16108
rect 4620 15988 4672 16040
rect 7656 16099 7708 16108
rect 7656 16065 7665 16099
rect 7665 16065 7699 16099
rect 7699 16065 7708 16099
rect 7656 16056 7708 16065
rect 7748 16099 7800 16108
rect 7748 16065 7757 16099
rect 7757 16065 7791 16099
rect 7791 16065 7800 16099
rect 7748 16056 7800 16065
rect 8116 16056 8168 16108
rect 8392 16056 8444 16108
rect 8484 16056 8536 16108
rect 9956 16056 10008 16108
rect 10232 16133 10241 16167
rect 10241 16133 10275 16167
rect 10275 16133 10284 16167
rect 10232 16124 10284 16133
rect 10784 16124 10836 16176
rect 10876 16167 10928 16176
rect 10876 16133 10885 16167
rect 10885 16133 10919 16167
rect 10919 16133 10928 16167
rect 10876 16124 10928 16133
rect 11060 16124 11112 16176
rect 13452 16167 13504 16176
rect 5448 15920 5500 15972
rect 6184 15895 6236 15904
rect 6184 15861 6193 15895
rect 6193 15861 6227 15895
rect 6227 15861 6236 15895
rect 6184 15852 6236 15861
rect 7196 15852 7248 15904
rect 8116 15852 8168 15904
rect 8300 15895 8352 15904
rect 8300 15861 8309 15895
rect 8309 15861 8343 15895
rect 8343 15861 8352 15895
rect 8300 15852 8352 15861
rect 8576 16031 8628 16040
rect 8576 15997 8585 16031
rect 8585 15997 8619 16031
rect 8619 15997 8628 16031
rect 8576 15988 8628 15997
rect 8852 15988 8904 16040
rect 10416 16099 10468 16108
rect 10416 16065 10461 16099
rect 10461 16065 10468 16099
rect 10416 16056 10468 16065
rect 10600 16099 10652 16108
rect 10600 16065 10609 16099
rect 10609 16065 10643 16099
rect 10643 16065 10652 16099
rect 10600 16056 10652 16065
rect 10692 16056 10744 16108
rect 9864 15852 9916 15904
rect 10416 15852 10468 15904
rect 10600 15852 10652 15904
rect 11336 15920 11388 15972
rect 11888 16056 11940 16108
rect 12808 16099 12860 16108
rect 12808 16065 12817 16099
rect 12817 16065 12851 16099
rect 12851 16065 12860 16099
rect 12808 16056 12860 16065
rect 13452 16133 13469 16167
rect 13469 16133 13504 16167
rect 13452 16124 13504 16133
rect 13820 16192 13872 16244
rect 14924 16192 14976 16244
rect 15200 16235 15252 16244
rect 15200 16201 15209 16235
rect 15209 16201 15243 16235
rect 15243 16201 15252 16235
rect 15200 16192 15252 16201
rect 19156 16192 19208 16244
rect 21824 16192 21876 16244
rect 13268 16099 13320 16108
rect 13268 16065 13277 16099
rect 13277 16065 13311 16099
rect 13311 16065 13320 16099
rect 13268 16056 13320 16065
rect 13544 16099 13596 16108
rect 13544 16065 13553 16099
rect 13553 16065 13587 16099
rect 13587 16065 13596 16099
rect 13544 16056 13596 16065
rect 17684 16124 17736 16176
rect 24952 16124 25004 16176
rect 25228 16124 25280 16176
rect 12900 16031 12952 16040
rect 12900 15997 12909 16031
rect 12909 15997 12943 16031
rect 12943 15997 12952 16031
rect 12900 15988 12952 15997
rect 11152 15852 11204 15904
rect 11796 15895 11848 15904
rect 11796 15861 11805 15895
rect 11805 15861 11839 15895
rect 11839 15861 11848 15895
rect 11796 15852 11848 15861
rect 13728 15920 13780 15972
rect 14280 16056 14332 16108
rect 15108 16099 15160 16108
rect 15108 16065 15117 16099
rect 15117 16065 15151 16099
rect 15151 16065 15160 16099
rect 15108 16056 15160 16065
rect 15844 16056 15896 16108
rect 16856 16099 16908 16108
rect 16856 16065 16865 16099
rect 16865 16065 16899 16099
rect 16899 16065 16908 16099
rect 16856 16056 16908 16065
rect 15016 15988 15068 16040
rect 17224 16056 17276 16108
rect 24584 16056 24636 16108
rect 24860 16099 24912 16108
rect 24860 16065 24869 16099
rect 24869 16065 24903 16099
rect 24903 16065 24912 16099
rect 24860 16056 24912 16065
rect 17132 16031 17184 16040
rect 17132 15997 17141 16031
rect 17141 15997 17175 16031
rect 17175 15997 17184 16031
rect 17132 15988 17184 15997
rect 25504 16099 25556 16108
rect 25504 16065 25513 16099
rect 25513 16065 25547 16099
rect 25547 16065 25556 16099
rect 25504 16056 25556 16065
rect 16396 15920 16448 15972
rect 17776 15920 17828 15972
rect 17408 15852 17460 15904
rect 25320 15852 25372 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 7748 15648 7800 15700
rect 11704 15648 11756 15700
rect 4620 15512 4672 15564
rect 2780 15444 2832 15496
rect 2504 15376 2556 15428
rect 2780 15308 2832 15360
rect 3976 15444 4028 15496
rect 4712 15444 4764 15496
rect 7656 15580 7708 15632
rect 11796 15580 11848 15632
rect 6184 15555 6236 15564
rect 6184 15521 6193 15555
rect 6193 15521 6227 15555
rect 6227 15521 6236 15555
rect 6184 15512 6236 15521
rect 8116 15512 8168 15564
rect 5724 15376 5776 15428
rect 6092 15487 6144 15496
rect 6092 15453 6101 15487
rect 6101 15453 6135 15487
rect 6135 15453 6144 15487
rect 6092 15444 6144 15453
rect 6552 15444 6604 15496
rect 8024 15487 8076 15496
rect 8024 15453 8033 15487
rect 8033 15453 8067 15487
rect 8067 15453 8076 15487
rect 8024 15444 8076 15453
rect 11980 15512 12032 15564
rect 13820 15512 13872 15564
rect 7656 15376 7708 15428
rect 8392 15444 8444 15496
rect 8484 15487 8536 15496
rect 8484 15453 8493 15487
rect 8493 15453 8527 15487
rect 8527 15453 8536 15487
rect 8484 15444 8536 15453
rect 12532 15444 12584 15496
rect 15016 15487 15068 15496
rect 15016 15453 15025 15487
rect 15025 15453 15059 15487
rect 15059 15453 15068 15487
rect 15016 15444 15068 15453
rect 17684 15648 17736 15700
rect 15752 15580 15804 15632
rect 15384 15444 15436 15496
rect 15476 15444 15528 15496
rect 17408 15487 17460 15496
rect 17408 15453 17417 15487
rect 17417 15453 17451 15487
rect 17451 15453 17460 15487
rect 17408 15444 17460 15453
rect 19248 15623 19300 15632
rect 19248 15589 19257 15623
rect 19257 15589 19291 15623
rect 19291 15589 19300 15623
rect 19248 15580 19300 15589
rect 17684 15512 17736 15564
rect 17592 15487 17644 15496
rect 17592 15453 17601 15487
rect 17601 15453 17635 15487
rect 17635 15453 17644 15487
rect 17592 15444 17644 15453
rect 20812 15648 20864 15700
rect 21640 15648 21692 15700
rect 22008 15648 22060 15700
rect 25504 15648 25556 15700
rect 20628 15580 20680 15632
rect 19432 15444 19484 15496
rect 8852 15376 8904 15428
rect 11152 15376 11204 15428
rect 15568 15376 15620 15428
rect 20352 15444 20404 15496
rect 20812 15487 20864 15496
rect 20812 15453 20820 15487
rect 20820 15453 20854 15487
rect 20854 15453 20864 15487
rect 20812 15444 20864 15453
rect 24676 15555 24728 15564
rect 24676 15521 24685 15555
rect 24685 15521 24719 15555
rect 24719 15521 24728 15555
rect 24676 15512 24728 15521
rect 25044 15512 25096 15564
rect 21272 15487 21324 15496
rect 21272 15453 21281 15487
rect 21281 15453 21315 15487
rect 21315 15453 21324 15487
rect 21272 15444 21324 15453
rect 21456 15487 21508 15496
rect 21456 15453 21465 15487
rect 21465 15453 21499 15487
rect 21499 15453 21508 15487
rect 21456 15444 21508 15453
rect 21548 15487 21600 15496
rect 21548 15453 21557 15487
rect 21557 15453 21591 15487
rect 21591 15453 21600 15487
rect 21548 15444 21600 15453
rect 21180 15376 21232 15428
rect 4804 15308 4856 15360
rect 5356 15308 5408 15360
rect 5540 15308 5592 15360
rect 8392 15351 8444 15360
rect 8392 15317 8401 15351
rect 8401 15317 8435 15351
rect 8435 15317 8444 15351
rect 8392 15308 8444 15317
rect 13268 15308 13320 15360
rect 13452 15308 13504 15360
rect 14096 15308 14148 15360
rect 15200 15308 15252 15360
rect 15384 15308 15436 15360
rect 15660 15308 15712 15360
rect 16396 15308 16448 15360
rect 17132 15308 17184 15360
rect 17868 15308 17920 15360
rect 20076 15308 20128 15360
rect 20720 15308 20772 15360
rect 22192 15444 22244 15496
rect 23572 15444 23624 15496
rect 24124 15487 24176 15496
rect 24124 15453 24133 15487
rect 24133 15453 24167 15487
rect 24167 15453 24176 15487
rect 24124 15444 24176 15453
rect 24216 15487 24268 15496
rect 24216 15453 24225 15487
rect 24225 15453 24259 15487
rect 24259 15453 24268 15487
rect 24216 15444 24268 15453
rect 25228 15487 25280 15496
rect 25228 15453 25237 15487
rect 25237 15453 25271 15487
rect 25271 15453 25280 15487
rect 25228 15444 25280 15453
rect 24952 15376 25004 15428
rect 25320 15376 25372 15428
rect 26424 15487 26476 15496
rect 26424 15453 26433 15487
rect 26433 15453 26467 15487
rect 26467 15453 26476 15487
rect 26424 15444 26476 15453
rect 24032 15308 24084 15360
rect 24584 15308 24636 15360
rect 25136 15308 25188 15360
rect 4874 15206 4926 15258
rect 4938 15206 4990 15258
rect 5002 15206 5054 15258
rect 5066 15206 5118 15258
rect 5130 15206 5182 15258
rect 2504 15147 2556 15156
rect 2504 15113 2513 15147
rect 2513 15113 2547 15147
rect 2547 15113 2556 15147
rect 2504 15104 2556 15113
rect 3884 15104 3936 15156
rect 2780 15036 2832 15088
rect 1952 15011 2004 15020
rect 1952 14977 1961 15011
rect 1961 14977 1995 15011
rect 1995 14977 2004 15011
rect 1952 14968 2004 14977
rect 2044 14968 2096 15020
rect 2320 15011 2372 15020
rect 2320 14977 2329 15011
rect 2329 14977 2363 15011
rect 2363 14977 2372 15011
rect 2320 14968 2372 14977
rect 3240 15011 3292 15020
rect 3240 14977 3249 15011
rect 3249 14977 3283 15011
rect 3283 14977 3292 15011
rect 3240 14968 3292 14977
rect 3884 15011 3936 15020
rect 3884 14977 3893 15011
rect 3893 14977 3927 15011
rect 3927 14977 3936 15011
rect 3884 14968 3936 14977
rect 8392 15104 8444 15156
rect 4068 14968 4120 15020
rect 4988 15011 5040 15020
rect 4988 14977 4997 15011
rect 4997 14977 5031 15011
rect 5031 14977 5040 15011
rect 4988 14968 5040 14977
rect 6000 15036 6052 15088
rect 7656 15036 7708 15088
rect 9036 15079 9088 15088
rect 9036 15045 9045 15079
rect 9045 15045 9079 15079
rect 9079 15045 9088 15079
rect 9036 15036 9088 15045
rect 5724 15011 5776 15020
rect 5724 14977 5733 15011
rect 5733 14977 5767 15011
rect 5767 14977 5776 15011
rect 5724 14968 5776 14977
rect 6092 14968 6144 15020
rect 7196 15011 7248 15020
rect 7196 14977 7205 15011
rect 7205 14977 7239 15011
rect 7239 14977 7248 15011
rect 7196 14968 7248 14977
rect 7288 15011 7340 15020
rect 7288 14977 7297 15011
rect 7297 14977 7331 15011
rect 7331 14977 7340 15011
rect 9680 15104 9732 15156
rect 10968 15104 11020 15156
rect 10692 15036 10744 15088
rect 11888 15104 11940 15156
rect 12348 15104 12400 15156
rect 14740 15147 14792 15156
rect 14740 15113 14749 15147
rect 14749 15113 14783 15147
rect 14783 15113 14792 15147
rect 14740 15104 14792 15113
rect 7288 14968 7340 14977
rect 9680 15011 9732 15020
rect 9680 14977 9689 15011
rect 9689 14977 9723 15011
rect 9723 14977 9732 15011
rect 9680 14968 9732 14977
rect 10600 15011 10652 15020
rect 10600 14977 10609 15011
rect 10609 14977 10643 15011
rect 10643 14977 10652 15011
rect 10600 14968 10652 14977
rect 4712 14900 4764 14952
rect 8852 14943 8904 14952
rect 8852 14909 8861 14943
rect 8861 14909 8895 14943
rect 8895 14909 8904 14943
rect 8852 14900 8904 14909
rect 4160 14875 4212 14884
rect 4160 14841 4169 14875
rect 4169 14841 4203 14875
rect 4203 14841 4212 14875
rect 4160 14832 4212 14841
rect 3976 14764 4028 14816
rect 4988 14832 5040 14884
rect 8760 14832 8812 14884
rect 8944 14832 8996 14884
rect 4620 14807 4672 14816
rect 4620 14773 4629 14807
rect 4629 14773 4663 14807
rect 4663 14773 4672 14807
rect 4620 14764 4672 14773
rect 5908 14807 5960 14816
rect 5908 14773 5917 14807
rect 5917 14773 5951 14807
rect 5951 14773 5960 14807
rect 5908 14764 5960 14773
rect 6368 14764 6420 14816
rect 6552 14807 6604 14816
rect 6552 14773 6561 14807
rect 6561 14773 6595 14807
rect 6595 14773 6604 14807
rect 6552 14764 6604 14773
rect 8668 14764 8720 14816
rect 9956 14943 10008 14952
rect 9956 14909 9965 14943
rect 9965 14909 9999 14943
rect 9999 14909 10008 14943
rect 9956 14900 10008 14909
rect 10140 14900 10192 14952
rect 10048 14832 10100 14884
rect 10508 14900 10560 14952
rect 10876 14900 10928 14952
rect 11060 15011 11112 15020
rect 11060 14977 11069 15011
rect 11069 14977 11103 15011
rect 11103 14977 11112 15011
rect 11060 14968 11112 14977
rect 11152 15011 11204 15020
rect 11152 14977 11161 15011
rect 11161 14977 11195 15011
rect 11195 14977 11204 15011
rect 11152 14968 11204 14977
rect 13728 15036 13780 15088
rect 13820 15079 13872 15088
rect 13820 15045 13829 15079
rect 13829 15045 13863 15079
rect 13863 15045 13872 15079
rect 13820 15036 13872 15045
rect 13268 15011 13320 15020
rect 13268 14977 13277 15011
rect 13277 14977 13311 15011
rect 13311 14977 13320 15011
rect 13268 14968 13320 14977
rect 10140 14764 10192 14816
rect 13176 14900 13228 14952
rect 13728 14943 13780 14952
rect 13728 14909 13737 14943
rect 13737 14909 13771 14943
rect 13771 14909 13780 14943
rect 13728 14900 13780 14909
rect 14004 15011 14056 15020
rect 14004 14977 14013 15011
rect 14013 14977 14047 15011
rect 14047 14977 14056 15011
rect 14004 14968 14056 14977
rect 14188 15011 14240 15020
rect 14188 14977 14197 15011
rect 14197 14977 14231 15011
rect 14231 14977 14240 15011
rect 14188 14968 14240 14977
rect 15108 15079 15160 15088
rect 15108 15045 15117 15079
rect 15117 15045 15151 15079
rect 15151 15045 15160 15079
rect 15108 15036 15160 15045
rect 15200 15079 15252 15088
rect 15200 15045 15235 15079
rect 15235 15045 15252 15079
rect 15844 15104 15896 15156
rect 16856 15104 16908 15156
rect 15200 15036 15252 15045
rect 16304 15036 16356 15088
rect 17776 15147 17828 15156
rect 17776 15113 17785 15147
rect 17785 15113 17819 15147
rect 17819 15113 17828 15147
rect 17776 15104 17828 15113
rect 20352 15104 20404 15156
rect 14740 14900 14792 14952
rect 15384 14943 15436 14952
rect 15384 14909 15393 14943
rect 15393 14909 15427 14943
rect 15427 14909 15436 14943
rect 15384 14900 15436 14909
rect 15660 15011 15712 15020
rect 15660 14977 15669 15011
rect 15669 14977 15703 15011
rect 15703 14977 15712 15011
rect 15660 14968 15712 14977
rect 15752 14968 15804 15020
rect 17684 15036 17736 15088
rect 20168 15036 20220 15088
rect 12716 14832 12768 14884
rect 13360 14832 13412 14884
rect 13820 14832 13872 14884
rect 16396 14900 16448 14952
rect 16764 14968 16816 15020
rect 17960 15011 18012 15020
rect 17960 14977 17969 15011
rect 17969 14977 18003 15011
rect 18003 14977 18012 15011
rect 17960 14968 18012 14977
rect 18144 15011 18196 15020
rect 18144 14977 18153 15011
rect 18153 14977 18187 15011
rect 18187 14977 18196 15011
rect 18144 14968 18196 14977
rect 18236 14968 18288 15020
rect 18788 14968 18840 15020
rect 18972 14968 19024 15020
rect 20076 15011 20128 15020
rect 20076 14977 20085 15011
rect 20085 14977 20119 15011
rect 20119 14977 20128 15011
rect 20076 14968 20128 14977
rect 22284 15104 22336 15156
rect 24124 15104 24176 15156
rect 24492 15104 24544 15156
rect 24860 15147 24912 15156
rect 24860 15113 24869 15147
rect 24869 15113 24903 15147
rect 24903 15113 24912 15147
rect 24860 15104 24912 15113
rect 25136 15147 25188 15156
rect 25136 15113 25145 15147
rect 25145 15113 25179 15147
rect 25179 15113 25188 15147
rect 25136 15104 25188 15113
rect 20904 15011 20956 15020
rect 20904 14977 20913 15011
rect 20913 14977 20947 15011
rect 20947 14977 20956 15011
rect 20904 14968 20956 14977
rect 20996 14968 21048 15020
rect 21180 15011 21232 15020
rect 21180 14977 21189 15011
rect 21189 14977 21223 15011
rect 21223 14977 21232 15011
rect 21180 14968 21232 14977
rect 21272 15011 21324 15020
rect 21272 14977 21281 15011
rect 21281 14977 21315 15011
rect 21315 14977 21324 15011
rect 21272 14968 21324 14977
rect 21640 15011 21692 15020
rect 21640 14977 21649 15011
rect 21649 14977 21683 15011
rect 21683 14977 21692 15011
rect 21640 14968 21692 14977
rect 21824 15011 21876 15020
rect 21824 14977 21833 15011
rect 21833 14977 21867 15011
rect 21867 14977 21876 15011
rect 21824 14968 21876 14977
rect 15568 14832 15620 14884
rect 17224 14832 17276 14884
rect 18972 14832 19024 14884
rect 19432 14832 19484 14884
rect 22008 14968 22060 15020
rect 22284 15011 22336 15020
rect 22284 14977 22293 15011
rect 22293 14977 22327 15011
rect 22327 14977 22336 15011
rect 22284 14968 22336 14977
rect 23204 14968 23256 15020
rect 23940 15011 23992 15020
rect 23940 14977 23949 15011
rect 23949 14977 23983 15011
rect 23983 14977 23992 15011
rect 23940 14968 23992 14977
rect 24676 15011 24728 15020
rect 24676 14977 24688 15011
rect 24688 14977 24722 15011
rect 24722 14977 24728 15011
rect 24676 14968 24728 14977
rect 22284 14832 22336 14884
rect 12992 14764 13044 14816
rect 14372 14807 14424 14816
rect 14372 14773 14381 14807
rect 14381 14773 14415 14807
rect 14415 14773 14424 14807
rect 14372 14764 14424 14773
rect 15384 14764 15436 14816
rect 15844 14807 15896 14816
rect 15844 14773 15853 14807
rect 15853 14773 15887 14807
rect 15887 14773 15896 14807
rect 15844 14764 15896 14773
rect 16028 14807 16080 14816
rect 16028 14773 16037 14807
rect 16037 14773 16071 14807
rect 16071 14773 16080 14807
rect 16028 14764 16080 14773
rect 16672 14764 16724 14816
rect 18420 14764 18472 14816
rect 18880 14764 18932 14816
rect 20628 14764 20680 14816
rect 24308 14807 24360 14816
rect 24308 14773 24317 14807
rect 24317 14773 24351 14807
rect 24351 14773 24360 14807
rect 24308 14764 24360 14773
rect 24584 14764 24636 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 1952 14603 2004 14612
rect 1952 14569 1961 14603
rect 1961 14569 1995 14603
rect 1995 14569 2004 14603
rect 1952 14560 2004 14569
rect 4988 14560 5040 14612
rect 5356 14560 5408 14612
rect 2780 14492 2832 14544
rect 3700 14492 3752 14544
rect 3976 14492 4028 14544
rect 3240 14424 3292 14476
rect 7196 14492 7248 14544
rect 1860 14356 1912 14408
rect 2136 14356 2188 14408
rect 3608 14399 3660 14408
rect 3608 14365 3617 14399
rect 3617 14365 3651 14399
rect 3651 14365 3660 14399
rect 3608 14356 3660 14365
rect 7380 14424 7432 14476
rect 7748 14424 7800 14476
rect 10140 14560 10192 14612
rect 10968 14560 11020 14612
rect 12992 14560 13044 14612
rect 13176 14603 13228 14612
rect 13176 14569 13185 14603
rect 13185 14569 13219 14603
rect 13219 14569 13228 14603
rect 13176 14560 13228 14569
rect 8852 14492 8904 14544
rect 8668 14467 8720 14476
rect 8668 14433 8677 14467
rect 8677 14433 8711 14467
rect 8711 14433 8720 14467
rect 8668 14424 8720 14433
rect 9036 14424 9088 14476
rect 10784 14535 10836 14544
rect 10784 14501 10793 14535
rect 10793 14501 10827 14535
rect 10827 14501 10836 14535
rect 10784 14492 10836 14501
rect 14004 14560 14056 14612
rect 14188 14560 14240 14612
rect 16028 14560 16080 14612
rect 18144 14560 18196 14612
rect 21180 14560 21232 14612
rect 13728 14492 13780 14544
rect 4068 14399 4120 14408
rect 4068 14365 4077 14399
rect 4077 14365 4111 14399
rect 4111 14365 4120 14399
rect 4068 14356 4120 14365
rect 4988 14356 5040 14408
rect 7288 14356 7340 14408
rect 8576 14399 8628 14408
rect 8576 14365 8585 14399
rect 8585 14365 8619 14399
rect 8619 14365 8628 14399
rect 8576 14356 8628 14365
rect 1400 14288 1452 14340
rect 2872 14288 2924 14340
rect 9680 14399 9732 14408
rect 9680 14365 9689 14399
rect 9689 14365 9723 14399
rect 9723 14365 9732 14399
rect 9680 14356 9732 14365
rect 9772 14288 9824 14340
rect 10048 14331 10100 14340
rect 10048 14297 10057 14331
rect 10057 14297 10091 14331
rect 10091 14297 10100 14331
rect 10048 14288 10100 14297
rect 11244 14356 11296 14408
rect 12900 14424 12952 14476
rect 14372 14424 14424 14476
rect 14740 14424 14792 14476
rect 20168 14492 20220 14544
rect 24124 14560 24176 14612
rect 24492 14603 24544 14612
rect 24492 14569 24501 14603
rect 24501 14569 24535 14603
rect 24535 14569 24544 14603
rect 24492 14560 24544 14569
rect 22744 14492 22796 14544
rect 23112 14492 23164 14544
rect 12808 14399 12860 14408
rect 12808 14365 12817 14399
rect 12817 14365 12851 14399
rect 12851 14365 12860 14399
rect 12808 14356 12860 14365
rect 12992 14399 13044 14408
rect 12992 14365 13001 14399
rect 13001 14365 13035 14399
rect 13035 14365 13044 14399
rect 12992 14356 13044 14365
rect 1768 14220 1820 14272
rect 2228 14220 2280 14272
rect 3884 14220 3936 14272
rect 4804 14220 4856 14272
rect 5448 14220 5500 14272
rect 5632 14220 5684 14272
rect 8208 14263 8260 14272
rect 8208 14229 8217 14263
rect 8217 14229 8251 14263
rect 8251 14229 8260 14263
rect 8208 14220 8260 14229
rect 9496 14263 9548 14272
rect 9496 14229 9505 14263
rect 9505 14229 9539 14263
rect 9539 14229 9548 14263
rect 9496 14220 9548 14229
rect 12348 14288 12400 14340
rect 15016 14399 15068 14408
rect 15016 14365 15025 14399
rect 15025 14365 15059 14399
rect 15059 14365 15068 14399
rect 15016 14356 15068 14365
rect 15844 14356 15896 14408
rect 16672 14356 16724 14408
rect 20444 14424 20496 14476
rect 20628 14424 20680 14476
rect 10416 14263 10468 14272
rect 10416 14229 10425 14263
rect 10425 14229 10459 14263
rect 10459 14229 10468 14263
rect 10416 14220 10468 14229
rect 10692 14220 10744 14272
rect 17592 14288 17644 14340
rect 18420 14399 18472 14408
rect 18420 14365 18429 14399
rect 18429 14365 18463 14399
rect 18463 14365 18472 14399
rect 18420 14356 18472 14365
rect 18604 14399 18656 14408
rect 18604 14365 18613 14399
rect 18613 14365 18647 14399
rect 18647 14365 18656 14399
rect 18604 14356 18656 14365
rect 20904 14356 20956 14408
rect 21732 14399 21784 14408
rect 21732 14365 21741 14399
rect 21741 14365 21775 14399
rect 21775 14365 21784 14399
rect 21732 14356 21784 14365
rect 23940 14424 23992 14476
rect 22284 14399 22336 14408
rect 22284 14365 22293 14399
rect 22293 14365 22327 14399
rect 22327 14365 22336 14399
rect 22284 14356 22336 14365
rect 22560 14356 22612 14408
rect 20352 14288 20404 14340
rect 22008 14288 22060 14340
rect 22836 14288 22888 14340
rect 23204 14288 23256 14340
rect 26608 14399 26660 14408
rect 26608 14365 26617 14399
rect 26617 14365 26651 14399
rect 26651 14365 26660 14399
rect 26608 14356 26660 14365
rect 26700 14399 26752 14408
rect 26700 14365 26709 14399
rect 26709 14365 26743 14399
rect 26743 14365 26752 14399
rect 26700 14356 26752 14365
rect 14280 14220 14332 14272
rect 16028 14263 16080 14272
rect 16028 14229 16037 14263
rect 16037 14229 16071 14263
rect 16071 14229 16080 14263
rect 16028 14220 16080 14229
rect 18144 14220 18196 14272
rect 18236 14263 18288 14272
rect 18236 14229 18245 14263
rect 18245 14229 18279 14263
rect 18279 14229 18288 14263
rect 18236 14220 18288 14229
rect 18880 14220 18932 14272
rect 20812 14220 20864 14272
rect 21180 14220 21232 14272
rect 24124 14220 24176 14272
rect 4874 14118 4926 14170
rect 4938 14118 4990 14170
rect 5002 14118 5054 14170
rect 5066 14118 5118 14170
rect 5130 14118 5182 14170
rect 2136 14016 2188 14068
rect 2228 13948 2280 14000
rect 4068 13948 4120 14000
rect 1400 13923 1452 13932
rect 1400 13889 1409 13923
rect 1409 13889 1443 13923
rect 1443 13889 1452 13923
rect 1400 13880 1452 13889
rect 1492 13923 1544 13932
rect 1492 13889 1501 13923
rect 1501 13889 1535 13923
rect 1535 13889 1544 13923
rect 1492 13880 1544 13889
rect 1676 13923 1728 13932
rect 1676 13889 1685 13923
rect 1685 13889 1719 13923
rect 1719 13889 1728 13923
rect 1676 13880 1728 13889
rect 1768 13923 1820 13932
rect 1768 13889 1777 13923
rect 1777 13889 1811 13923
rect 1811 13889 1820 13923
rect 1768 13880 1820 13889
rect 2320 13880 2372 13932
rect 4712 14016 4764 14068
rect 4804 13991 4856 14000
rect 4804 13957 4813 13991
rect 4813 13957 4847 13991
rect 4847 13957 4856 13991
rect 4804 13948 4856 13957
rect 5908 14016 5960 14068
rect 6368 14059 6420 14068
rect 6368 14025 6377 14059
rect 6377 14025 6411 14059
rect 6411 14025 6420 14059
rect 6368 14016 6420 14025
rect 7656 14016 7708 14068
rect 8576 14016 8628 14068
rect 2044 13812 2096 13864
rect 2412 13855 2464 13864
rect 2412 13821 2421 13855
rect 2421 13821 2455 13855
rect 2455 13821 2464 13855
rect 2412 13812 2464 13821
rect 7656 13923 7708 13932
rect 7656 13889 7665 13923
rect 7665 13889 7699 13923
rect 7699 13889 7708 13923
rect 7656 13880 7708 13889
rect 9772 13948 9824 14000
rect 10692 13948 10744 14000
rect 13728 13948 13780 14000
rect 14096 13991 14148 14000
rect 14096 13957 14131 13991
rect 14131 13957 14148 13991
rect 16764 14016 16816 14068
rect 17960 14059 18012 14068
rect 14096 13948 14148 13957
rect 4620 13812 4672 13864
rect 5632 13812 5684 13864
rect 6092 13855 6144 13864
rect 6092 13821 6101 13855
rect 6101 13821 6135 13855
rect 6135 13821 6144 13855
rect 6092 13812 6144 13821
rect 5540 13744 5592 13796
rect 6920 13812 6972 13864
rect 9864 13812 9916 13864
rect 10508 13923 10560 13932
rect 10508 13889 10517 13923
rect 10517 13889 10551 13923
rect 10551 13889 10560 13923
rect 10508 13880 10560 13889
rect 7196 13744 7248 13796
rect 7840 13744 7892 13796
rect 8760 13744 8812 13796
rect 1676 13676 1728 13728
rect 3608 13676 3660 13728
rect 3976 13676 4028 13728
rect 4620 13676 4672 13728
rect 7932 13719 7984 13728
rect 7932 13685 7941 13719
rect 7941 13685 7975 13719
rect 7975 13685 7984 13719
rect 7932 13676 7984 13685
rect 8024 13719 8076 13728
rect 8024 13685 8033 13719
rect 8033 13685 8067 13719
rect 8067 13685 8076 13719
rect 8024 13676 8076 13685
rect 10140 13744 10192 13796
rect 10600 13812 10652 13864
rect 11060 13812 11112 13864
rect 12348 13880 12400 13932
rect 13452 13880 13504 13932
rect 13820 13923 13872 13932
rect 13820 13889 13829 13923
rect 13829 13889 13863 13923
rect 13863 13889 13872 13923
rect 13820 13880 13872 13889
rect 13912 13923 13964 13932
rect 13912 13889 13921 13923
rect 13921 13889 13955 13923
rect 13955 13889 13964 13923
rect 13912 13880 13964 13889
rect 14280 13923 14332 13932
rect 14280 13889 14289 13923
rect 14289 13889 14323 13923
rect 14323 13889 14332 13923
rect 14280 13880 14332 13889
rect 14556 13923 14608 13932
rect 14556 13889 14565 13923
rect 14565 13889 14599 13923
rect 14599 13889 14608 13923
rect 14556 13880 14608 13889
rect 16304 13948 16356 14000
rect 17224 13923 17276 13932
rect 17224 13889 17233 13923
rect 17233 13889 17267 13923
rect 17267 13889 17276 13923
rect 17224 13880 17276 13889
rect 17960 14025 17969 14059
rect 17969 14025 18003 14059
rect 18003 14025 18012 14059
rect 17960 14016 18012 14025
rect 18604 14016 18656 14068
rect 17592 13923 17644 13932
rect 17592 13889 17601 13923
rect 17601 13889 17635 13923
rect 17635 13889 17644 13923
rect 17592 13880 17644 13889
rect 17776 13880 17828 13932
rect 18144 13880 18196 13932
rect 19340 13948 19392 14000
rect 19156 13923 19208 13932
rect 19156 13889 19165 13923
rect 19165 13889 19199 13923
rect 19199 13889 19208 13923
rect 19156 13880 19208 13889
rect 19432 13957 19484 13966
rect 19432 13923 19441 13957
rect 19441 13923 19475 13957
rect 19475 13923 19484 13957
rect 19432 13914 19484 13923
rect 19892 13948 19944 14000
rect 20720 14016 20772 14068
rect 20996 14016 21048 14068
rect 21548 14016 21600 14068
rect 22560 14059 22612 14068
rect 22560 14025 22569 14059
rect 22569 14025 22603 14059
rect 22603 14025 22612 14059
rect 22560 14016 22612 14025
rect 26608 14016 26660 14068
rect 19616 13880 19668 13932
rect 9128 13676 9180 13728
rect 10324 13719 10376 13728
rect 10324 13685 10333 13719
rect 10333 13685 10367 13719
rect 10367 13685 10376 13719
rect 10324 13676 10376 13685
rect 13912 13676 13964 13728
rect 19432 13812 19484 13864
rect 19340 13744 19392 13796
rect 19524 13744 19576 13796
rect 20168 13880 20220 13932
rect 20352 13923 20404 13932
rect 20352 13889 20369 13923
rect 20369 13889 20403 13923
rect 20403 13889 20404 13923
rect 22928 13991 22980 14000
rect 22928 13957 22937 13991
rect 22937 13957 22971 13991
rect 22971 13957 22980 13991
rect 22928 13948 22980 13957
rect 20352 13880 20404 13889
rect 21180 13923 21232 13932
rect 21180 13889 21189 13923
rect 21189 13889 21223 13923
rect 21223 13889 21232 13923
rect 21180 13880 21232 13889
rect 21456 13923 21508 13932
rect 21456 13889 21465 13923
rect 21465 13889 21499 13923
rect 21499 13889 21508 13923
rect 21456 13880 21508 13889
rect 23020 13923 23072 13932
rect 23020 13889 23029 13923
rect 23029 13889 23063 13923
rect 23063 13889 23072 13923
rect 23020 13880 23072 13889
rect 23388 13923 23440 13932
rect 23388 13889 23397 13923
rect 23397 13889 23431 13923
rect 23431 13889 23440 13923
rect 23388 13880 23440 13889
rect 25044 13923 25096 13932
rect 25044 13889 25053 13923
rect 25053 13889 25087 13923
rect 25087 13889 25096 13923
rect 25044 13880 25096 13889
rect 25228 13923 25280 13932
rect 25228 13889 25237 13923
rect 25237 13889 25271 13923
rect 25271 13889 25280 13923
rect 25228 13880 25280 13889
rect 26424 13880 26476 13932
rect 23296 13812 23348 13864
rect 19800 13744 19852 13796
rect 14372 13719 14424 13728
rect 14372 13685 14381 13719
rect 14381 13685 14415 13719
rect 14415 13685 14424 13719
rect 14372 13676 14424 13685
rect 15844 13676 15896 13728
rect 16304 13719 16356 13728
rect 16304 13685 16313 13719
rect 16313 13685 16347 13719
rect 16347 13685 16356 13719
rect 16304 13676 16356 13685
rect 19432 13719 19484 13728
rect 19432 13685 19441 13719
rect 19441 13685 19475 13719
rect 19475 13685 19484 13719
rect 19432 13676 19484 13685
rect 22284 13744 22336 13796
rect 25412 13812 25464 13864
rect 25596 13855 25648 13864
rect 25596 13821 25605 13855
rect 25605 13821 25639 13855
rect 25639 13821 25648 13855
rect 25596 13812 25648 13821
rect 26240 13812 26292 13864
rect 26332 13855 26384 13864
rect 26332 13821 26341 13855
rect 26341 13821 26375 13855
rect 26375 13821 26384 13855
rect 26332 13812 26384 13821
rect 25780 13744 25832 13796
rect 20168 13676 20220 13728
rect 21272 13676 21324 13728
rect 26424 13676 26476 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 1676 13472 1728 13524
rect 5264 13472 5316 13524
rect 7932 13472 7984 13524
rect 8760 13472 8812 13524
rect 11060 13515 11112 13524
rect 11060 13481 11069 13515
rect 11069 13481 11103 13515
rect 11103 13481 11112 13515
rect 11060 13472 11112 13481
rect 1860 13447 1912 13456
rect 1860 13413 1869 13447
rect 1869 13413 1903 13447
rect 1903 13413 1912 13447
rect 1860 13404 1912 13413
rect 5540 13404 5592 13456
rect 7196 13447 7248 13456
rect 7196 13413 7205 13447
rect 7205 13413 7239 13447
rect 7239 13413 7248 13447
rect 7196 13404 7248 13413
rect 8024 13404 8076 13456
rect 1492 13268 1544 13320
rect 1400 13200 1452 13252
rect 2688 13200 2740 13252
rect 5632 13268 5684 13320
rect 10600 13336 10652 13388
rect 13820 13472 13872 13524
rect 14280 13515 14332 13524
rect 14280 13481 14289 13515
rect 14289 13481 14323 13515
rect 14323 13481 14332 13515
rect 14280 13472 14332 13481
rect 16396 13472 16448 13524
rect 19616 13472 19668 13524
rect 21180 13472 21232 13524
rect 22928 13515 22980 13524
rect 22928 13481 22937 13515
rect 22937 13481 22971 13515
rect 22971 13481 22980 13515
rect 22928 13472 22980 13481
rect 24124 13472 24176 13524
rect 25596 13472 25648 13524
rect 15384 13404 15436 13456
rect 8944 13311 8996 13320
rect 8944 13277 8953 13311
rect 8953 13277 8987 13311
rect 8987 13277 8996 13311
rect 8944 13268 8996 13277
rect 9128 13311 9180 13320
rect 9128 13277 9137 13311
rect 9137 13277 9171 13311
rect 9171 13277 9180 13311
rect 9128 13268 9180 13277
rect 9772 13268 9824 13320
rect 10140 13311 10192 13320
rect 10140 13277 10149 13311
rect 10149 13277 10183 13311
rect 10183 13277 10192 13311
rect 10140 13268 10192 13277
rect 10324 13311 10376 13320
rect 10324 13277 10333 13311
rect 10333 13277 10367 13311
rect 10367 13277 10376 13311
rect 10324 13268 10376 13277
rect 10508 13268 10560 13320
rect 14372 13311 14424 13320
rect 14372 13277 14381 13311
rect 14381 13277 14415 13311
rect 14415 13277 14424 13311
rect 14372 13268 14424 13277
rect 14556 13268 14608 13320
rect 16028 13336 16080 13388
rect 20628 13404 20680 13456
rect 19340 13336 19392 13388
rect 19432 13336 19484 13388
rect 20260 13379 20312 13388
rect 20260 13345 20269 13379
rect 20269 13345 20303 13379
rect 20303 13345 20312 13379
rect 20260 13336 20312 13345
rect 20352 13379 20404 13388
rect 20352 13345 20361 13379
rect 20361 13345 20395 13379
rect 20395 13345 20404 13379
rect 20352 13336 20404 13345
rect 3976 13132 4028 13184
rect 5264 13132 5316 13184
rect 7288 13175 7340 13184
rect 7288 13141 7297 13175
rect 7297 13141 7331 13175
rect 7331 13141 7340 13175
rect 7288 13132 7340 13141
rect 7656 13175 7708 13184
rect 7656 13141 7665 13175
rect 7665 13141 7699 13175
rect 7699 13141 7708 13175
rect 7656 13132 7708 13141
rect 8116 13132 8168 13184
rect 9036 13175 9088 13184
rect 9036 13141 9045 13175
rect 9045 13141 9079 13175
rect 9079 13141 9088 13175
rect 9036 13132 9088 13141
rect 10140 13175 10192 13184
rect 10140 13141 10149 13175
rect 10149 13141 10183 13175
rect 10183 13141 10192 13175
rect 10140 13132 10192 13141
rect 10692 13132 10744 13184
rect 11796 13175 11848 13184
rect 11796 13141 11805 13175
rect 11805 13141 11839 13175
rect 11839 13141 11848 13175
rect 11796 13132 11848 13141
rect 14556 13175 14608 13184
rect 14556 13141 14565 13175
rect 14565 13141 14599 13175
rect 14599 13141 14608 13175
rect 14556 13132 14608 13141
rect 15292 13311 15344 13320
rect 15292 13277 15301 13311
rect 15301 13277 15335 13311
rect 15335 13277 15344 13311
rect 15292 13268 15344 13277
rect 14832 13243 14884 13252
rect 14832 13209 14841 13243
rect 14841 13209 14875 13243
rect 14875 13209 14884 13243
rect 14832 13200 14884 13209
rect 15108 13200 15160 13252
rect 16304 13311 16356 13320
rect 16304 13277 16313 13311
rect 16313 13277 16347 13311
rect 16347 13277 16356 13311
rect 16304 13268 16356 13277
rect 19156 13268 19208 13320
rect 19708 13268 19760 13320
rect 21272 13404 21324 13456
rect 15752 13200 15804 13252
rect 19340 13200 19392 13252
rect 20168 13200 20220 13252
rect 16948 13132 17000 13184
rect 19524 13132 19576 13184
rect 20996 13268 21048 13320
rect 21456 13311 21508 13320
rect 21456 13277 21465 13311
rect 21465 13277 21499 13311
rect 21499 13277 21508 13311
rect 21456 13268 21508 13277
rect 25320 13404 25372 13456
rect 26148 13404 26200 13456
rect 25780 13336 25832 13388
rect 26332 13336 26384 13388
rect 20628 13200 20680 13252
rect 20536 13132 20588 13184
rect 22928 13175 22980 13184
rect 22928 13141 22955 13175
rect 22955 13141 22980 13175
rect 22928 13132 22980 13141
rect 23296 13200 23348 13252
rect 23848 13200 23900 13252
rect 24768 13200 24820 13252
rect 24952 13200 25004 13252
rect 26148 13311 26200 13320
rect 26148 13277 26157 13311
rect 26157 13277 26191 13311
rect 26191 13277 26200 13311
rect 26148 13268 26200 13277
rect 26700 13200 26752 13252
rect 23388 13132 23440 13184
rect 4874 13030 4926 13082
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 10324 12928 10376 12980
rect 14832 12971 14884 12980
rect 14832 12937 14841 12971
rect 14841 12937 14875 12971
rect 14875 12937 14884 12971
rect 14832 12928 14884 12937
rect 2688 12792 2740 12844
rect 3792 12835 3844 12844
rect 3792 12801 3801 12835
rect 3801 12801 3835 12835
rect 3835 12801 3844 12835
rect 3792 12792 3844 12801
rect 3976 12835 4028 12844
rect 3976 12801 3985 12835
rect 3985 12801 4019 12835
rect 4019 12801 4028 12835
rect 3976 12792 4028 12801
rect 5540 12792 5592 12844
rect 8024 12792 8076 12844
rect 8392 12835 8444 12844
rect 8392 12801 8401 12835
rect 8401 12801 8435 12835
rect 8435 12801 8444 12835
rect 10784 12860 10836 12912
rect 15752 12928 15804 12980
rect 15384 12860 15436 12912
rect 8392 12792 8444 12801
rect 10140 12835 10192 12844
rect 10140 12801 10149 12835
rect 10149 12801 10183 12835
rect 10183 12801 10192 12835
rect 10140 12792 10192 12801
rect 10324 12835 10376 12844
rect 10324 12801 10333 12835
rect 10333 12801 10367 12835
rect 10367 12801 10376 12835
rect 10324 12792 10376 12801
rect 10416 12835 10468 12844
rect 10416 12801 10425 12835
rect 10425 12801 10459 12835
rect 10459 12801 10468 12835
rect 10416 12792 10468 12801
rect 4068 12724 4120 12776
rect 6368 12767 6420 12776
rect 6368 12733 6377 12767
rect 6377 12733 6411 12767
rect 6411 12733 6420 12767
rect 6368 12724 6420 12733
rect 6920 12767 6972 12776
rect 6920 12733 6929 12767
rect 6929 12733 6963 12767
rect 6963 12733 6972 12767
rect 6920 12724 6972 12733
rect 10692 12835 10744 12844
rect 10692 12801 10701 12835
rect 10701 12801 10735 12835
rect 10735 12801 10744 12835
rect 10692 12792 10744 12801
rect 3792 12656 3844 12708
rect 5356 12656 5408 12708
rect 8392 12656 8444 12708
rect 13544 12835 13596 12844
rect 13544 12801 13553 12835
rect 13553 12801 13587 12835
rect 13587 12801 13596 12835
rect 13544 12792 13596 12801
rect 14556 12792 14608 12844
rect 15292 12792 15344 12844
rect 14004 12724 14056 12776
rect 14648 12767 14700 12776
rect 14648 12733 14657 12767
rect 14657 12733 14691 12767
rect 14691 12733 14700 12767
rect 14648 12724 14700 12733
rect 15660 12903 15712 12912
rect 15660 12869 15669 12903
rect 15669 12869 15703 12903
rect 15703 12869 15712 12903
rect 15660 12860 15712 12869
rect 19156 12928 19208 12980
rect 20352 12928 20404 12980
rect 20720 12928 20772 12980
rect 14096 12656 14148 12708
rect 16120 12724 16172 12776
rect 16304 12835 16356 12844
rect 16304 12801 16313 12835
rect 16313 12801 16347 12835
rect 16347 12801 16356 12835
rect 16304 12792 16356 12801
rect 16948 12835 17000 12844
rect 16948 12801 16957 12835
rect 16957 12801 16991 12835
rect 16991 12801 17000 12835
rect 16948 12792 17000 12801
rect 16396 12724 16448 12776
rect 17316 12767 17368 12776
rect 17316 12733 17325 12767
rect 17325 12733 17359 12767
rect 17359 12733 17368 12767
rect 17316 12724 17368 12733
rect 17868 12767 17920 12776
rect 17868 12733 17877 12767
rect 17877 12733 17911 12767
rect 17911 12733 17920 12767
rect 17868 12724 17920 12733
rect 18880 12835 18932 12844
rect 18880 12801 18889 12835
rect 18889 12801 18923 12835
rect 18923 12801 18932 12835
rect 18880 12792 18932 12801
rect 19340 12860 19392 12912
rect 19708 12860 19760 12912
rect 23848 12860 23900 12912
rect 24860 12928 24912 12980
rect 24676 12860 24728 12912
rect 26332 12928 26384 12980
rect 20260 12792 20312 12844
rect 21824 12792 21876 12844
rect 26240 12860 26292 12912
rect 26608 12903 26660 12912
rect 26608 12869 26617 12903
rect 26617 12869 26651 12903
rect 26651 12869 26660 12903
rect 26608 12860 26660 12869
rect 15108 12656 15160 12708
rect 17776 12656 17828 12708
rect 20536 12767 20588 12776
rect 20536 12733 20545 12767
rect 20545 12733 20579 12767
rect 20579 12733 20588 12767
rect 20536 12724 20588 12733
rect 20628 12656 20680 12708
rect 4620 12588 4672 12640
rect 7932 12631 7984 12640
rect 7932 12597 7941 12631
rect 7941 12597 7975 12631
rect 7975 12597 7984 12631
rect 7932 12588 7984 12597
rect 8116 12631 8168 12640
rect 8116 12597 8125 12631
rect 8125 12597 8159 12631
rect 8159 12597 8168 12631
rect 8116 12588 8168 12597
rect 10876 12631 10928 12640
rect 10876 12597 10885 12631
rect 10885 12597 10919 12631
rect 10919 12597 10928 12631
rect 10876 12588 10928 12597
rect 11244 12631 11296 12640
rect 11244 12597 11253 12631
rect 11253 12597 11287 12631
rect 11287 12597 11296 12631
rect 11244 12588 11296 12597
rect 13176 12631 13228 12640
rect 13176 12597 13185 12631
rect 13185 12597 13219 12631
rect 13219 12597 13228 12631
rect 13176 12588 13228 12597
rect 15292 12631 15344 12640
rect 15292 12597 15301 12631
rect 15301 12597 15335 12631
rect 15335 12597 15344 12631
rect 15292 12588 15344 12597
rect 20444 12588 20496 12640
rect 24860 12724 24912 12776
rect 25688 12835 25740 12844
rect 25688 12801 25697 12835
rect 25697 12801 25731 12835
rect 25731 12801 25740 12835
rect 25688 12792 25740 12801
rect 26148 12792 26200 12844
rect 26700 12792 26752 12844
rect 26056 12724 26108 12776
rect 25780 12656 25832 12708
rect 24400 12588 24452 12640
rect 24676 12588 24728 12640
rect 24768 12631 24820 12640
rect 24768 12597 24777 12631
rect 24777 12597 24811 12631
rect 24811 12597 24820 12631
rect 24768 12588 24820 12597
rect 24952 12588 25004 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 4252 12427 4304 12436
rect 4252 12393 4261 12427
rect 4261 12393 4295 12427
rect 4295 12393 4304 12427
rect 4252 12384 4304 12393
rect 3700 12316 3752 12368
rect 5356 12316 5408 12368
rect 4068 12248 4120 12300
rect 2136 12223 2188 12232
rect 2136 12189 2145 12223
rect 2145 12189 2179 12223
rect 2179 12189 2188 12223
rect 2136 12180 2188 12189
rect 2320 12180 2372 12232
rect 2504 12180 2556 12232
rect 1676 12044 1728 12096
rect 2872 12223 2924 12232
rect 2872 12189 2881 12223
rect 2881 12189 2915 12223
rect 2915 12189 2924 12223
rect 2872 12180 2924 12189
rect 3792 12223 3844 12232
rect 3792 12189 3801 12223
rect 3801 12189 3835 12223
rect 3835 12189 3844 12223
rect 3792 12180 3844 12189
rect 4160 12112 4212 12164
rect 4712 12248 4764 12300
rect 3240 12044 3292 12096
rect 4620 12180 4672 12232
rect 5356 12223 5408 12232
rect 5356 12189 5365 12223
rect 5365 12189 5399 12223
rect 5399 12189 5408 12223
rect 5356 12180 5408 12189
rect 6736 12384 6788 12436
rect 7288 12248 7340 12300
rect 8024 12384 8076 12436
rect 8392 12384 8444 12436
rect 8576 12384 8628 12436
rect 7012 12223 7064 12232
rect 7012 12189 7021 12223
rect 7021 12189 7055 12223
rect 7055 12189 7064 12223
rect 7012 12180 7064 12189
rect 7380 12223 7432 12232
rect 7380 12189 7389 12223
rect 7389 12189 7423 12223
rect 7423 12189 7432 12223
rect 7380 12180 7432 12189
rect 7564 12223 7616 12232
rect 7564 12189 7573 12223
rect 7573 12189 7607 12223
rect 7607 12189 7616 12223
rect 7564 12180 7616 12189
rect 8208 12248 8260 12300
rect 8392 12223 8444 12232
rect 8392 12189 8401 12223
rect 8401 12189 8435 12223
rect 8435 12189 8444 12223
rect 8392 12180 8444 12189
rect 8668 12223 8720 12232
rect 8668 12189 8677 12223
rect 8677 12189 8711 12223
rect 8711 12189 8720 12223
rect 8668 12180 8720 12189
rect 9128 12316 9180 12368
rect 9772 12384 9824 12436
rect 16120 12384 16172 12436
rect 17316 12384 17368 12436
rect 19616 12427 19668 12436
rect 19616 12393 19625 12427
rect 19625 12393 19659 12427
rect 19659 12393 19668 12427
rect 19616 12384 19668 12393
rect 20628 12384 20680 12436
rect 21732 12384 21784 12436
rect 25780 12384 25832 12436
rect 9496 12180 9548 12232
rect 9772 12223 9824 12232
rect 9772 12189 9781 12223
rect 9781 12189 9815 12223
rect 9815 12189 9824 12223
rect 9772 12180 9824 12189
rect 9036 12112 9088 12164
rect 10232 12180 10284 12232
rect 10784 12180 10836 12232
rect 11612 12223 11664 12232
rect 11612 12189 11621 12223
rect 11621 12189 11655 12223
rect 11655 12189 11664 12223
rect 11612 12180 11664 12189
rect 11796 12223 11848 12232
rect 11796 12189 11805 12223
rect 11805 12189 11839 12223
rect 11839 12189 11848 12223
rect 11796 12180 11848 12189
rect 12164 12223 12216 12232
rect 12164 12189 12173 12223
rect 12173 12189 12207 12223
rect 12207 12189 12216 12223
rect 12164 12180 12216 12189
rect 15476 12291 15528 12300
rect 15476 12257 15485 12291
rect 15485 12257 15519 12291
rect 15519 12257 15528 12291
rect 15476 12248 15528 12257
rect 15292 12180 15344 12232
rect 17224 12180 17276 12232
rect 17776 12223 17828 12232
rect 17776 12189 17785 12223
rect 17785 12189 17819 12223
rect 17819 12189 17828 12223
rect 17776 12180 17828 12189
rect 18236 12180 18288 12232
rect 4804 12087 4856 12096
rect 4804 12053 4813 12087
rect 4813 12053 4847 12087
rect 4847 12053 4856 12087
rect 4804 12044 4856 12053
rect 6828 12044 6880 12096
rect 7012 12044 7064 12096
rect 8024 12044 8076 12096
rect 8116 12087 8168 12096
rect 8116 12053 8125 12087
rect 8125 12053 8159 12087
rect 8159 12053 8168 12087
rect 8116 12044 8168 12053
rect 11336 12044 11388 12096
rect 12440 12044 12492 12096
rect 12624 12044 12676 12096
rect 24492 12248 24544 12300
rect 27160 12316 27212 12368
rect 25688 12248 25740 12300
rect 23020 12223 23072 12232
rect 23020 12189 23029 12223
rect 23029 12189 23063 12223
rect 23063 12189 23072 12223
rect 23020 12180 23072 12189
rect 23204 12223 23256 12232
rect 23204 12189 23213 12223
rect 23213 12189 23247 12223
rect 23247 12189 23256 12223
rect 23204 12180 23256 12189
rect 23388 12223 23440 12232
rect 23388 12189 23397 12223
rect 23397 12189 23431 12223
rect 23431 12189 23440 12223
rect 23388 12180 23440 12189
rect 25504 12223 25556 12232
rect 25504 12189 25513 12223
rect 25513 12189 25547 12223
rect 25547 12189 25556 12223
rect 25504 12180 25556 12189
rect 25964 12180 26016 12232
rect 24032 12112 24084 12164
rect 25228 12112 25280 12164
rect 22928 12044 22980 12096
rect 23940 12044 23992 12096
rect 25412 12087 25464 12096
rect 25412 12053 25421 12087
rect 25421 12053 25455 12087
rect 25455 12053 25464 12087
rect 25412 12044 25464 12053
rect 25688 12044 25740 12096
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 2504 11840 2556 11892
rect 2412 11772 2464 11824
rect 1676 11747 1728 11756
rect 1676 11713 1710 11747
rect 1710 11713 1728 11747
rect 1676 11704 1728 11713
rect 12164 11840 12216 11892
rect 14648 11883 14700 11892
rect 14648 11849 14657 11883
rect 14657 11849 14691 11883
rect 14691 11849 14700 11883
rect 14648 11840 14700 11849
rect 19984 11840 20036 11892
rect 23204 11840 23256 11892
rect 24492 11840 24544 11892
rect 24860 11840 24912 11892
rect 3240 11679 3292 11688
rect 3240 11645 3249 11679
rect 3249 11645 3283 11679
rect 3283 11645 3292 11679
rect 3240 11636 3292 11645
rect 3884 11747 3936 11756
rect 3884 11713 3893 11747
rect 3893 11713 3927 11747
rect 3927 11713 3936 11747
rect 3884 11704 3936 11713
rect 4160 11704 4212 11756
rect 5172 11704 5224 11756
rect 5356 11772 5408 11824
rect 8116 11772 8168 11824
rect 5540 11747 5592 11756
rect 5540 11713 5549 11747
rect 5549 11713 5583 11747
rect 5583 11713 5592 11747
rect 5540 11704 5592 11713
rect 5724 11747 5776 11756
rect 5724 11713 5733 11747
rect 5733 11713 5767 11747
rect 5767 11713 5776 11747
rect 5724 11704 5776 11713
rect 4804 11636 4856 11688
rect 3516 11611 3568 11620
rect 3516 11577 3525 11611
rect 3525 11577 3559 11611
rect 3559 11577 3568 11611
rect 3516 11568 3568 11577
rect 6184 11500 6236 11552
rect 6644 11704 6696 11756
rect 6920 11747 6972 11756
rect 6920 11713 6929 11747
rect 6929 11713 6963 11747
rect 6963 11713 6972 11747
rect 6920 11704 6972 11713
rect 6828 11636 6880 11688
rect 6552 11568 6604 11620
rect 8668 11704 8720 11756
rect 9128 11747 9180 11756
rect 9128 11713 9137 11747
rect 9137 11713 9171 11747
rect 9171 11713 9180 11747
rect 9128 11704 9180 11713
rect 9404 11704 9456 11756
rect 7472 11636 7524 11688
rect 10324 11747 10376 11756
rect 10324 11713 10333 11747
rect 10333 11713 10367 11747
rect 10367 11713 10376 11747
rect 10324 11704 10376 11713
rect 10784 11704 10836 11756
rect 11704 11704 11756 11756
rect 11796 11747 11848 11756
rect 11796 11713 11805 11747
rect 11805 11713 11839 11747
rect 11839 11713 11848 11747
rect 11796 11704 11848 11713
rect 13176 11772 13228 11824
rect 18052 11772 18104 11824
rect 19248 11772 19300 11824
rect 23020 11772 23072 11824
rect 23940 11815 23992 11824
rect 23940 11781 23949 11815
rect 23949 11781 23983 11815
rect 23983 11781 23992 11815
rect 23940 11772 23992 11781
rect 25412 11815 25464 11824
rect 25412 11781 25421 11815
rect 25421 11781 25455 11815
rect 25455 11781 25464 11815
rect 25412 11772 25464 11781
rect 12440 11747 12492 11756
rect 10968 11636 11020 11688
rect 11520 11636 11572 11688
rect 12440 11713 12449 11747
rect 12449 11713 12483 11747
rect 12483 11713 12492 11747
rect 12440 11704 12492 11713
rect 12624 11747 12676 11756
rect 12624 11713 12633 11747
rect 12633 11713 12667 11747
rect 12667 11713 12676 11747
rect 12624 11704 12676 11713
rect 13360 11704 13412 11756
rect 18604 11747 18656 11756
rect 18604 11713 18613 11747
rect 18613 11713 18647 11747
rect 18647 11713 18656 11747
rect 18604 11704 18656 11713
rect 20536 11704 20588 11756
rect 23480 11747 23532 11756
rect 23480 11713 23489 11747
rect 23489 11713 23523 11747
rect 23523 11713 23532 11747
rect 23480 11704 23532 11713
rect 24400 11747 24452 11756
rect 24400 11713 24409 11747
rect 24409 11713 24443 11747
rect 24443 11713 24452 11747
rect 24400 11704 24452 11713
rect 24952 11704 25004 11756
rect 25504 11704 25556 11756
rect 27160 11747 27212 11756
rect 27160 11713 27169 11747
rect 27169 11713 27203 11747
rect 27203 11713 27212 11747
rect 27160 11704 27212 11713
rect 27252 11747 27304 11756
rect 27252 11713 27261 11747
rect 27261 11713 27295 11747
rect 27295 11713 27304 11747
rect 27252 11704 27304 11713
rect 20904 11679 20956 11688
rect 20904 11645 20913 11679
rect 20913 11645 20947 11679
rect 20947 11645 20956 11679
rect 20904 11636 20956 11645
rect 22744 11636 22796 11688
rect 23572 11636 23624 11688
rect 23848 11679 23900 11688
rect 23848 11645 23857 11679
rect 23857 11645 23891 11679
rect 23891 11645 23900 11679
rect 23848 11636 23900 11645
rect 26056 11679 26108 11688
rect 26056 11645 26065 11679
rect 26065 11645 26099 11679
rect 26099 11645 26108 11679
rect 26056 11636 26108 11645
rect 12532 11568 12584 11620
rect 25688 11611 25740 11620
rect 25688 11577 25697 11611
rect 25697 11577 25731 11611
rect 25731 11577 25740 11611
rect 25688 11568 25740 11577
rect 7932 11500 7984 11552
rect 8208 11500 8260 11552
rect 11612 11500 11664 11552
rect 12624 11500 12676 11552
rect 23388 11500 23440 11552
rect 26516 11543 26568 11552
rect 26516 11509 26525 11543
rect 26525 11509 26559 11543
rect 26559 11509 26568 11543
rect 26516 11500 26568 11509
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 4804 11339 4856 11348
rect 4804 11305 4813 11339
rect 4813 11305 4847 11339
rect 4847 11305 4856 11339
rect 4804 11296 4856 11305
rect 8300 11339 8352 11348
rect 8300 11305 8309 11339
rect 8309 11305 8343 11339
rect 8343 11305 8352 11339
rect 8300 11296 8352 11305
rect 8392 11296 8444 11348
rect 8576 11296 8628 11348
rect 7564 11160 7616 11212
rect 8208 11228 8260 11280
rect 4344 11092 4396 11144
rect 4620 11092 4672 11144
rect 4804 11092 4856 11144
rect 5172 11092 5224 11144
rect 5540 11135 5592 11144
rect 5540 11101 5549 11135
rect 5549 11101 5583 11135
rect 5583 11101 5592 11135
rect 5540 11092 5592 11101
rect 5724 11135 5776 11144
rect 5724 11101 5733 11135
rect 5733 11101 5767 11135
rect 5767 11101 5776 11135
rect 5724 11092 5776 11101
rect 6552 11024 6604 11076
rect 4712 10956 4764 11008
rect 4896 10956 4948 11008
rect 5356 10956 5408 11008
rect 8392 11135 8444 11144
rect 8392 11101 8401 11135
rect 8401 11101 8435 11135
rect 8435 11101 8444 11135
rect 8392 11092 8444 11101
rect 9036 11203 9088 11212
rect 9036 11169 9045 11203
rect 9045 11169 9079 11203
rect 9079 11169 9088 11203
rect 9036 11160 9088 11169
rect 9404 11092 9456 11144
rect 11704 11296 11756 11348
rect 19248 11339 19300 11348
rect 19248 11305 19257 11339
rect 19257 11305 19291 11339
rect 19291 11305 19300 11339
rect 19248 11296 19300 11305
rect 23112 11296 23164 11348
rect 24308 11296 24360 11348
rect 26056 11296 26108 11348
rect 15476 11228 15528 11280
rect 12624 11160 12676 11212
rect 9036 11024 9088 11076
rect 9772 11067 9824 11076
rect 9772 11033 9781 11067
rect 9781 11033 9815 11067
rect 9815 11033 9824 11067
rect 9772 11024 9824 11033
rect 8300 10956 8352 11008
rect 9128 10956 9180 11008
rect 10876 11092 10928 11144
rect 10968 11092 11020 11144
rect 11336 11135 11388 11144
rect 11336 11101 11345 11135
rect 11345 11101 11379 11135
rect 11379 11101 11388 11135
rect 11336 11092 11388 11101
rect 12532 11135 12584 11144
rect 12532 11101 12541 11135
rect 12541 11101 12575 11135
rect 12575 11101 12584 11135
rect 12532 11092 12584 11101
rect 12992 11203 13044 11212
rect 12992 11169 13001 11203
rect 13001 11169 13035 11203
rect 13035 11169 13044 11203
rect 12992 11160 13044 11169
rect 14924 11160 14976 11212
rect 16120 11160 16172 11212
rect 11796 11024 11848 11076
rect 14188 11092 14240 11144
rect 14832 11092 14884 11144
rect 15108 11092 15160 11144
rect 17132 11092 17184 11144
rect 17500 11092 17552 11144
rect 17776 11135 17828 11144
rect 16212 11024 16264 11076
rect 17776 11101 17798 11135
rect 17798 11101 17828 11135
rect 17776 11092 17828 11101
rect 18052 11135 18104 11144
rect 10324 10956 10376 11008
rect 12716 10956 12768 11008
rect 13912 10999 13964 11008
rect 13912 10965 13921 10999
rect 13921 10965 13955 10999
rect 13955 10965 13964 10999
rect 13912 10956 13964 10965
rect 18052 11101 18061 11135
rect 18061 11101 18095 11135
rect 18095 11101 18104 11135
rect 18052 11092 18104 11101
rect 23480 11160 23532 11212
rect 23756 11160 23808 11212
rect 27160 11228 27212 11280
rect 18604 11092 18656 11144
rect 19892 11092 19944 11144
rect 22376 11135 22428 11144
rect 22376 11101 22385 11135
rect 22385 11101 22419 11135
rect 22419 11101 22428 11135
rect 22376 11092 22428 11101
rect 24584 11092 24636 11144
rect 26608 11160 26660 11212
rect 27252 11160 27304 11212
rect 25412 11092 25464 11144
rect 19340 11024 19392 11076
rect 21180 11024 21232 11076
rect 19800 10956 19852 11008
rect 22284 10999 22336 11008
rect 22284 10965 22293 10999
rect 22293 10965 22327 10999
rect 22327 10965 22336 10999
rect 22284 10956 22336 10965
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 3516 10752 3568 10804
rect 3884 10684 3936 10736
rect 9036 10684 9088 10736
rect 18604 10752 18656 10804
rect 20352 10752 20404 10804
rect 20904 10752 20956 10804
rect 4160 10591 4212 10600
rect 4160 10557 4169 10591
rect 4169 10557 4203 10591
rect 4203 10557 4212 10591
rect 4160 10548 4212 10557
rect 4804 10616 4856 10668
rect 5264 10616 5316 10668
rect 6644 10659 6696 10668
rect 6644 10625 6653 10659
rect 6653 10625 6687 10659
rect 6687 10625 6696 10659
rect 6644 10616 6696 10625
rect 7472 10616 7524 10668
rect 9128 10659 9180 10668
rect 9128 10625 9137 10659
rect 9137 10625 9171 10659
rect 9171 10625 9180 10659
rect 9128 10616 9180 10625
rect 9312 10659 9364 10668
rect 9312 10625 9321 10659
rect 9321 10625 9355 10659
rect 9355 10625 9364 10659
rect 9312 10616 9364 10625
rect 9496 10659 9548 10668
rect 9496 10625 9505 10659
rect 9505 10625 9539 10659
rect 9539 10625 9548 10659
rect 9496 10616 9548 10625
rect 12348 10659 12400 10668
rect 12348 10625 12357 10659
rect 12357 10625 12391 10659
rect 12391 10625 12400 10659
rect 12348 10616 12400 10625
rect 12440 10659 12492 10668
rect 12440 10625 12449 10659
rect 12449 10625 12483 10659
rect 12483 10625 12492 10659
rect 12440 10616 12492 10625
rect 12624 10659 12676 10668
rect 12624 10625 12633 10659
rect 12633 10625 12667 10659
rect 12667 10625 12676 10659
rect 12624 10616 12676 10625
rect 12716 10659 12768 10668
rect 12716 10625 12725 10659
rect 12725 10625 12759 10659
rect 12759 10625 12768 10659
rect 12716 10616 12768 10625
rect 4344 10480 4396 10532
rect 5356 10548 5408 10600
rect 6276 10548 6328 10600
rect 8392 10548 8444 10600
rect 15476 10616 15528 10668
rect 16212 10616 16264 10668
rect 16488 10616 16540 10668
rect 17040 10659 17092 10668
rect 17040 10625 17049 10659
rect 17049 10625 17083 10659
rect 17083 10625 17092 10659
rect 17040 10616 17092 10625
rect 15384 10548 15436 10600
rect 16764 10548 16816 10600
rect 17776 10727 17828 10736
rect 17776 10693 17811 10727
rect 17811 10693 17828 10727
rect 17776 10684 17828 10693
rect 17960 10727 18012 10736
rect 17960 10693 17985 10727
rect 17985 10693 18012 10727
rect 17960 10684 18012 10693
rect 19708 10684 19760 10736
rect 17684 10659 17736 10668
rect 17684 10625 17693 10659
rect 17693 10625 17727 10659
rect 17727 10625 17736 10659
rect 17684 10616 17736 10625
rect 19800 10616 19852 10668
rect 20536 10616 20588 10668
rect 21088 10616 21140 10668
rect 21456 10616 21508 10668
rect 22008 10659 22060 10668
rect 22008 10625 22017 10659
rect 22017 10625 22051 10659
rect 22051 10625 22060 10659
rect 22008 10616 22060 10625
rect 22192 10616 22244 10668
rect 22560 10616 22612 10668
rect 25688 10727 25740 10736
rect 25688 10693 25697 10727
rect 25697 10693 25731 10727
rect 25731 10693 25740 10727
rect 25688 10684 25740 10693
rect 24216 10616 24268 10668
rect 24308 10659 24360 10668
rect 24308 10625 24317 10659
rect 24317 10625 24351 10659
rect 24351 10625 24360 10659
rect 24308 10616 24360 10625
rect 24492 10659 24544 10668
rect 24492 10625 24501 10659
rect 24501 10625 24535 10659
rect 24535 10625 24544 10659
rect 24492 10616 24544 10625
rect 24676 10659 24728 10668
rect 24676 10625 24685 10659
rect 24685 10625 24719 10659
rect 24719 10625 24728 10659
rect 24676 10616 24728 10625
rect 12992 10480 13044 10532
rect 17316 10480 17368 10532
rect 4620 10412 4672 10464
rect 7196 10412 7248 10464
rect 9864 10412 9916 10464
rect 11796 10412 11848 10464
rect 17500 10412 17552 10464
rect 19340 10548 19392 10600
rect 19892 10548 19944 10600
rect 21180 10591 21232 10600
rect 21180 10557 21189 10591
rect 21189 10557 21223 10591
rect 21223 10557 21232 10591
rect 21180 10548 21232 10557
rect 21824 10591 21876 10600
rect 21824 10557 21833 10591
rect 21833 10557 21867 10591
rect 21867 10557 21876 10591
rect 21824 10548 21876 10557
rect 22836 10548 22888 10600
rect 19524 10412 19576 10464
rect 19984 10412 20036 10464
rect 20444 10412 20496 10464
rect 20628 10455 20680 10464
rect 20628 10421 20637 10455
rect 20637 10421 20671 10455
rect 20671 10421 20680 10455
rect 20628 10412 20680 10421
rect 21640 10412 21692 10464
rect 22284 10412 22336 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 6276 10251 6328 10260
rect 6276 10217 6285 10251
rect 6285 10217 6319 10251
rect 6319 10217 6328 10251
rect 6276 10208 6328 10217
rect 11888 10251 11940 10260
rect 11888 10217 11897 10251
rect 11897 10217 11931 10251
rect 11931 10217 11940 10251
rect 11888 10208 11940 10217
rect 15108 10208 15160 10260
rect 15476 10251 15528 10260
rect 15476 10217 15485 10251
rect 15485 10217 15519 10251
rect 15519 10217 15528 10251
rect 15476 10208 15528 10217
rect 16764 10251 16816 10260
rect 16764 10217 16773 10251
rect 16773 10217 16807 10251
rect 16807 10217 16816 10251
rect 16764 10208 16816 10217
rect 17040 10208 17092 10260
rect 19524 10208 19576 10260
rect 21272 10208 21324 10260
rect 21824 10251 21876 10260
rect 21824 10217 21833 10251
rect 21833 10217 21867 10251
rect 21867 10217 21876 10251
rect 21824 10208 21876 10217
rect 4712 10004 4764 10056
rect 5540 10072 5592 10124
rect 5908 10004 5960 10056
rect 7472 10072 7524 10124
rect 9312 10115 9364 10124
rect 9312 10081 9321 10115
rect 9321 10081 9355 10115
rect 9355 10081 9364 10115
rect 9312 10072 9364 10081
rect 6828 10047 6880 10056
rect 6828 10013 6837 10047
rect 6837 10013 6871 10047
rect 6871 10013 6880 10047
rect 6828 10004 6880 10013
rect 6184 9936 6236 9988
rect 6552 9979 6604 9988
rect 6552 9945 6561 9979
rect 6561 9945 6595 9979
rect 6595 9945 6604 9979
rect 6552 9936 6604 9945
rect 6644 9979 6696 9988
rect 6644 9945 6653 9979
rect 6653 9945 6687 9979
rect 6687 9945 6696 9979
rect 6644 9936 6696 9945
rect 8208 10047 8260 10056
rect 8208 10013 8217 10047
rect 8217 10013 8251 10047
rect 8251 10013 8260 10047
rect 8208 10004 8260 10013
rect 9496 10004 9548 10056
rect 10784 10047 10836 10056
rect 10784 10013 10793 10047
rect 10793 10013 10827 10047
rect 10827 10013 10836 10047
rect 10784 10004 10836 10013
rect 13912 10004 13964 10056
rect 14372 10004 14424 10056
rect 15200 10047 15252 10056
rect 15200 10013 15209 10047
rect 15209 10013 15243 10047
rect 15243 10013 15252 10047
rect 15200 10004 15252 10013
rect 15384 10047 15436 10056
rect 15384 10013 15393 10047
rect 15393 10013 15427 10047
rect 15427 10013 15436 10047
rect 15384 10004 15436 10013
rect 15568 10115 15620 10124
rect 15568 10081 15577 10115
rect 15577 10081 15611 10115
rect 15611 10081 15620 10115
rect 15568 10072 15620 10081
rect 16120 10115 16172 10124
rect 16120 10081 16129 10115
rect 16129 10081 16163 10115
rect 16163 10081 16172 10115
rect 16120 10072 16172 10081
rect 16028 10047 16080 10056
rect 16028 10013 16037 10047
rect 16037 10013 16071 10047
rect 16071 10013 16080 10047
rect 16028 10004 16080 10013
rect 17684 10140 17736 10192
rect 19708 10140 19760 10192
rect 21088 10140 21140 10192
rect 22008 10140 22060 10192
rect 16488 10004 16540 10056
rect 8300 9936 8352 9988
rect 8760 9936 8812 9988
rect 5356 9868 5408 9920
rect 5816 9911 5868 9920
rect 5816 9877 5825 9911
rect 5825 9877 5859 9911
rect 5859 9877 5868 9911
rect 5816 9868 5868 9877
rect 7472 9868 7524 9920
rect 8116 9868 8168 9920
rect 8208 9868 8260 9920
rect 14924 9936 14976 9988
rect 17040 10047 17092 10056
rect 17040 10013 17049 10047
rect 17049 10013 17083 10047
rect 17083 10013 17092 10047
rect 17040 10004 17092 10013
rect 17224 10004 17276 10056
rect 17316 10047 17368 10056
rect 17316 10013 17325 10047
rect 17325 10013 17359 10047
rect 17359 10013 17368 10047
rect 17316 10004 17368 10013
rect 10048 9911 10100 9920
rect 10048 9877 10057 9911
rect 10057 9877 10091 9911
rect 10091 9877 10100 9911
rect 10048 9868 10100 9877
rect 14096 9911 14148 9920
rect 14096 9877 14105 9911
rect 14105 9877 14139 9911
rect 14139 9877 14148 9911
rect 14096 9868 14148 9877
rect 14464 9911 14516 9920
rect 14464 9877 14473 9911
rect 14473 9877 14507 9911
rect 14507 9877 14516 9911
rect 14464 9868 14516 9877
rect 16212 9868 16264 9920
rect 16396 9911 16448 9920
rect 16396 9877 16405 9911
rect 16405 9877 16439 9911
rect 16439 9877 16448 9911
rect 16396 9868 16448 9877
rect 19984 10115 20036 10124
rect 19984 10081 19993 10115
rect 19993 10081 20027 10115
rect 20027 10081 20036 10115
rect 19984 10072 20036 10081
rect 20628 10072 20680 10124
rect 19708 10047 19760 10056
rect 19708 10013 19717 10047
rect 19717 10013 19751 10047
rect 19751 10013 19760 10047
rect 19708 10004 19760 10013
rect 20168 10047 20220 10056
rect 20168 10013 20177 10047
rect 20177 10013 20211 10047
rect 20211 10013 20220 10047
rect 20168 10004 20220 10013
rect 20352 10047 20404 10056
rect 20352 10013 20361 10047
rect 20361 10013 20395 10047
rect 20395 10013 20404 10047
rect 20352 10004 20404 10013
rect 20444 10004 20496 10056
rect 21088 10047 21140 10056
rect 21088 10013 21097 10047
rect 21097 10013 21131 10047
rect 21131 10013 21140 10047
rect 21088 10004 21140 10013
rect 21272 10047 21324 10056
rect 21272 10013 21281 10047
rect 21281 10013 21315 10047
rect 21315 10013 21324 10047
rect 21272 10004 21324 10013
rect 21456 10115 21508 10124
rect 21456 10081 21465 10115
rect 21465 10081 21499 10115
rect 21499 10081 21508 10115
rect 21456 10072 21508 10081
rect 21640 10047 21692 10056
rect 21640 10013 21649 10047
rect 21649 10013 21683 10047
rect 21683 10013 21692 10047
rect 21640 10004 21692 10013
rect 22560 10251 22612 10260
rect 22560 10217 22569 10251
rect 22569 10217 22603 10251
rect 22603 10217 22612 10251
rect 22560 10208 22612 10217
rect 25964 10251 26016 10260
rect 25964 10217 25973 10251
rect 25973 10217 26007 10251
rect 26007 10217 26016 10251
rect 25964 10208 26016 10217
rect 26332 10251 26384 10260
rect 26332 10217 26341 10251
rect 26341 10217 26375 10251
rect 26375 10217 26384 10251
rect 26332 10208 26384 10217
rect 26424 10251 26476 10260
rect 26424 10217 26433 10251
rect 26433 10217 26467 10251
rect 26467 10217 26476 10251
rect 26424 10208 26476 10217
rect 24400 10140 24452 10192
rect 25688 10140 25740 10192
rect 23572 10115 23624 10124
rect 23572 10081 23581 10115
rect 23581 10081 23615 10115
rect 23615 10081 23624 10115
rect 23572 10072 23624 10081
rect 21180 9936 21232 9988
rect 21364 9979 21416 9988
rect 21364 9945 21373 9979
rect 21373 9945 21407 9979
rect 21407 9945 21416 9979
rect 21364 9936 21416 9945
rect 17592 9868 17644 9920
rect 17684 9911 17736 9920
rect 17684 9877 17693 9911
rect 17693 9877 17727 9911
rect 17727 9877 17736 9911
rect 17684 9868 17736 9877
rect 22284 10047 22336 10056
rect 22284 10013 22293 10047
rect 22293 10013 22327 10047
rect 22327 10013 22336 10047
rect 22284 10004 22336 10013
rect 22376 10047 22428 10056
rect 22376 10013 22390 10047
rect 22390 10013 22424 10047
rect 22424 10013 22428 10047
rect 22376 10004 22428 10013
rect 23480 10047 23532 10056
rect 23480 10013 23489 10047
rect 23489 10013 23523 10047
rect 23523 10013 23532 10047
rect 23480 10004 23532 10013
rect 23940 10047 23992 10056
rect 23940 10013 23949 10047
rect 23949 10013 23983 10047
rect 23983 10013 23992 10047
rect 23940 10004 23992 10013
rect 22100 9868 22152 9920
rect 22928 9936 22980 9988
rect 25504 10047 25556 10056
rect 25504 10013 25513 10047
rect 25513 10013 25547 10047
rect 25547 10013 25556 10047
rect 25504 10004 25556 10013
rect 25688 10004 25740 10056
rect 26424 10072 26476 10124
rect 26516 10004 26568 10056
rect 24032 9911 24084 9920
rect 24032 9877 24041 9911
rect 24041 9877 24075 9911
rect 24075 9877 24084 9911
rect 24032 9868 24084 9877
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 4712 9664 4764 9716
rect 5356 9664 5408 9716
rect 8208 9664 8260 9716
rect 9312 9707 9364 9716
rect 9312 9673 9321 9707
rect 9321 9673 9355 9707
rect 9355 9673 9364 9707
rect 9312 9664 9364 9673
rect 17224 9664 17276 9716
rect 17684 9664 17736 9716
rect 23572 9664 23624 9716
rect 3884 9571 3936 9580
rect 3884 9537 3893 9571
rect 3893 9537 3927 9571
rect 3927 9537 3936 9571
rect 3884 9528 3936 9537
rect 6552 9596 6604 9648
rect 4620 9503 4672 9512
rect 4620 9469 4629 9503
rect 4629 9469 4663 9503
rect 4663 9469 4672 9503
rect 4620 9460 4672 9469
rect 4712 9503 4764 9512
rect 4712 9469 4721 9503
rect 4721 9469 4755 9503
rect 4755 9469 4764 9503
rect 4712 9460 4764 9469
rect 5356 9528 5408 9580
rect 5540 9528 5592 9580
rect 5632 9571 5684 9580
rect 5632 9537 5651 9571
rect 5651 9537 5684 9571
rect 5632 9528 5684 9537
rect 6644 9528 6696 9580
rect 7196 9571 7248 9580
rect 7196 9537 7205 9571
rect 7205 9537 7239 9571
rect 7239 9537 7248 9571
rect 7196 9528 7248 9537
rect 7472 9639 7524 9648
rect 7472 9605 7481 9639
rect 7481 9605 7515 9639
rect 7515 9605 7524 9639
rect 7472 9596 7524 9605
rect 8760 9639 8812 9648
rect 8760 9605 8769 9639
rect 8769 9605 8803 9639
rect 8803 9605 8812 9639
rect 8760 9596 8812 9605
rect 11888 9596 11940 9648
rect 4988 9503 5040 9512
rect 4988 9469 4997 9503
rect 4997 9469 5031 9503
rect 5031 9469 5040 9503
rect 4988 9460 5040 9469
rect 3424 9367 3476 9376
rect 3424 9333 3433 9367
rect 3433 9333 3467 9367
rect 3467 9333 3476 9367
rect 3424 9324 3476 9333
rect 3792 9324 3844 9376
rect 4712 9324 4764 9376
rect 5816 9392 5868 9444
rect 7840 9460 7892 9512
rect 10324 9528 10376 9580
rect 11704 9571 11756 9580
rect 11704 9537 11713 9571
rect 11713 9537 11747 9571
rect 11747 9537 11756 9571
rect 11704 9528 11756 9537
rect 12808 9571 12860 9580
rect 12808 9537 12817 9571
rect 12817 9537 12851 9571
rect 12851 9537 12860 9571
rect 12808 9528 12860 9537
rect 13912 9528 13964 9580
rect 15200 9528 15252 9580
rect 15476 9571 15528 9580
rect 15476 9537 15485 9571
rect 15485 9537 15519 9571
rect 15519 9537 15528 9571
rect 15476 9528 15528 9537
rect 16488 9528 16540 9580
rect 17408 9528 17460 9580
rect 19524 9571 19576 9580
rect 19524 9537 19533 9571
rect 19533 9537 19567 9571
rect 19567 9537 19576 9571
rect 19524 9528 19576 9537
rect 19708 9596 19760 9648
rect 19800 9571 19852 9580
rect 19800 9537 19809 9571
rect 19809 9537 19843 9571
rect 19843 9537 19852 9571
rect 19800 9528 19852 9537
rect 24584 9596 24636 9648
rect 23756 9571 23808 9580
rect 23756 9537 23765 9571
rect 23765 9537 23799 9571
rect 23799 9537 23808 9571
rect 23756 9528 23808 9537
rect 23848 9528 23900 9580
rect 24032 9571 24084 9580
rect 24032 9537 24041 9571
rect 24041 9537 24075 9571
rect 24075 9537 24084 9571
rect 24032 9528 24084 9537
rect 8576 9503 8628 9512
rect 8576 9469 8585 9503
rect 8585 9469 8619 9503
rect 8619 9469 8628 9503
rect 8576 9460 8628 9469
rect 9404 9503 9456 9512
rect 9404 9469 9413 9503
rect 9413 9469 9447 9503
rect 9447 9469 9456 9503
rect 9404 9460 9456 9469
rect 11796 9503 11848 9512
rect 11796 9469 11805 9503
rect 11805 9469 11839 9503
rect 11839 9469 11848 9503
rect 11796 9460 11848 9469
rect 14464 9503 14516 9512
rect 14464 9469 14473 9503
rect 14473 9469 14507 9503
rect 14507 9469 14516 9503
rect 14464 9460 14516 9469
rect 5540 9367 5592 9376
rect 5540 9333 5549 9367
rect 5549 9333 5583 9367
rect 5583 9333 5592 9367
rect 5540 9324 5592 9333
rect 6552 9367 6604 9376
rect 6552 9333 6561 9367
rect 6561 9333 6595 9367
rect 6595 9333 6604 9367
rect 6552 9324 6604 9333
rect 7196 9324 7248 9376
rect 12072 9435 12124 9444
rect 12072 9401 12081 9435
rect 12081 9401 12115 9435
rect 12115 9401 12124 9435
rect 12072 9392 12124 9401
rect 13636 9392 13688 9444
rect 14188 9324 14240 9376
rect 16028 9460 16080 9512
rect 19892 9460 19944 9512
rect 25780 9460 25832 9512
rect 17316 9392 17368 9444
rect 16856 9367 16908 9376
rect 16856 9333 16865 9367
rect 16865 9333 16899 9367
rect 16899 9333 16908 9367
rect 16856 9324 16908 9333
rect 19524 9324 19576 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 8208 9120 8260 9172
rect 12808 9163 12860 9172
rect 12808 9129 12817 9163
rect 12817 9129 12851 9163
rect 12851 9129 12860 9163
rect 12808 9120 12860 9129
rect 16396 9120 16448 9172
rect 20168 9120 20220 9172
rect 21456 9120 21508 9172
rect 21640 9120 21692 9172
rect 4988 9052 5040 9104
rect 5264 9052 5316 9104
rect 3424 8984 3476 9036
rect 3792 8959 3844 8968
rect 3792 8925 3801 8959
rect 3801 8925 3835 8959
rect 3835 8925 3844 8959
rect 3792 8916 3844 8925
rect 5448 8916 5500 8968
rect 5540 8916 5592 8968
rect 11428 9052 11480 9104
rect 6552 9027 6604 9036
rect 6552 8993 6561 9027
rect 6561 8993 6595 9027
rect 6595 8993 6604 9027
rect 6552 8984 6604 8993
rect 9772 8984 9824 9036
rect 6736 8959 6788 8968
rect 6736 8925 6745 8959
rect 6745 8925 6779 8959
rect 6779 8925 6788 8959
rect 6736 8916 6788 8925
rect 7840 8916 7892 8968
rect 8116 8959 8168 8968
rect 8116 8925 8125 8959
rect 8125 8925 8159 8959
rect 8159 8925 8168 8959
rect 8116 8916 8168 8925
rect 10140 8984 10192 9036
rect 11244 8984 11296 9036
rect 13636 9027 13688 9036
rect 13636 8993 13645 9027
rect 13645 8993 13679 9027
rect 13679 8993 13688 9027
rect 13636 8984 13688 8993
rect 13820 8984 13872 9036
rect 15108 8984 15160 9036
rect 15568 8984 15620 9036
rect 16856 9027 16908 9036
rect 16856 8993 16865 9027
rect 16865 8993 16899 9027
rect 16899 8993 16908 9027
rect 16856 8984 16908 8993
rect 22100 9052 22152 9104
rect 11060 8959 11112 8968
rect 11060 8925 11069 8959
rect 11069 8925 11103 8959
rect 11103 8925 11112 8959
rect 11060 8916 11112 8925
rect 11152 8916 11204 8968
rect 11612 8916 11664 8968
rect 12348 8959 12400 8968
rect 12348 8925 12357 8959
rect 12357 8925 12391 8959
rect 12391 8925 12400 8959
rect 12348 8916 12400 8925
rect 12624 8959 12676 8968
rect 12624 8925 12633 8959
rect 12633 8925 12667 8959
rect 12667 8925 12676 8959
rect 12624 8916 12676 8925
rect 14096 8916 14148 8968
rect 14280 8959 14332 8968
rect 14280 8925 14289 8959
rect 14289 8925 14323 8959
rect 14323 8925 14332 8959
rect 14280 8916 14332 8925
rect 14464 8959 14516 8968
rect 14464 8925 14473 8959
rect 14473 8925 14507 8959
rect 14507 8925 14516 8959
rect 14464 8916 14516 8925
rect 11244 8848 11296 8900
rect 17040 8916 17092 8968
rect 17684 8959 17736 8968
rect 17684 8925 17693 8959
rect 17693 8925 17727 8959
rect 17727 8925 17736 8959
rect 17684 8916 17736 8925
rect 17868 8959 17920 8968
rect 17868 8925 17877 8959
rect 17877 8925 17911 8959
rect 17911 8925 17920 8959
rect 17868 8916 17920 8925
rect 16212 8891 16264 8900
rect 16212 8857 16237 8891
rect 16237 8857 16264 8891
rect 18144 8959 18196 8968
rect 18144 8925 18153 8959
rect 18153 8925 18187 8959
rect 18187 8925 18196 8959
rect 18144 8916 18196 8925
rect 24584 9052 24636 9104
rect 25596 9052 25648 9104
rect 20260 8959 20312 8968
rect 20260 8925 20269 8959
rect 20269 8925 20303 8959
rect 20303 8925 20312 8959
rect 20260 8916 20312 8925
rect 21364 8916 21416 8968
rect 21640 8916 21692 8968
rect 22284 8984 22336 9036
rect 21916 8916 21968 8968
rect 22008 8959 22060 8968
rect 22008 8925 22017 8959
rect 22017 8925 22051 8959
rect 22051 8925 22060 8959
rect 22008 8916 22060 8925
rect 16212 8848 16264 8857
rect 4804 8780 4856 8832
rect 5908 8780 5960 8832
rect 7472 8823 7524 8832
rect 7472 8789 7481 8823
rect 7481 8789 7515 8823
rect 7515 8789 7524 8823
rect 7472 8780 7524 8789
rect 7748 8823 7800 8832
rect 7748 8789 7757 8823
rect 7757 8789 7791 8823
rect 7791 8789 7800 8823
rect 7748 8780 7800 8789
rect 11060 8780 11112 8832
rect 19524 8891 19576 8900
rect 19524 8857 19533 8891
rect 19533 8857 19567 8891
rect 19567 8857 19576 8891
rect 19524 8848 19576 8857
rect 22192 8916 22244 8968
rect 22376 8959 22428 8968
rect 22376 8925 22385 8959
rect 22385 8925 22419 8959
rect 22419 8925 22428 8959
rect 22376 8916 22428 8925
rect 23848 8984 23900 9036
rect 23296 8916 23348 8968
rect 24216 8959 24268 8968
rect 24216 8925 24225 8959
rect 24225 8925 24259 8959
rect 24259 8925 24268 8959
rect 24216 8916 24268 8925
rect 24400 8959 24452 8968
rect 24400 8925 24409 8959
rect 24409 8925 24443 8959
rect 24443 8925 24452 8959
rect 24400 8916 24452 8925
rect 24676 8959 24728 8968
rect 24676 8925 24685 8959
rect 24685 8925 24719 8959
rect 24719 8925 24728 8959
rect 24676 8916 24728 8925
rect 25780 8916 25832 8968
rect 17408 8780 17460 8832
rect 17868 8780 17920 8832
rect 18052 8823 18104 8832
rect 18052 8789 18061 8823
rect 18061 8789 18095 8823
rect 18095 8789 18104 8823
rect 18052 8780 18104 8789
rect 19708 8823 19760 8832
rect 19708 8789 19733 8823
rect 19733 8789 19760 8823
rect 19708 8780 19760 8789
rect 20352 8780 20404 8832
rect 20444 8780 20496 8832
rect 22192 8780 22244 8832
rect 22652 8823 22704 8832
rect 22652 8789 22661 8823
rect 22661 8789 22695 8823
rect 22695 8789 22704 8823
rect 22652 8780 22704 8789
rect 22744 8823 22796 8832
rect 22744 8789 22753 8823
rect 22753 8789 22787 8823
rect 22787 8789 22796 8823
rect 22744 8780 22796 8789
rect 24124 8823 24176 8832
rect 24124 8789 24133 8823
rect 24133 8789 24167 8823
rect 24167 8789 24176 8823
rect 24124 8780 24176 8789
rect 24492 8780 24544 8832
rect 25136 8780 25188 8832
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 4896 8576 4948 8628
rect 10140 8619 10192 8628
rect 10140 8585 10149 8619
rect 10149 8585 10183 8619
rect 10183 8585 10192 8619
rect 10140 8576 10192 8585
rect 6828 8508 6880 8560
rect 3516 8483 3568 8492
rect 3516 8449 3525 8483
rect 3525 8449 3559 8483
rect 3559 8449 3568 8483
rect 3516 8440 3568 8449
rect 4620 8483 4672 8492
rect 4620 8449 4629 8483
rect 4629 8449 4663 8483
rect 4663 8449 4672 8483
rect 4620 8440 4672 8449
rect 4712 8440 4764 8492
rect 5080 8440 5132 8492
rect 3424 8415 3476 8424
rect 3424 8381 3433 8415
rect 3433 8381 3467 8415
rect 3467 8381 3476 8415
rect 3424 8372 3476 8381
rect 4988 8372 5040 8424
rect 6736 8372 6788 8424
rect 4712 8304 4764 8356
rect 5264 8236 5316 8288
rect 10140 8440 10192 8492
rect 11152 8440 11204 8492
rect 11244 8483 11296 8492
rect 11244 8449 11253 8483
rect 11253 8449 11287 8483
rect 11287 8449 11296 8483
rect 11244 8440 11296 8449
rect 12624 8483 12676 8492
rect 12624 8449 12633 8483
rect 12633 8449 12667 8483
rect 12667 8449 12676 8483
rect 12624 8440 12676 8449
rect 9772 8372 9824 8424
rect 9864 8372 9916 8424
rect 14188 8483 14240 8492
rect 14188 8449 14197 8483
rect 14197 8449 14231 8483
rect 14231 8449 14240 8483
rect 14188 8440 14240 8449
rect 15476 8576 15528 8628
rect 20260 8619 20312 8628
rect 20260 8585 20269 8619
rect 20269 8585 20303 8619
rect 20303 8585 20312 8619
rect 20260 8576 20312 8585
rect 21640 8576 21692 8628
rect 16028 8508 16080 8560
rect 15016 8440 15068 8492
rect 16396 8440 16448 8492
rect 17040 8483 17092 8492
rect 17040 8449 17049 8483
rect 17049 8449 17083 8483
rect 17083 8449 17092 8483
rect 17040 8440 17092 8449
rect 18144 8508 18196 8560
rect 17592 8440 17644 8492
rect 16212 8372 16264 8424
rect 17132 8415 17184 8424
rect 17132 8381 17141 8415
rect 17141 8381 17175 8415
rect 17175 8381 17184 8415
rect 17132 8372 17184 8381
rect 19524 8440 19576 8492
rect 17868 8372 17920 8424
rect 20352 8440 20404 8492
rect 20536 8440 20588 8492
rect 22008 8483 22060 8492
rect 22008 8449 22017 8483
rect 22017 8449 22051 8483
rect 22051 8449 22060 8483
rect 22008 8440 22060 8449
rect 22376 8576 22428 8628
rect 24216 8508 24268 8560
rect 24676 8508 24728 8560
rect 22192 8440 22244 8492
rect 22744 8483 22796 8492
rect 22744 8449 22753 8483
rect 22753 8449 22787 8483
rect 22787 8449 22796 8483
rect 22744 8440 22796 8449
rect 23296 8483 23348 8492
rect 23296 8449 23305 8483
rect 23305 8449 23339 8483
rect 23339 8449 23348 8483
rect 23296 8440 23348 8449
rect 24400 8440 24452 8492
rect 9220 8304 9272 8356
rect 16304 8304 16356 8356
rect 17500 8304 17552 8356
rect 20720 8304 20772 8356
rect 25136 8415 25188 8424
rect 25136 8381 25145 8415
rect 25145 8381 25179 8415
rect 25179 8381 25188 8415
rect 25136 8372 25188 8381
rect 8300 8236 8352 8288
rect 9772 8279 9824 8288
rect 9772 8245 9781 8279
rect 9781 8245 9815 8279
rect 9815 8245 9824 8279
rect 9772 8236 9824 8245
rect 10048 8236 10100 8288
rect 11244 8236 11296 8288
rect 14004 8279 14056 8288
rect 14004 8245 14013 8279
rect 14013 8245 14047 8279
rect 14047 8245 14056 8279
rect 14004 8236 14056 8245
rect 19800 8236 19852 8288
rect 21916 8304 21968 8356
rect 23388 8304 23440 8356
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 4712 7964 4764 8016
rect 4620 7896 4672 7948
rect 5448 8007 5500 8016
rect 5448 7973 5457 8007
rect 5457 7973 5491 8007
rect 5491 7973 5500 8007
rect 5448 7964 5500 7973
rect 7840 8032 7892 8084
rect 8944 8032 8996 8084
rect 11152 8032 11204 8084
rect 12900 8032 12952 8084
rect 13176 8032 13228 8084
rect 14188 8032 14240 8084
rect 17132 8032 17184 8084
rect 20352 8032 20404 8084
rect 21272 8032 21324 8084
rect 24400 8032 24452 8084
rect 5264 7871 5316 7880
rect 5264 7837 5273 7871
rect 5273 7837 5307 7871
rect 5307 7837 5316 7871
rect 5264 7828 5316 7837
rect 12440 7964 12492 8016
rect 14280 7964 14332 8016
rect 7656 7871 7708 7880
rect 7656 7837 7665 7871
rect 7665 7837 7699 7871
rect 7699 7837 7708 7871
rect 7656 7828 7708 7837
rect 7840 7871 7892 7880
rect 7840 7837 7849 7871
rect 7849 7837 7883 7871
rect 7883 7837 7892 7871
rect 7840 7828 7892 7837
rect 8116 7828 8168 7880
rect 8484 7871 8536 7880
rect 8484 7837 8493 7871
rect 8493 7837 8527 7871
rect 8527 7837 8536 7871
rect 8484 7828 8536 7837
rect 8576 7871 8628 7880
rect 8576 7837 8585 7871
rect 8585 7837 8619 7871
rect 8619 7837 8628 7871
rect 8576 7828 8628 7837
rect 8944 7871 8996 7880
rect 8944 7837 8953 7871
rect 8953 7837 8987 7871
rect 8987 7837 8996 7871
rect 8944 7828 8996 7837
rect 9220 7896 9272 7948
rect 11428 7939 11480 7948
rect 11428 7905 11437 7939
rect 11437 7905 11471 7939
rect 11471 7905 11480 7939
rect 11428 7896 11480 7905
rect 9772 7871 9824 7880
rect 9772 7837 9781 7871
rect 9781 7837 9815 7871
rect 9815 7837 9824 7871
rect 9772 7828 9824 7837
rect 9864 7871 9916 7880
rect 9864 7837 9873 7871
rect 9873 7837 9907 7871
rect 9907 7837 9916 7871
rect 9864 7828 9916 7837
rect 4896 7760 4948 7812
rect 5356 7760 5408 7812
rect 5632 7803 5684 7812
rect 5632 7769 5641 7803
rect 5641 7769 5675 7803
rect 5675 7769 5684 7803
rect 5632 7760 5684 7769
rect 4436 7692 4488 7744
rect 4988 7692 5040 7744
rect 5080 7692 5132 7744
rect 5264 7692 5316 7744
rect 6736 7760 6788 7812
rect 9588 7760 9640 7812
rect 10048 7828 10100 7880
rect 11336 7871 11388 7880
rect 11336 7837 11345 7871
rect 11345 7837 11379 7871
rect 11379 7837 11388 7871
rect 11336 7828 11388 7837
rect 12532 7803 12584 7812
rect 12532 7769 12541 7803
rect 12541 7769 12575 7803
rect 12575 7769 12584 7803
rect 12532 7760 12584 7769
rect 13452 7896 13504 7948
rect 14004 7896 14056 7948
rect 20444 7896 20496 7948
rect 24216 7896 24268 7948
rect 12900 7828 12952 7880
rect 6552 7692 6604 7744
rect 8668 7692 8720 7744
rect 9496 7735 9548 7744
rect 9496 7701 9505 7735
rect 9505 7701 9539 7735
rect 9539 7701 9548 7735
rect 9496 7692 9548 7701
rect 12164 7692 12216 7744
rect 13268 7760 13320 7812
rect 13636 7828 13688 7880
rect 13728 7760 13780 7812
rect 14832 7803 14884 7812
rect 14832 7769 14841 7803
rect 14841 7769 14875 7803
rect 14875 7769 14884 7803
rect 14832 7760 14884 7769
rect 14924 7692 14976 7744
rect 17592 7871 17644 7880
rect 17592 7837 17601 7871
rect 17601 7837 17635 7871
rect 17635 7837 17644 7871
rect 17592 7828 17644 7837
rect 18052 7828 18104 7880
rect 19616 7871 19668 7880
rect 19616 7837 19625 7871
rect 19625 7837 19659 7871
rect 19659 7837 19668 7871
rect 19616 7828 19668 7837
rect 19800 7871 19852 7880
rect 19800 7837 19809 7871
rect 19809 7837 19843 7871
rect 19843 7837 19852 7871
rect 19800 7828 19852 7837
rect 21272 7828 21324 7880
rect 22284 7871 22336 7880
rect 22284 7837 22293 7871
rect 22293 7837 22327 7871
rect 22327 7837 22336 7871
rect 22284 7828 22336 7837
rect 22376 7828 22428 7880
rect 23480 7828 23532 7880
rect 17316 7760 17368 7812
rect 17500 7760 17552 7812
rect 21088 7760 21140 7812
rect 24308 7760 24360 7812
rect 18052 7735 18104 7744
rect 18052 7701 18061 7735
rect 18061 7701 18095 7735
rect 18095 7701 18104 7735
rect 18052 7692 18104 7701
rect 19984 7735 20036 7744
rect 19984 7701 19993 7735
rect 19993 7701 20027 7735
rect 20027 7701 20036 7735
rect 19984 7692 20036 7701
rect 22928 7692 22980 7744
rect 23848 7735 23900 7744
rect 23848 7701 23857 7735
rect 23857 7701 23891 7735
rect 23891 7701 23900 7735
rect 23848 7692 23900 7701
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 4620 7488 4672 7540
rect 5264 7488 5316 7540
rect 4160 7420 4212 7472
rect 6644 7488 6696 7540
rect 11060 7531 11112 7540
rect 4436 7395 4488 7404
rect 4436 7361 4445 7395
rect 4445 7361 4479 7395
rect 4479 7361 4488 7395
rect 4436 7352 4488 7361
rect 4620 7395 4672 7404
rect 4620 7361 4629 7395
rect 4629 7361 4663 7395
rect 4663 7361 4672 7395
rect 4620 7352 4672 7361
rect 5724 7352 5776 7404
rect 4712 7216 4764 7268
rect 5816 7284 5868 7336
rect 6552 7395 6604 7404
rect 6552 7361 6561 7395
rect 6561 7361 6595 7395
rect 6595 7361 6604 7395
rect 6552 7352 6604 7361
rect 5356 7216 5408 7268
rect 6276 7216 6328 7268
rect 6552 7216 6604 7268
rect 6736 7352 6788 7404
rect 7472 7352 7524 7404
rect 8392 7420 8444 7472
rect 11060 7497 11069 7531
rect 11069 7497 11103 7531
rect 11103 7497 11112 7531
rect 11060 7488 11112 7497
rect 15016 7488 15068 7540
rect 17592 7488 17644 7540
rect 19616 7488 19668 7540
rect 21180 7531 21232 7540
rect 21180 7497 21189 7531
rect 21189 7497 21223 7531
rect 21223 7497 21232 7531
rect 21180 7488 21232 7497
rect 22376 7488 22428 7540
rect 23480 7488 23532 7540
rect 24952 7531 25004 7540
rect 24952 7497 24961 7531
rect 24961 7497 24995 7531
rect 24995 7497 25004 7531
rect 24952 7488 25004 7497
rect 25780 7488 25832 7540
rect 7656 7327 7708 7336
rect 7656 7293 7665 7327
rect 7665 7293 7699 7327
rect 7699 7293 7708 7327
rect 7656 7284 7708 7293
rect 8300 7395 8352 7404
rect 8300 7361 8309 7395
rect 8309 7361 8343 7395
rect 8343 7361 8352 7395
rect 8300 7352 8352 7361
rect 8116 7284 8168 7336
rect 9496 7420 9548 7472
rect 9864 7420 9916 7472
rect 11244 7463 11296 7472
rect 8668 7395 8720 7404
rect 8668 7361 8677 7395
rect 8677 7361 8711 7395
rect 8711 7361 8720 7395
rect 8668 7352 8720 7361
rect 10048 7352 10100 7404
rect 11244 7429 11253 7463
rect 11253 7429 11287 7463
rect 11287 7429 11296 7463
rect 11244 7420 11296 7429
rect 12992 7420 13044 7472
rect 14832 7420 14884 7472
rect 10968 7395 11020 7404
rect 10968 7361 10977 7395
rect 10977 7361 11011 7395
rect 11011 7361 11020 7395
rect 10968 7352 11020 7361
rect 12072 7352 12124 7404
rect 13176 7395 13228 7404
rect 13176 7361 13185 7395
rect 13185 7361 13219 7395
rect 13219 7361 13228 7395
rect 13176 7352 13228 7361
rect 13268 7395 13320 7404
rect 13268 7361 13277 7395
rect 13277 7361 13311 7395
rect 13311 7361 13320 7395
rect 13268 7352 13320 7361
rect 10968 7216 11020 7268
rect 12900 7284 12952 7336
rect 13544 7352 13596 7404
rect 13636 7352 13688 7404
rect 13452 7327 13504 7336
rect 13452 7293 13461 7327
rect 13461 7293 13495 7327
rect 13495 7293 13504 7327
rect 13452 7284 13504 7293
rect 13728 7284 13780 7336
rect 14924 7284 14976 7336
rect 12716 7216 12768 7268
rect 13268 7216 13320 7268
rect 17224 7395 17276 7404
rect 17224 7361 17233 7395
rect 17233 7361 17267 7395
rect 17267 7361 17276 7395
rect 17224 7352 17276 7361
rect 17316 7395 17368 7404
rect 17316 7361 17325 7395
rect 17325 7361 17359 7395
rect 17359 7361 17368 7395
rect 17316 7352 17368 7361
rect 16120 7284 16172 7336
rect 17868 7352 17920 7404
rect 19800 7395 19852 7404
rect 19800 7361 19809 7395
rect 19809 7361 19843 7395
rect 19843 7361 19852 7395
rect 19800 7352 19852 7361
rect 19984 7395 20036 7404
rect 19984 7361 19993 7395
rect 19993 7361 20027 7395
rect 20027 7361 20036 7395
rect 19984 7352 20036 7361
rect 21088 7395 21140 7404
rect 21088 7361 21127 7395
rect 21127 7361 21140 7395
rect 21088 7352 21140 7361
rect 22652 7420 22704 7472
rect 22928 7420 22980 7472
rect 25228 7420 25280 7472
rect 18052 7327 18104 7336
rect 18052 7293 18061 7327
rect 18061 7293 18095 7327
rect 18095 7293 18104 7327
rect 18052 7284 18104 7293
rect 21640 7327 21692 7336
rect 21640 7293 21649 7327
rect 21649 7293 21683 7327
rect 21683 7293 21692 7327
rect 21640 7284 21692 7293
rect 8852 7191 8904 7200
rect 8852 7157 8861 7191
rect 8861 7157 8895 7191
rect 8895 7157 8904 7191
rect 8852 7148 8904 7157
rect 10692 7148 10744 7200
rect 10876 7191 10928 7200
rect 10876 7157 10885 7191
rect 10885 7157 10919 7191
rect 10919 7157 10928 7191
rect 10876 7148 10928 7157
rect 13176 7148 13228 7200
rect 13728 7148 13780 7200
rect 17040 7191 17092 7200
rect 17040 7157 17049 7191
rect 17049 7157 17083 7191
rect 17083 7157 17092 7191
rect 17040 7148 17092 7157
rect 22100 7216 22152 7268
rect 22284 7216 22336 7268
rect 23848 7352 23900 7404
rect 24124 7395 24176 7404
rect 24124 7361 24133 7395
rect 24133 7361 24167 7395
rect 24167 7361 24176 7395
rect 24124 7352 24176 7361
rect 24308 7395 24360 7404
rect 24308 7361 24317 7395
rect 24317 7361 24351 7395
rect 24351 7361 24360 7395
rect 24308 7352 24360 7361
rect 25136 7352 25188 7404
rect 25596 7395 25648 7404
rect 25596 7361 25605 7395
rect 25605 7361 25639 7395
rect 25639 7361 25648 7395
rect 25596 7352 25648 7361
rect 23756 7284 23808 7336
rect 24492 7284 24544 7336
rect 25872 7259 25924 7268
rect 25872 7225 25881 7259
rect 25881 7225 25915 7259
rect 25915 7225 25924 7259
rect 25872 7216 25924 7225
rect 23388 7191 23440 7200
rect 23388 7157 23397 7191
rect 23397 7157 23431 7191
rect 23431 7157 23440 7191
rect 23388 7148 23440 7157
rect 25228 7148 25280 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 21180 6944 21232 6996
rect 21548 6987 21600 6996
rect 21548 6953 21557 6987
rect 21557 6953 21591 6987
rect 21591 6953 21600 6987
rect 21548 6944 21600 6953
rect 23756 6987 23808 6996
rect 23756 6953 23765 6987
rect 23765 6953 23799 6987
rect 23799 6953 23808 6987
rect 23756 6944 23808 6953
rect 25044 6944 25096 6996
rect 25596 6944 25648 6996
rect 6276 6876 6328 6928
rect 8300 6876 8352 6928
rect 10416 6876 10468 6928
rect 11060 6876 11112 6928
rect 12164 6876 12216 6928
rect 13268 6876 13320 6928
rect 6368 6740 6420 6792
rect 8852 6740 8904 6792
rect 7656 6672 7708 6724
rect 10416 6783 10468 6792
rect 10416 6749 10425 6783
rect 10425 6749 10459 6783
rect 10459 6749 10468 6783
rect 10416 6740 10468 6749
rect 9772 6672 9824 6724
rect 10692 6783 10744 6792
rect 10692 6749 10701 6783
rect 10701 6749 10735 6783
rect 10735 6749 10744 6783
rect 10692 6740 10744 6749
rect 10876 6740 10928 6792
rect 12348 6740 12400 6792
rect 15936 6783 15988 6792
rect 15936 6749 15945 6783
rect 15945 6749 15979 6783
rect 15979 6749 15988 6783
rect 15936 6740 15988 6749
rect 16120 6783 16172 6792
rect 16120 6749 16129 6783
rect 16129 6749 16163 6783
rect 16163 6749 16172 6783
rect 16120 6740 16172 6749
rect 16304 6783 16356 6792
rect 16304 6749 16313 6783
rect 16313 6749 16347 6783
rect 16347 6749 16356 6783
rect 16304 6740 16356 6749
rect 17040 6783 17092 6792
rect 17040 6749 17049 6783
rect 17049 6749 17083 6783
rect 17083 6749 17092 6783
rect 17040 6740 17092 6749
rect 16856 6672 16908 6724
rect 17408 6783 17460 6792
rect 17408 6749 17417 6783
rect 17417 6749 17451 6783
rect 17451 6749 17460 6783
rect 17408 6740 17460 6749
rect 18604 6740 18656 6792
rect 19616 6740 19668 6792
rect 19892 6783 19944 6792
rect 19892 6749 19901 6783
rect 19901 6749 19935 6783
rect 19935 6749 19944 6783
rect 19892 6740 19944 6749
rect 21640 6876 21692 6928
rect 21364 6851 21416 6860
rect 21364 6817 21373 6851
rect 21373 6817 21407 6851
rect 21407 6817 21416 6851
rect 21364 6808 21416 6817
rect 22376 6919 22428 6928
rect 22376 6885 22385 6919
rect 22385 6885 22419 6919
rect 22419 6885 22428 6919
rect 22376 6876 22428 6885
rect 24952 6808 25004 6860
rect 25780 6876 25832 6928
rect 20260 6740 20312 6792
rect 18696 6672 18748 6724
rect 6184 6647 6236 6656
rect 6184 6613 6193 6647
rect 6193 6613 6227 6647
rect 6227 6613 6236 6647
rect 6184 6604 6236 6613
rect 6736 6604 6788 6656
rect 10232 6604 10284 6656
rect 10416 6604 10468 6656
rect 11060 6604 11112 6656
rect 16120 6604 16172 6656
rect 19800 6604 19852 6656
rect 20260 6604 20312 6656
rect 20352 6647 20404 6656
rect 20352 6613 20361 6647
rect 20361 6613 20395 6647
rect 20395 6613 20404 6647
rect 20352 6604 20404 6613
rect 20720 6715 20772 6724
rect 20720 6681 20729 6715
rect 20729 6681 20763 6715
rect 20763 6681 20772 6715
rect 20720 6672 20772 6681
rect 20904 6715 20956 6724
rect 20904 6681 20913 6715
rect 20913 6681 20947 6715
rect 20947 6681 20956 6715
rect 20904 6672 20956 6681
rect 20996 6672 21048 6724
rect 23388 6740 23440 6792
rect 23572 6783 23624 6792
rect 23572 6749 23581 6783
rect 23581 6749 23615 6783
rect 23615 6749 23624 6783
rect 23572 6740 23624 6749
rect 23756 6783 23808 6792
rect 23756 6749 23765 6783
rect 23765 6749 23799 6783
rect 23799 6749 23808 6783
rect 23756 6740 23808 6749
rect 25044 6783 25096 6792
rect 25044 6749 25053 6783
rect 25053 6749 25087 6783
rect 25087 6749 25096 6783
rect 25044 6740 25096 6749
rect 25228 6740 25280 6792
rect 25596 6740 25648 6792
rect 25872 6783 25924 6792
rect 25872 6749 25881 6783
rect 25881 6749 25915 6783
rect 25915 6749 25924 6783
rect 25872 6740 25924 6749
rect 25780 6715 25832 6724
rect 25780 6681 25789 6715
rect 25789 6681 25823 6715
rect 25823 6681 25832 6715
rect 25780 6672 25832 6681
rect 23664 6604 23716 6656
rect 25136 6604 25188 6656
rect 26148 6604 26200 6656
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 5632 6443 5684 6452
rect 5632 6409 5641 6443
rect 5641 6409 5675 6443
rect 5675 6409 5684 6443
rect 5632 6400 5684 6409
rect 6736 6400 6788 6452
rect 7656 6400 7708 6452
rect 5264 6264 5316 6316
rect 6644 6375 6696 6384
rect 6644 6341 6653 6375
rect 6653 6341 6687 6375
rect 6687 6341 6696 6375
rect 6644 6332 6696 6341
rect 5540 6307 5592 6316
rect 5540 6273 5549 6307
rect 5549 6273 5583 6307
rect 5583 6273 5592 6307
rect 5540 6264 5592 6273
rect 5724 6264 5776 6316
rect 6184 6264 6236 6316
rect 6000 6196 6052 6248
rect 5724 6128 5776 6180
rect 6828 6264 6880 6316
rect 7564 6307 7616 6316
rect 7564 6273 7573 6307
rect 7573 6273 7607 6307
rect 7607 6273 7616 6307
rect 7564 6264 7616 6273
rect 7748 6307 7800 6316
rect 7748 6273 7757 6307
rect 7757 6273 7791 6307
rect 7791 6273 7800 6307
rect 7748 6264 7800 6273
rect 10048 6264 10100 6316
rect 12072 6332 12124 6384
rect 11980 6264 12032 6316
rect 12624 6264 12676 6316
rect 12992 6400 13044 6452
rect 13820 6400 13872 6452
rect 14832 6400 14884 6452
rect 10416 6239 10468 6248
rect 10416 6205 10425 6239
rect 10425 6205 10459 6239
rect 10459 6205 10468 6239
rect 10416 6196 10468 6205
rect 11888 6239 11940 6248
rect 11888 6205 11897 6239
rect 11897 6205 11931 6239
rect 11931 6205 11940 6239
rect 11888 6196 11940 6205
rect 9956 6128 10008 6180
rect 4804 6103 4856 6112
rect 4804 6069 4813 6103
rect 4813 6069 4847 6103
rect 4847 6069 4856 6103
rect 4804 6060 4856 6069
rect 11796 6103 11848 6112
rect 11796 6069 11805 6103
rect 11805 6069 11839 6103
rect 11839 6069 11848 6103
rect 11796 6060 11848 6069
rect 14372 6332 14424 6384
rect 15936 6400 15988 6452
rect 16304 6400 16356 6452
rect 20996 6443 21048 6452
rect 20996 6409 21005 6443
rect 21005 6409 21039 6443
rect 21039 6409 21048 6443
rect 20996 6400 21048 6409
rect 23572 6400 23624 6452
rect 18696 6375 18748 6384
rect 18696 6341 18705 6375
rect 18705 6341 18739 6375
rect 18739 6341 18748 6375
rect 18696 6332 18748 6341
rect 12992 6307 13044 6316
rect 12992 6273 13001 6307
rect 13001 6273 13035 6307
rect 13035 6273 13044 6307
rect 12992 6264 13044 6273
rect 13176 6264 13228 6316
rect 13268 6307 13320 6316
rect 13268 6273 13277 6307
rect 13277 6273 13311 6307
rect 13311 6273 13320 6307
rect 13268 6264 13320 6273
rect 14096 6264 14148 6316
rect 15200 6307 15252 6316
rect 15200 6273 15209 6307
rect 15209 6273 15243 6307
rect 15243 6273 15252 6307
rect 15200 6264 15252 6273
rect 15844 6307 15896 6316
rect 15844 6273 15853 6307
rect 15853 6273 15887 6307
rect 15887 6273 15896 6307
rect 15844 6264 15896 6273
rect 16120 6307 16172 6316
rect 16120 6273 16129 6307
rect 16129 6273 16163 6307
rect 16163 6273 16172 6307
rect 16120 6264 16172 6273
rect 18420 6264 18472 6316
rect 18604 6307 18656 6316
rect 18604 6273 18613 6307
rect 18613 6273 18647 6307
rect 18647 6273 18656 6307
rect 18604 6264 18656 6273
rect 20904 6332 20956 6384
rect 13084 6128 13136 6180
rect 12808 6060 12860 6112
rect 12900 6103 12952 6112
rect 12900 6069 12909 6103
rect 12909 6069 12943 6103
rect 12943 6069 12952 6103
rect 12900 6060 12952 6069
rect 13728 6103 13780 6112
rect 13728 6069 13737 6103
rect 13737 6069 13771 6103
rect 13771 6069 13780 6103
rect 14372 6239 14424 6248
rect 14372 6205 14381 6239
rect 14381 6205 14415 6239
rect 14415 6205 14424 6239
rect 14372 6196 14424 6205
rect 14464 6128 14516 6180
rect 18328 6239 18380 6248
rect 18328 6205 18337 6239
rect 18337 6205 18371 6239
rect 18371 6205 18380 6239
rect 18328 6196 18380 6205
rect 13728 6060 13780 6069
rect 15568 6060 15620 6112
rect 20720 6264 20772 6316
rect 21548 6264 21600 6316
rect 21916 6264 21968 6316
rect 23204 6307 23256 6316
rect 23204 6273 23213 6307
rect 23213 6273 23247 6307
rect 23247 6273 23256 6307
rect 23204 6264 23256 6273
rect 23480 6307 23532 6316
rect 23480 6273 23489 6307
rect 23489 6273 23523 6307
rect 23523 6273 23532 6307
rect 23480 6264 23532 6273
rect 25780 6400 25832 6452
rect 25136 6196 25188 6248
rect 21364 6128 21416 6180
rect 21824 6128 21876 6180
rect 23480 6128 23532 6180
rect 25596 6128 25648 6180
rect 21088 6103 21140 6112
rect 21088 6069 21097 6103
rect 21097 6069 21131 6103
rect 21131 6069 21140 6103
rect 21088 6060 21140 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 11980 5856 12032 5908
rect 12624 5899 12676 5908
rect 12624 5865 12633 5899
rect 12633 5865 12667 5899
rect 12667 5865 12676 5899
rect 12624 5856 12676 5865
rect 12716 5899 12768 5908
rect 12716 5865 12725 5899
rect 12725 5865 12759 5899
rect 12759 5865 12768 5899
rect 12716 5856 12768 5865
rect 13084 5899 13136 5908
rect 13084 5865 13093 5899
rect 13093 5865 13127 5899
rect 13127 5865 13136 5899
rect 13084 5856 13136 5865
rect 14832 5899 14884 5908
rect 14832 5865 14841 5899
rect 14841 5865 14875 5899
rect 14875 5865 14884 5899
rect 14832 5856 14884 5865
rect 16304 5856 16356 5908
rect 7656 5720 7708 5772
rect 7932 5720 7984 5772
rect 9772 5720 9824 5772
rect 5908 5695 5960 5704
rect 5908 5661 5917 5695
rect 5917 5661 5951 5695
rect 5951 5661 5960 5695
rect 5908 5652 5960 5661
rect 6092 5695 6144 5704
rect 6092 5661 6101 5695
rect 6101 5661 6135 5695
rect 6135 5661 6144 5695
rect 6092 5652 6144 5661
rect 7564 5652 7616 5704
rect 8760 5652 8812 5704
rect 9588 5695 9640 5704
rect 9588 5661 9597 5695
rect 9597 5661 9631 5695
rect 9631 5661 9640 5695
rect 9588 5652 9640 5661
rect 10232 5788 10284 5840
rect 10968 5788 11020 5840
rect 11796 5788 11848 5840
rect 12164 5831 12216 5840
rect 12164 5797 12173 5831
rect 12173 5797 12207 5831
rect 12207 5797 12216 5831
rect 12164 5788 12216 5797
rect 13176 5788 13228 5840
rect 16856 5788 16908 5840
rect 12532 5763 12584 5772
rect 12532 5729 12541 5763
rect 12541 5729 12575 5763
rect 12575 5729 12584 5763
rect 12532 5720 12584 5729
rect 11888 5652 11940 5704
rect 12348 5695 12400 5704
rect 12348 5661 12357 5695
rect 12357 5661 12391 5695
rect 12391 5661 12400 5695
rect 12348 5652 12400 5661
rect 12808 5695 12860 5704
rect 12808 5661 12817 5695
rect 12817 5661 12851 5695
rect 12851 5661 12860 5695
rect 12808 5652 12860 5661
rect 14096 5652 14148 5704
rect 14464 5695 14516 5704
rect 14464 5661 14473 5695
rect 14473 5661 14507 5695
rect 14507 5661 14516 5695
rect 14464 5652 14516 5661
rect 15844 5652 15896 5704
rect 16856 5695 16908 5704
rect 16856 5661 16865 5695
rect 16865 5661 16899 5695
rect 16899 5661 16908 5695
rect 16856 5652 16908 5661
rect 17316 5652 17368 5704
rect 8392 5584 8444 5636
rect 9036 5584 9088 5636
rect 12716 5584 12768 5636
rect 15200 5584 15252 5636
rect 17960 5695 18012 5704
rect 17960 5661 17969 5695
rect 17969 5661 18003 5695
rect 18003 5661 18012 5695
rect 17960 5652 18012 5661
rect 18420 5899 18472 5908
rect 18420 5865 18429 5899
rect 18429 5865 18463 5899
rect 18463 5865 18472 5899
rect 18420 5856 18472 5865
rect 18696 5788 18748 5840
rect 20260 5763 20312 5772
rect 20260 5729 20269 5763
rect 20269 5729 20303 5763
rect 20303 5729 20312 5763
rect 20260 5720 20312 5729
rect 6000 5559 6052 5568
rect 6000 5525 6009 5559
rect 6009 5525 6043 5559
rect 6043 5525 6052 5559
rect 6000 5516 6052 5525
rect 6644 5516 6696 5568
rect 11888 5559 11940 5568
rect 11888 5525 11897 5559
rect 11897 5525 11931 5559
rect 11931 5525 11940 5559
rect 11888 5516 11940 5525
rect 16672 5516 16724 5568
rect 17316 5516 17368 5568
rect 18604 5584 18656 5636
rect 20352 5695 20404 5704
rect 20352 5661 20361 5695
rect 20361 5661 20395 5695
rect 20395 5661 20404 5695
rect 20352 5652 20404 5661
rect 20720 5720 20772 5772
rect 21272 5788 21324 5840
rect 23204 5856 23256 5908
rect 22192 5788 22244 5840
rect 22376 5788 22428 5840
rect 23572 5788 23624 5840
rect 24308 5788 24360 5840
rect 19892 5584 19944 5636
rect 21640 5695 21692 5704
rect 21640 5661 21649 5695
rect 21649 5661 21683 5695
rect 21683 5661 21692 5695
rect 21640 5652 21692 5661
rect 22284 5720 22336 5772
rect 25228 5720 25280 5772
rect 21180 5627 21232 5636
rect 21180 5593 21189 5627
rect 21189 5593 21223 5627
rect 21223 5593 21232 5627
rect 21180 5584 21232 5593
rect 22192 5695 22244 5704
rect 22192 5661 22201 5695
rect 22201 5661 22235 5695
rect 22235 5661 22244 5695
rect 22192 5652 22244 5661
rect 22928 5652 22980 5704
rect 23756 5695 23808 5704
rect 23756 5661 23765 5695
rect 23765 5661 23799 5695
rect 23799 5661 23808 5695
rect 23756 5652 23808 5661
rect 24032 5695 24084 5704
rect 24032 5661 24041 5695
rect 24041 5661 24075 5695
rect 24075 5661 24084 5695
rect 24032 5652 24084 5661
rect 24952 5695 25004 5704
rect 24952 5661 24994 5695
rect 24994 5661 25004 5695
rect 24952 5652 25004 5661
rect 18052 5559 18104 5568
rect 18052 5525 18061 5559
rect 18061 5525 18095 5559
rect 18095 5525 18104 5559
rect 18052 5516 18104 5525
rect 20444 5516 20496 5568
rect 20904 5516 20956 5568
rect 22560 5584 22612 5636
rect 23204 5516 23256 5568
rect 23480 5516 23532 5568
rect 24860 5559 24912 5568
rect 24860 5525 24869 5559
rect 24869 5525 24903 5559
rect 24903 5525 24912 5559
rect 24860 5516 24912 5525
rect 25044 5559 25096 5568
rect 25044 5525 25053 5559
rect 25053 5525 25087 5559
rect 25087 5525 25096 5559
rect 25044 5516 25096 5525
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 6092 5312 6144 5364
rect 10508 5312 10560 5364
rect 11796 5312 11848 5364
rect 11888 5355 11940 5364
rect 11888 5321 11897 5355
rect 11897 5321 11931 5355
rect 11931 5321 11940 5355
rect 11888 5312 11940 5321
rect 12072 5312 12124 5364
rect 4804 5244 4856 5296
rect 4712 5176 4764 5228
rect 5724 5219 5776 5228
rect 5724 5185 5733 5219
rect 5733 5185 5767 5219
rect 5767 5185 5776 5219
rect 5724 5176 5776 5185
rect 5908 5176 5960 5228
rect 6644 5219 6696 5228
rect 6644 5185 6653 5219
rect 6653 5185 6687 5219
rect 6687 5185 6696 5219
rect 6644 5176 6696 5185
rect 6736 5219 6788 5228
rect 6736 5185 6745 5219
rect 6745 5185 6779 5219
rect 6779 5185 6788 5219
rect 6736 5176 6788 5185
rect 7932 5219 7984 5228
rect 7932 5185 7941 5219
rect 7941 5185 7975 5219
rect 7975 5185 7984 5219
rect 7932 5176 7984 5185
rect 6828 5108 6880 5160
rect 8760 5219 8812 5228
rect 8760 5185 8769 5219
rect 8769 5185 8803 5219
rect 8803 5185 8812 5219
rect 8760 5176 8812 5185
rect 9772 5176 9824 5228
rect 11704 5219 11756 5228
rect 11704 5185 11713 5219
rect 11713 5185 11747 5219
rect 11747 5185 11756 5219
rect 11704 5176 11756 5185
rect 12072 5219 12124 5228
rect 12072 5185 12081 5219
rect 12081 5185 12115 5219
rect 12115 5185 12124 5219
rect 12072 5176 12124 5185
rect 12900 5176 12952 5228
rect 4804 5040 4856 5092
rect 11060 5040 11112 5092
rect 4896 5015 4948 5024
rect 4896 4981 4905 5015
rect 4905 4981 4939 5015
rect 4939 4981 4948 5015
rect 4896 4972 4948 4981
rect 5448 5015 5500 5024
rect 5448 4981 5457 5015
rect 5457 4981 5491 5015
rect 5491 4981 5500 5015
rect 5448 4972 5500 4981
rect 8484 5015 8536 5024
rect 8484 4981 8493 5015
rect 8493 4981 8527 5015
rect 8527 4981 8536 5015
rect 8484 4972 8536 4981
rect 11520 5015 11572 5024
rect 11520 4981 11529 5015
rect 11529 4981 11563 5015
rect 11563 4981 11572 5015
rect 11520 4972 11572 4981
rect 11888 4972 11940 5024
rect 12532 5040 12584 5092
rect 13728 5219 13780 5228
rect 13728 5185 13737 5219
rect 13737 5185 13771 5219
rect 13771 5185 13780 5219
rect 13728 5176 13780 5185
rect 13912 5176 13964 5228
rect 14372 5176 14424 5228
rect 17960 5312 18012 5364
rect 16304 5219 16356 5228
rect 16304 5185 16313 5219
rect 16313 5185 16347 5219
rect 16347 5185 16356 5219
rect 16304 5176 16356 5185
rect 16672 5219 16724 5228
rect 16672 5185 16681 5219
rect 16681 5185 16715 5219
rect 16715 5185 16724 5219
rect 16672 5176 16724 5185
rect 17224 5176 17276 5228
rect 17592 5176 17644 5228
rect 18052 5219 18104 5228
rect 18052 5185 18061 5219
rect 18061 5185 18095 5219
rect 18095 5185 18104 5219
rect 18052 5176 18104 5185
rect 18696 5312 18748 5364
rect 19892 5355 19944 5364
rect 19892 5321 19901 5355
rect 19901 5321 19935 5355
rect 19935 5321 19944 5355
rect 19892 5312 19944 5321
rect 22100 5312 22152 5364
rect 21916 5244 21968 5296
rect 19800 5219 19852 5228
rect 19800 5185 19809 5219
rect 19809 5185 19843 5219
rect 19843 5185 19852 5219
rect 19800 5176 19852 5185
rect 19984 5219 20036 5228
rect 19984 5185 19993 5219
rect 19993 5185 20027 5219
rect 20027 5185 20036 5219
rect 19984 5176 20036 5185
rect 16488 5040 16540 5092
rect 13912 4972 13964 5024
rect 14004 5015 14056 5024
rect 14004 4981 14013 5015
rect 14013 4981 14047 5015
rect 14047 4981 14056 5015
rect 14004 4972 14056 4981
rect 22376 5176 22428 5228
rect 22560 5219 22612 5228
rect 22560 5185 22569 5219
rect 22569 5185 22603 5219
rect 22603 5185 22612 5219
rect 22560 5176 22612 5185
rect 22928 5355 22980 5364
rect 22928 5321 22937 5355
rect 22937 5321 22971 5355
rect 22971 5321 22980 5355
rect 22928 5312 22980 5321
rect 24032 5312 24084 5364
rect 25320 5355 25372 5364
rect 25320 5321 25329 5355
rect 25329 5321 25363 5355
rect 25363 5321 25372 5355
rect 25320 5312 25372 5321
rect 23756 5176 23808 5228
rect 24860 5219 24912 5228
rect 24860 5185 24869 5219
rect 24869 5185 24903 5219
rect 24903 5185 24912 5219
rect 24860 5176 24912 5185
rect 25136 5219 25188 5228
rect 25136 5185 25145 5219
rect 25145 5185 25179 5219
rect 25179 5185 25188 5219
rect 25136 5176 25188 5185
rect 22928 5108 22980 5160
rect 23204 5151 23256 5160
rect 23204 5117 23213 5151
rect 23213 5117 23247 5151
rect 23247 5117 23256 5151
rect 23204 5108 23256 5117
rect 18328 5040 18380 5092
rect 19984 5040 20036 5092
rect 22100 5040 22152 5092
rect 17592 4972 17644 5024
rect 21824 4972 21876 5024
rect 22376 5015 22428 5024
rect 22376 4981 22385 5015
rect 22385 4981 22419 5015
rect 22419 4981 22428 5015
rect 22376 4972 22428 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 7656 4768 7708 4820
rect 10692 4768 10744 4820
rect 16304 4768 16356 4820
rect 19800 4768 19852 4820
rect 20444 4811 20496 4820
rect 20444 4777 20453 4811
rect 20453 4777 20487 4811
rect 20487 4777 20496 4811
rect 20444 4768 20496 4777
rect 22376 4768 22428 4820
rect 23572 4768 23624 4820
rect 24308 4768 24360 4820
rect 25044 4768 25096 4820
rect 6552 4743 6604 4752
rect 6552 4709 6561 4743
rect 6561 4709 6595 4743
rect 6595 4709 6604 4743
rect 6552 4700 6604 4709
rect 5724 4632 5776 4684
rect 10968 4700 11020 4752
rect 4620 4564 4672 4616
rect 4896 4564 4948 4616
rect 5448 4607 5500 4616
rect 5448 4573 5457 4607
rect 5457 4573 5491 4607
rect 5491 4573 5500 4607
rect 5448 4564 5500 4573
rect 6184 4607 6236 4616
rect 6184 4573 6193 4607
rect 6193 4573 6227 4607
rect 6227 4573 6236 4607
rect 6184 4564 6236 4573
rect 7472 4607 7524 4616
rect 7472 4573 7481 4607
rect 7481 4573 7515 4607
rect 7515 4573 7524 4607
rect 7472 4564 7524 4573
rect 7656 4496 7708 4548
rect 8484 4496 8536 4548
rect 9588 4632 9640 4684
rect 12348 4632 12400 4684
rect 21916 4700 21968 4752
rect 25504 4700 25556 4752
rect 9588 4496 9640 4548
rect 10508 4607 10560 4616
rect 10508 4573 10517 4607
rect 10517 4573 10551 4607
rect 10551 4573 10560 4607
rect 10508 4564 10560 4573
rect 10692 4607 10744 4616
rect 10692 4573 10701 4607
rect 10701 4573 10735 4607
rect 10735 4573 10744 4607
rect 10692 4564 10744 4573
rect 14004 4496 14056 4548
rect 18328 4632 18380 4684
rect 20536 4675 20588 4684
rect 20536 4641 20545 4675
rect 20545 4641 20579 4675
rect 20579 4641 20588 4675
rect 20536 4632 20588 4641
rect 25136 4632 25188 4684
rect 15568 4607 15620 4616
rect 15568 4573 15577 4607
rect 15577 4573 15611 4607
rect 15611 4573 15620 4607
rect 15568 4564 15620 4573
rect 15660 4607 15712 4616
rect 15660 4573 15669 4607
rect 15669 4573 15703 4607
rect 15703 4573 15712 4607
rect 15660 4564 15712 4573
rect 8024 4428 8076 4480
rect 9496 4471 9548 4480
rect 9496 4437 9505 4471
rect 9505 4437 9539 4471
rect 9539 4437 9548 4471
rect 9496 4428 9548 4437
rect 11152 4428 11204 4480
rect 11520 4428 11572 4480
rect 12808 4428 12860 4480
rect 16488 4607 16540 4616
rect 16488 4573 16497 4607
rect 16497 4573 16531 4607
rect 16531 4573 16540 4607
rect 16488 4564 16540 4573
rect 20076 4564 20128 4616
rect 20260 4607 20312 4616
rect 20260 4573 20269 4607
rect 20269 4573 20303 4607
rect 20303 4573 20312 4607
rect 20260 4564 20312 4573
rect 21732 4564 21784 4616
rect 24400 4607 24452 4616
rect 24400 4573 24409 4607
rect 24409 4573 24443 4607
rect 24443 4573 24452 4607
rect 24400 4564 24452 4573
rect 24676 4564 24728 4616
rect 16212 4428 16264 4480
rect 20628 4428 20680 4480
rect 21640 4428 21692 4480
rect 21824 4428 21876 4480
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 6552 4224 6604 4276
rect 8024 4156 8076 4208
rect 9956 4224 10008 4276
rect 10232 4156 10284 4208
rect 9956 4131 10008 4140
rect 9956 4097 9965 4131
rect 9965 4097 9999 4131
rect 9999 4097 10008 4131
rect 9956 4088 10008 4097
rect 10784 4088 10836 4140
rect 10876 4131 10928 4140
rect 10876 4097 10885 4131
rect 10885 4097 10919 4131
rect 10919 4097 10928 4131
rect 10876 4088 10928 4097
rect 11704 4224 11756 4276
rect 12808 4224 12860 4276
rect 13452 4224 13504 4276
rect 14556 4224 14608 4276
rect 19800 4224 19852 4276
rect 20076 4224 20128 4276
rect 20352 4224 20404 4276
rect 20536 4224 20588 4276
rect 11612 4156 11664 4208
rect 17776 4156 17828 4208
rect 20444 4156 20496 4208
rect 11152 4131 11204 4140
rect 11152 4097 11161 4131
rect 11161 4097 11195 4131
rect 11195 4097 11204 4131
rect 11152 4088 11204 4097
rect 10416 3995 10468 4004
rect 10416 3961 10425 3995
rect 10425 3961 10459 3995
rect 10459 3961 10468 3995
rect 10416 3952 10468 3961
rect 11428 4020 11480 4072
rect 13268 4088 13320 4140
rect 15200 4131 15252 4140
rect 15200 4097 15209 4131
rect 15209 4097 15243 4131
rect 15243 4097 15252 4131
rect 15200 4088 15252 4097
rect 15292 4131 15344 4140
rect 15292 4097 15301 4131
rect 15301 4097 15335 4131
rect 15335 4097 15344 4131
rect 15292 4088 15344 4097
rect 15476 4131 15528 4140
rect 15476 4097 15485 4131
rect 15485 4097 15519 4131
rect 15519 4097 15528 4131
rect 15476 4088 15528 4097
rect 15660 4088 15712 4140
rect 17224 4088 17276 4140
rect 15384 4020 15436 4072
rect 16580 4020 16632 4072
rect 17592 4088 17644 4140
rect 19708 4088 19760 4140
rect 20076 4131 20128 4140
rect 20076 4097 20085 4131
rect 20085 4097 20119 4131
rect 20119 4097 20128 4131
rect 20076 4088 20128 4097
rect 20260 4131 20312 4140
rect 20260 4097 20269 4131
rect 20269 4097 20303 4131
rect 20303 4097 20312 4131
rect 20260 4088 20312 4097
rect 20536 4131 20588 4140
rect 20536 4097 20545 4131
rect 20545 4097 20579 4131
rect 20579 4097 20588 4131
rect 20536 4088 20588 4097
rect 22284 4131 22336 4140
rect 22284 4097 22293 4131
rect 22293 4097 22327 4131
rect 22327 4097 22336 4131
rect 22284 4088 22336 4097
rect 22376 4088 22428 4140
rect 23204 4131 23256 4140
rect 23204 4097 23213 4131
rect 23213 4097 23247 4131
rect 23247 4097 23256 4131
rect 23204 4088 23256 4097
rect 21824 4063 21876 4072
rect 21824 4029 21833 4063
rect 21833 4029 21867 4063
rect 21867 4029 21876 4063
rect 21824 4020 21876 4029
rect 10508 3884 10560 3936
rect 10692 3884 10744 3936
rect 17684 3952 17736 4004
rect 20628 3952 20680 4004
rect 21456 3952 21508 4004
rect 23480 4131 23532 4140
rect 23480 4097 23489 4131
rect 23489 4097 23523 4131
rect 23523 4097 23532 4131
rect 23480 4088 23532 4097
rect 24308 4131 24360 4140
rect 24308 4097 24317 4131
rect 24317 4097 24351 4131
rect 24351 4097 24360 4131
rect 24308 4088 24360 4097
rect 23664 4063 23716 4072
rect 23664 4029 23673 4063
rect 23673 4029 23707 4063
rect 23707 4029 23716 4063
rect 23664 4020 23716 4029
rect 24676 4131 24728 4140
rect 24676 4097 24685 4131
rect 24685 4097 24719 4131
rect 24719 4097 24728 4131
rect 24676 4088 24728 4097
rect 25136 4224 25188 4276
rect 24952 4088 25004 4140
rect 23480 3952 23532 4004
rect 25504 4131 25556 4140
rect 25504 4097 25513 4131
rect 25513 4097 25547 4131
rect 25547 4097 25556 4131
rect 25504 4088 25556 4097
rect 11796 3927 11848 3936
rect 11796 3893 11805 3927
rect 11805 3893 11839 3927
rect 11839 3893 11848 3927
rect 11796 3884 11848 3893
rect 16580 3884 16632 3936
rect 16948 3927 17000 3936
rect 16948 3893 16957 3927
rect 16957 3893 16991 3927
rect 16991 3893 17000 3927
rect 16948 3884 17000 3893
rect 24400 3884 24452 3936
rect 24860 3927 24912 3936
rect 24860 3893 24869 3927
rect 24869 3893 24903 3927
rect 24903 3893 24912 3927
rect 24860 3884 24912 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 10140 3680 10192 3732
rect 15200 3612 15252 3664
rect 15384 3612 15436 3664
rect 10416 3544 10468 3596
rect 9036 3519 9088 3528
rect 9036 3485 9045 3519
rect 9045 3485 9079 3519
rect 9079 3485 9088 3519
rect 9036 3476 9088 3485
rect 9496 3476 9548 3528
rect 11244 3519 11296 3528
rect 11244 3485 11253 3519
rect 11253 3485 11287 3519
rect 11287 3485 11296 3519
rect 11244 3476 11296 3485
rect 11428 3519 11480 3528
rect 11428 3485 11437 3519
rect 11437 3485 11471 3519
rect 11471 3485 11480 3519
rect 11428 3476 11480 3485
rect 11888 3519 11940 3528
rect 11888 3485 11897 3519
rect 11897 3485 11931 3519
rect 11931 3485 11940 3519
rect 11888 3476 11940 3485
rect 11152 3408 11204 3460
rect 13452 3476 13504 3528
rect 13544 3519 13596 3528
rect 13544 3485 13553 3519
rect 13553 3485 13587 3519
rect 13587 3485 13596 3519
rect 13544 3476 13596 3485
rect 16028 3544 16080 3596
rect 16304 3680 16356 3732
rect 18880 3680 18932 3732
rect 19800 3723 19852 3732
rect 19800 3689 19809 3723
rect 19809 3689 19843 3723
rect 19843 3689 19852 3723
rect 19800 3680 19852 3689
rect 20444 3723 20496 3732
rect 20444 3689 20453 3723
rect 20453 3689 20487 3723
rect 20487 3689 20496 3723
rect 20444 3680 20496 3689
rect 21916 3723 21968 3732
rect 21916 3689 21925 3723
rect 21925 3689 21959 3723
rect 21959 3689 21968 3723
rect 21916 3680 21968 3689
rect 23204 3680 23256 3732
rect 25504 3680 25556 3732
rect 16212 3612 16264 3664
rect 13268 3408 13320 3460
rect 14556 3519 14608 3528
rect 14556 3485 14565 3519
rect 14565 3485 14599 3519
rect 14599 3485 14608 3519
rect 14556 3476 14608 3485
rect 13728 3408 13780 3460
rect 10876 3340 10928 3392
rect 13544 3340 13596 3392
rect 15660 3476 15712 3528
rect 16304 3476 16356 3528
rect 16396 3519 16448 3528
rect 16396 3485 16405 3519
rect 16405 3485 16439 3519
rect 16439 3485 16448 3519
rect 16396 3476 16448 3485
rect 16948 3544 17000 3596
rect 16580 3476 16632 3528
rect 21272 3612 21324 3664
rect 15568 3408 15620 3460
rect 18420 3544 18472 3596
rect 20628 3587 20680 3596
rect 20628 3553 20637 3587
rect 20637 3553 20671 3587
rect 20671 3553 20680 3587
rect 20628 3544 20680 3553
rect 17316 3519 17368 3528
rect 17316 3485 17325 3519
rect 17325 3485 17359 3519
rect 17359 3485 17368 3519
rect 17316 3476 17368 3485
rect 17592 3476 17644 3528
rect 18236 3476 18288 3528
rect 20076 3519 20128 3528
rect 20076 3485 20085 3519
rect 20085 3485 20119 3519
rect 20119 3485 20128 3519
rect 20076 3476 20128 3485
rect 20260 3476 20312 3528
rect 20352 3476 20404 3528
rect 20536 3340 20588 3392
rect 21824 3544 21876 3596
rect 22376 3612 22428 3664
rect 21272 3519 21324 3528
rect 21272 3485 21281 3519
rect 21281 3485 21315 3519
rect 21315 3485 21324 3519
rect 21272 3476 21324 3485
rect 21640 3476 21692 3528
rect 22376 3519 22428 3528
rect 22376 3485 22385 3519
rect 22385 3485 22419 3519
rect 22419 3485 22428 3519
rect 22376 3476 22428 3485
rect 21456 3451 21508 3460
rect 21456 3417 21465 3451
rect 21465 3417 21499 3451
rect 21499 3417 21508 3451
rect 21456 3408 21508 3417
rect 22468 3451 22520 3460
rect 22468 3417 22477 3451
rect 22477 3417 22511 3451
rect 22511 3417 22520 3451
rect 22468 3408 22520 3417
rect 21916 3340 21968 3392
rect 23480 3408 23532 3460
rect 23664 3519 23716 3528
rect 23664 3485 23673 3519
rect 23673 3485 23707 3519
rect 23707 3485 23716 3519
rect 23664 3476 23716 3485
rect 24860 3612 24912 3664
rect 25688 3612 25740 3664
rect 24676 3408 24728 3460
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 10140 3179 10192 3188
rect 10140 3145 10149 3179
rect 10149 3145 10183 3179
rect 10183 3145 10192 3179
rect 10140 3136 10192 3145
rect 11152 3136 11204 3188
rect 10508 3111 10560 3120
rect 10508 3077 10517 3111
rect 10517 3077 10551 3111
rect 10551 3077 10560 3111
rect 10508 3068 10560 3077
rect 11612 3068 11664 3120
rect 9956 3000 10008 3052
rect 10232 3043 10284 3052
rect 10232 3009 10241 3043
rect 10241 3009 10275 3043
rect 10275 3009 10284 3043
rect 10232 3000 10284 3009
rect 848 2932 900 2984
rect 10416 2932 10468 2984
rect 10876 3000 10928 3052
rect 11152 3000 11204 3052
rect 11796 3000 11848 3052
rect 12072 2975 12124 2984
rect 12072 2941 12081 2975
rect 12081 2941 12115 2975
rect 12115 2941 12124 2975
rect 13268 3043 13320 3052
rect 13268 3009 13277 3043
rect 13277 3009 13311 3043
rect 13311 3009 13320 3043
rect 13268 3000 13320 3009
rect 15660 3136 15712 3188
rect 15936 3179 15988 3188
rect 15936 3145 15945 3179
rect 15945 3145 15979 3179
rect 15979 3145 15988 3179
rect 15936 3136 15988 3145
rect 16580 3136 16632 3188
rect 15292 3068 15344 3120
rect 15752 3068 15804 3120
rect 16212 3111 16264 3120
rect 16212 3077 16221 3111
rect 16221 3077 16255 3111
rect 16255 3077 16264 3111
rect 16212 3068 16264 3077
rect 20076 3136 20128 3188
rect 20168 3136 20220 3188
rect 21732 3136 21784 3188
rect 15200 3043 15252 3052
rect 15200 3009 15209 3043
rect 15209 3009 15243 3043
rect 15243 3009 15252 3043
rect 15200 3000 15252 3009
rect 15568 3043 15620 3052
rect 15568 3009 15577 3043
rect 15577 3009 15611 3043
rect 15611 3009 15620 3043
rect 15568 3000 15620 3009
rect 15660 3000 15712 3052
rect 17132 3000 17184 3052
rect 17776 3000 17828 3052
rect 18236 3000 18288 3052
rect 18420 3043 18472 3052
rect 18420 3009 18429 3043
rect 18429 3009 18463 3043
rect 18463 3009 18472 3043
rect 18420 3000 18472 3009
rect 18696 3043 18748 3052
rect 18696 3009 18705 3043
rect 18705 3009 18739 3043
rect 18739 3009 18748 3043
rect 18696 3000 18748 3009
rect 18880 3043 18932 3052
rect 18880 3009 18889 3043
rect 18889 3009 18923 3043
rect 18923 3009 18932 3043
rect 18880 3000 18932 3009
rect 12072 2932 12124 2941
rect 9956 2796 10008 2848
rect 13636 2864 13688 2916
rect 13452 2796 13504 2848
rect 17132 2907 17184 2916
rect 17132 2873 17141 2907
rect 17141 2873 17175 2907
rect 17175 2873 17184 2907
rect 17132 2864 17184 2873
rect 17500 2975 17552 2984
rect 17500 2941 17509 2975
rect 17509 2941 17543 2975
rect 17543 2941 17552 2975
rect 17500 2932 17552 2941
rect 18696 2864 18748 2916
rect 22468 3136 22520 3188
rect 23664 3136 23716 3188
rect 21916 2975 21968 2984
rect 21916 2941 21925 2975
rect 21925 2941 21959 2975
rect 21959 2941 21968 2975
rect 21916 2932 21968 2941
rect 27528 2975 27580 2984
rect 27528 2941 27537 2975
rect 27537 2941 27571 2975
rect 27571 2941 27580 2975
rect 27528 2932 27580 2941
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 10416 2635 10468 2644
rect 10416 2601 10425 2635
rect 10425 2601 10459 2635
rect 10459 2601 10468 2635
rect 10416 2592 10468 2601
rect 12072 2635 12124 2644
rect 12072 2601 12081 2635
rect 12081 2601 12115 2635
rect 12115 2601 12124 2635
rect 12072 2592 12124 2601
rect 13544 2635 13596 2644
rect 13544 2601 13553 2635
rect 13553 2601 13587 2635
rect 13587 2601 13596 2635
rect 13544 2592 13596 2601
rect 16396 2592 16448 2644
rect 18696 2592 18748 2644
rect 15200 2524 15252 2576
rect 10968 2456 11020 2508
rect 15752 2567 15804 2576
rect 15752 2533 15761 2567
rect 15761 2533 15795 2567
rect 15795 2533 15804 2567
rect 15752 2524 15804 2533
rect 11244 2388 11296 2440
rect 11612 2431 11664 2440
rect 11612 2397 11621 2431
rect 11621 2397 11655 2431
rect 11655 2397 11664 2431
rect 11612 2388 11664 2397
rect 13452 2431 13504 2440
rect 13452 2397 13461 2431
rect 13461 2397 13495 2431
rect 13495 2397 13504 2431
rect 13452 2388 13504 2397
rect 13636 2431 13688 2440
rect 13636 2397 13645 2431
rect 13645 2397 13679 2431
rect 13679 2397 13688 2431
rect 13636 2388 13688 2397
rect 15384 2388 15436 2440
rect 15844 2431 15896 2440
rect 15844 2397 15853 2431
rect 15853 2397 15887 2431
rect 15887 2397 15896 2431
rect 15844 2388 15896 2397
rect 16948 2388 17000 2440
rect 17776 2388 17828 2440
rect 15568 2320 15620 2372
rect 11888 2252 11940 2304
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
<< metal2 >>
rect 3238 30364 3294 31164
rect 5814 30364 5870 31164
rect 6458 30364 6514 31164
rect 7102 30364 7158 31164
rect 8390 30364 8446 31164
rect 9034 30364 9090 31164
rect 3252 28626 3280 30364
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 5828 28762 5856 30364
rect 6472 28762 6500 30364
rect 5816 28756 5868 28762
rect 5816 28698 5868 28704
rect 6460 28756 6512 28762
rect 6460 28698 6512 28704
rect 3240 28620 3292 28626
rect 3240 28562 3292 28568
rect 4620 28552 4672 28558
rect 4620 28494 4672 28500
rect 5540 28552 5592 28558
rect 5540 28494 5592 28500
rect 6184 28552 6236 28558
rect 6184 28494 6236 28500
rect 2964 28144 3016 28150
rect 2964 28086 3016 28092
rect 1768 28076 1820 28082
rect 1768 28018 1820 28024
rect 1860 28076 1912 28082
rect 1860 28018 1912 28024
rect 1400 28008 1452 28014
rect 1306 27976 1362 27985
rect 1400 27950 1452 27956
rect 1306 27911 1362 27920
rect 1214 26616 1270 26625
rect 1214 26551 1216 26560
rect 1268 26551 1270 26560
rect 1216 26522 1268 26528
rect 848 25424 900 25430
rect 846 25392 848 25401
rect 900 25392 902 25401
rect 846 25327 902 25336
rect 846 24712 902 24721
rect 846 24647 848 24656
rect 900 24647 902 24656
rect 848 24618 900 24624
rect 1214 23896 1270 23905
rect 1214 23831 1216 23840
rect 1268 23831 1270 23840
rect 1216 23802 1268 23808
rect 848 21548 900 21554
rect 848 21490 900 21496
rect 860 21321 888 21490
rect 846 21312 902 21321
rect 846 21247 902 21256
rect 1320 20058 1348 27911
rect 1412 27538 1440 27950
rect 1676 27872 1728 27878
rect 1676 27814 1728 27820
rect 1400 27532 1452 27538
rect 1400 27474 1452 27480
rect 1412 24274 1440 27474
rect 1688 27470 1716 27814
rect 1676 27464 1728 27470
rect 1676 27406 1728 27412
rect 1780 27130 1808 28018
rect 1872 27130 1900 28018
rect 2412 27532 2464 27538
rect 2412 27474 2464 27480
rect 1768 27124 1820 27130
rect 1768 27066 1820 27072
rect 1860 27124 1912 27130
rect 1860 27066 1912 27072
rect 2424 26994 2452 27474
rect 2596 27396 2648 27402
rect 2596 27338 2648 27344
rect 2608 26994 2636 27338
rect 2044 26988 2096 26994
rect 2044 26930 2096 26936
rect 2412 26988 2464 26994
rect 2412 26930 2464 26936
rect 2596 26988 2648 26994
rect 2596 26930 2648 26936
rect 2056 26874 2084 26930
rect 1964 26846 2084 26874
rect 1964 26790 1992 26846
rect 1952 26784 2004 26790
rect 1952 26726 2004 26732
rect 1860 26376 1912 26382
rect 1860 26318 1912 26324
rect 1492 26240 1544 26246
rect 1492 26182 1544 26188
rect 1504 25945 1532 26182
rect 1490 25936 1546 25945
rect 1872 25906 1900 26318
rect 1490 25871 1546 25880
rect 1860 25900 1912 25906
rect 1860 25842 1912 25848
rect 1768 25696 1820 25702
rect 1768 25638 1820 25644
rect 1780 25294 1808 25638
rect 1768 25288 1820 25294
rect 1768 25230 1820 25236
rect 1964 24886 1992 26726
rect 2608 26042 2636 26930
rect 2872 26920 2924 26926
rect 2872 26862 2924 26868
rect 2780 26240 2832 26246
rect 2780 26182 2832 26188
rect 2596 26036 2648 26042
rect 2596 25978 2648 25984
rect 2608 25922 2636 25978
rect 2792 25974 2820 26182
rect 2516 25906 2636 25922
rect 2780 25968 2832 25974
rect 2780 25910 2832 25916
rect 2504 25900 2636 25906
rect 2556 25894 2636 25900
rect 2504 25842 2556 25848
rect 2884 24970 2912 26862
rect 2976 26790 3004 28086
rect 3332 28076 3384 28082
rect 3332 28018 3384 28024
rect 3148 27668 3200 27674
rect 3148 27610 3200 27616
rect 2964 26784 3016 26790
rect 2964 26726 3016 26732
rect 3160 26382 3188 27610
rect 3344 27470 3372 28018
rect 3884 27872 3936 27878
rect 3884 27814 3936 27820
rect 3332 27464 3384 27470
rect 3332 27406 3384 27412
rect 3424 27464 3476 27470
rect 3424 27406 3476 27412
rect 3700 27464 3752 27470
rect 3700 27406 3752 27412
rect 3344 26382 3372 27406
rect 3436 27334 3464 27406
rect 3424 27328 3476 27334
rect 3424 27270 3476 27276
rect 2964 26376 3016 26382
rect 2964 26318 3016 26324
rect 3148 26376 3200 26382
rect 3148 26318 3200 26324
rect 3332 26376 3384 26382
rect 3332 26318 3384 26324
rect 2976 25906 3004 26318
rect 3436 25906 3464 27270
rect 3712 26568 3740 27406
rect 3896 27402 3924 27814
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4632 27606 4660 28494
rect 4712 28484 4764 28490
rect 4712 28426 4764 28432
rect 4724 28218 4752 28426
rect 4874 28316 5182 28325
rect 4874 28314 4880 28316
rect 4936 28314 4960 28316
rect 5016 28314 5040 28316
rect 5096 28314 5120 28316
rect 5176 28314 5182 28316
rect 4936 28262 4938 28314
rect 5118 28262 5120 28314
rect 4874 28260 4880 28262
rect 4936 28260 4960 28262
rect 5016 28260 5040 28262
rect 5096 28260 5120 28262
rect 5176 28260 5182 28262
rect 4874 28251 5182 28260
rect 4712 28212 4764 28218
rect 4712 28154 4764 28160
rect 4724 27674 4752 28154
rect 4804 28144 4856 28150
rect 4804 28086 4856 28092
rect 4816 27878 4844 28086
rect 4896 28076 4948 28082
rect 4896 28018 4948 28024
rect 4804 27872 4856 27878
rect 4804 27814 4856 27820
rect 4712 27668 4764 27674
rect 4712 27610 4764 27616
rect 4620 27600 4672 27606
rect 4620 27542 4672 27548
rect 4816 27470 4844 27814
rect 4804 27464 4856 27470
rect 4804 27406 4856 27412
rect 3884 27396 3936 27402
rect 3884 27338 3936 27344
rect 3792 27328 3844 27334
rect 4908 27316 4936 28018
rect 3792 27270 3844 27276
rect 4816 27288 4936 27316
rect 3804 27130 3832 27270
rect 3792 27124 3844 27130
rect 3792 27066 3844 27072
rect 4816 27062 4844 27288
rect 4874 27228 5182 27237
rect 4874 27226 4880 27228
rect 4936 27226 4960 27228
rect 5016 27226 5040 27228
rect 5096 27226 5120 27228
rect 5176 27226 5182 27228
rect 4936 27174 4938 27226
rect 5118 27174 5120 27226
rect 4874 27172 4880 27174
rect 4936 27172 4960 27174
rect 5016 27172 5040 27174
rect 5096 27172 5120 27174
rect 5176 27172 5182 27174
rect 4874 27163 5182 27172
rect 4160 27056 4212 27062
rect 4160 26998 4212 27004
rect 4804 27056 4856 27062
rect 4804 26998 4856 27004
rect 4172 26772 4200 26998
rect 4620 26988 4672 26994
rect 4620 26930 4672 26936
rect 3988 26744 4200 26772
rect 3792 26580 3844 26586
rect 3620 26540 3792 26568
rect 3620 25974 3648 26540
rect 3792 26522 3844 26528
rect 3700 26376 3752 26382
rect 3700 26318 3752 26324
rect 3608 25968 3660 25974
rect 3608 25910 3660 25916
rect 2964 25900 3016 25906
rect 2964 25842 3016 25848
rect 3424 25900 3476 25906
rect 3424 25842 3476 25848
rect 3240 25832 3292 25838
rect 3240 25774 3292 25780
rect 2884 24942 3096 24970
rect 1952 24880 2004 24886
rect 1952 24822 2004 24828
rect 2872 24880 2924 24886
rect 2872 24822 2924 24828
rect 2044 24608 2096 24614
rect 2044 24550 2096 24556
rect 2228 24608 2280 24614
rect 2228 24550 2280 24556
rect 1400 24268 1452 24274
rect 1400 24210 1452 24216
rect 1412 22642 1440 24210
rect 2056 24206 2084 24550
rect 2044 24200 2096 24206
rect 2044 24142 2096 24148
rect 2240 23798 2268 24550
rect 2884 24290 2912 24822
rect 2964 24812 3016 24818
rect 2964 24754 3016 24760
rect 2976 24410 3004 24754
rect 2964 24404 3016 24410
rect 2964 24346 3016 24352
rect 2884 24262 3004 24290
rect 2780 24200 2832 24206
rect 2780 24142 2832 24148
rect 2792 23866 2820 24142
rect 2780 23860 2832 23866
rect 2780 23802 2832 23808
rect 2228 23792 2280 23798
rect 2228 23734 2280 23740
rect 2976 23730 3004 24262
rect 3068 24070 3096 24942
rect 3148 24880 3200 24886
rect 3148 24822 3200 24828
rect 3160 24342 3188 24822
rect 3148 24336 3200 24342
rect 3148 24278 3200 24284
rect 3252 24206 3280 25774
rect 3712 25702 3740 26318
rect 3700 25696 3752 25702
rect 3700 25638 3752 25644
rect 3712 25294 3740 25638
rect 3700 25288 3752 25294
rect 3700 25230 3752 25236
rect 3712 24886 3740 25230
rect 3804 25226 3832 26522
rect 3884 26444 3936 26450
rect 3884 26386 3936 26392
rect 3896 26042 3924 26386
rect 3884 26036 3936 26042
rect 3884 25978 3936 25984
rect 3988 25974 4016 26744
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4632 26586 4660 26930
rect 4804 26784 4856 26790
rect 4804 26726 4856 26732
rect 5172 26784 5224 26790
rect 5172 26726 5224 26732
rect 4620 26580 4672 26586
rect 4620 26522 4672 26528
rect 4436 26376 4488 26382
rect 4436 26318 4488 26324
rect 4068 26308 4120 26314
rect 4068 26250 4120 26256
rect 4080 26042 4108 26250
rect 4068 26036 4120 26042
rect 4068 25978 4120 25984
rect 4448 25974 4476 26318
rect 3976 25968 4028 25974
rect 3976 25910 4028 25916
rect 4436 25968 4488 25974
rect 4436 25910 4488 25916
rect 3988 25786 4016 25910
rect 4632 25906 4660 26522
rect 4816 26382 4844 26726
rect 5184 26518 5212 26726
rect 5172 26512 5224 26518
rect 4986 26480 5042 26489
rect 5172 26454 5224 26460
rect 5356 26512 5408 26518
rect 5356 26454 5408 26460
rect 4986 26415 5042 26424
rect 5264 26444 5316 26450
rect 5000 26382 5028 26415
rect 5264 26386 5316 26392
rect 4804 26376 4856 26382
rect 4804 26318 4856 26324
rect 4988 26376 5040 26382
rect 4988 26318 5040 26324
rect 4712 25968 4764 25974
rect 4712 25910 4764 25916
rect 4068 25900 4120 25906
rect 4068 25842 4120 25848
rect 4620 25900 4672 25906
rect 4620 25842 4672 25848
rect 3896 25770 4016 25786
rect 3884 25764 4016 25770
rect 3936 25758 4016 25764
rect 3884 25706 3936 25712
rect 3988 25498 4016 25758
rect 3976 25492 4028 25498
rect 3976 25434 4028 25440
rect 3792 25220 3844 25226
rect 3792 25162 3844 25168
rect 3700 24880 3752 24886
rect 3700 24822 3752 24828
rect 3988 24614 4016 25434
rect 4080 25294 4108 25842
rect 4620 25764 4672 25770
rect 4620 25706 4672 25712
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4344 25424 4396 25430
rect 4344 25366 4396 25372
rect 4068 25288 4120 25294
rect 4068 25230 4120 25236
rect 4356 24750 4384 25366
rect 4632 24834 4660 25706
rect 4724 25498 4752 25910
rect 4816 25838 4844 26318
rect 4874 26140 5182 26149
rect 4874 26138 4880 26140
rect 4936 26138 4960 26140
rect 5016 26138 5040 26140
rect 5096 26138 5120 26140
rect 5176 26138 5182 26140
rect 4936 26086 4938 26138
rect 5118 26086 5120 26138
rect 4874 26084 4880 26086
rect 4936 26084 4960 26086
rect 5016 26084 5040 26086
rect 5096 26084 5120 26086
rect 5176 26084 5182 26086
rect 4874 26075 5182 26084
rect 4988 26036 5040 26042
rect 4988 25978 5040 25984
rect 4804 25832 4856 25838
rect 4804 25774 4856 25780
rect 4896 25696 4948 25702
rect 4896 25638 4948 25644
rect 4712 25492 4764 25498
rect 4712 25434 4764 25440
rect 4908 25294 4936 25638
rect 5000 25294 5028 25978
rect 5276 25888 5304 26386
rect 5368 25974 5396 26454
rect 5552 26042 5580 28494
rect 6196 28218 6224 28494
rect 6552 28416 6604 28422
rect 6552 28358 6604 28364
rect 6184 28212 6236 28218
rect 6184 28154 6236 28160
rect 6564 28150 6592 28358
rect 7116 28218 7144 30364
rect 8404 28558 8432 30364
rect 9048 28762 9076 30364
rect 9036 28756 9088 28762
rect 9036 28698 9088 28704
rect 8392 28552 8444 28558
rect 8392 28494 8444 28500
rect 9128 28552 9180 28558
rect 9128 28494 9180 28500
rect 9680 28552 9732 28558
rect 9680 28494 9732 28500
rect 12532 28552 12584 28558
rect 12532 28494 12584 28500
rect 17040 28552 17092 28558
rect 17040 28494 17092 28500
rect 7748 28484 7800 28490
rect 7748 28426 7800 28432
rect 7288 28416 7340 28422
rect 7288 28358 7340 28364
rect 7104 28212 7156 28218
rect 7104 28154 7156 28160
rect 6552 28144 6604 28150
rect 6552 28086 6604 28092
rect 5632 28076 5684 28082
rect 5632 28018 5684 28024
rect 5816 28076 5868 28082
rect 5816 28018 5868 28024
rect 5908 28076 5960 28082
rect 5908 28018 5960 28024
rect 6644 28076 6696 28082
rect 6644 28018 6696 28024
rect 6736 28076 6788 28082
rect 6736 28018 6788 28024
rect 5644 26586 5672 28018
rect 5828 27878 5856 28018
rect 5816 27872 5868 27878
rect 5816 27814 5868 27820
rect 5828 26994 5856 27814
rect 5920 27606 5948 28018
rect 6276 28008 6328 28014
rect 6276 27950 6328 27956
rect 6288 27878 6316 27950
rect 6276 27872 6328 27878
rect 6276 27814 6328 27820
rect 6288 27606 6316 27814
rect 6656 27674 6684 28018
rect 6644 27668 6696 27674
rect 6644 27610 6696 27616
rect 5908 27600 5960 27606
rect 5908 27542 5960 27548
rect 6276 27600 6328 27606
rect 6276 27542 6328 27548
rect 6184 27464 6236 27470
rect 6184 27406 6236 27412
rect 5816 26988 5868 26994
rect 5816 26930 5868 26936
rect 5632 26580 5684 26586
rect 5632 26522 5684 26528
rect 5724 26376 5776 26382
rect 5724 26318 5776 26324
rect 5540 26036 5592 26042
rect 5540 25978 5592 25984
rect 5356 25968 5408 25974
rect 5356 25910 5408 25916
rect 5184 25860 5304 25888
rect 4896 25288 4948 25294
rect 4896 25230 4948 25236
rect 4988 25288 5040 25294
rect 4988 25230 5040 25236
rect 4712 25152 4764 25158
rect 5184 25140 5212 25860
rect 5264 25764 5316 25770
rect 5264 25706 5316 25712
rect 4712 25094 4764 25100
rect 4816 25112 5212 25140
rect 4540 24818 4660 24834
rect 4528 24812 4660 24818
rect 4580 24806 4660 24812
rect 4528 24754 4580 24760
rect 4724 24750 4752 25094
rect 4344 24744 4396 24750
rect 4344 24686 4396 24692
rect 4712 24744 4764 24750
rect 4712 24686 4764 24692
rect 4816 24682 4844 25112
rect 4874 25052 5182 25061
rect 4874 25050 4880 25052
rect 4936 25050 4960 25052
rect 5016 25050 5040 25052
rect 5096 25050 5120 25052
rect 5176 25050 5182 25052
rect 4936 24998 4938 25050
rect 5118 24998 5120 25050
rect 4874 24996 4880 24998
rect 4936 24996 4960 24998
rect 5016 24996 5040 24998
rect 5096 24996 5120 24998
rect 5176 24996 5182 24998
rect 4874 24987 5182 24996
rect 5276 24682 5304 25706
rect 5368 25498 5396 25910
rect 5356 25492 5408 25498
rect 5356 25434 5408 25440
rect 5448 25288 5500 25294
rect 5448 25230 5500 25236
rect 5632 25288 5684 25294
rect 5736 25276 5764 26318
rect 5828 25514 5856 26930
rect 5908 26308 5960 26314
rect 5908 26250 5960 26256
rect 5920 26042 5948 26250
rect 6000 26240 6052 26246
rect 6000 26182 6052 26188
rect 5908 26036 5960 26042
rect 5908 25978 5960 25984
rect 6012 25838 6040 26182
rect 6000 25832 6052 25838
rect 6000 25774 6052 25780
rect 6196 25770 6224 27406
rect 6288 26382 6316 27542
rect 6368 27328 6420 27334
rect 6368 27270 6420 27276
rect 6380 26450 6408 27270
rect 6644 26988 6696 26994
rect 6644 26930 6696 26936
rect 6460 26580 6512 26586
rect 6460 26522 6512 26528
rect 6368 26444 6420 26450
rect 6368 26386 6420 26392
rect 6276 26376 6328 26382
rect 6276 26318 6328 26324
rect 6472 26364 6500 26522
rect 6552 26376 6604 26382
rect 6472 26336 6552 26364
rect 6368 26308 6420 26314
rect 6368 26250 6420 26256
rect 6276 25900 6328 25906
rect 6276 25842 6328 25848
rect 6184 25764 6236 25770
rect 6184 25706 6236 25712
rect 5828 25498 5948 25514
rect 5828 25492 5960 25498
rect 5828 25486 5908 25492
rect 5908 25434 5960 25440
rect 6184 25492 6236 25498
rect 6184 25434 6236 25440
rect 6196 25294 6224 25434
rect 5816 25288 5868 25294
rect 5736 25248 5816 25276
rect 5632 25230 5684 25236
rect 5816 25230 5868 25236
rect 6184 25288 6236 25294
rect 6184 25230 6236 25236
rect 5356 25152 5408 25158
rect 5356 25094 5408 25100
rect 5368 24818 5396 25094
rect 5356 24812 5408 24818
rect 5356 24754 5408 24760
rect 5460 24750 5488 25230
rect 5644 25140 5672 25230
rect 5644 25112 5856 25140
rect 5828 24818 5856 25112
rect 6288 24818 6316 25842
rect 6380 24818 6408 26250
rect 6472 25974 6500 26336
rect 6552 26318 6604 26324
rect 6656 26246 6684 26930
rect 6748 26586 6776 28018
rect 6828 27396 6880 27402
rect 6828 27338 6880 27344
rect 6736 26580 6788 26586
rect 6736 26522 6788 26528
rect 6644 26240 6696 26246
rect 6644 26182 6696 26188
rect 6460 25968 6512 25974
rect 6460 25910 6512 25916
rect 6552 25900 6604 25906
rect 6656 25888 6684 26182
rect 6736 26036 6788 26042
rect 6736 25978 6788 25984
rect 6604 25860 6684 25888
rect 6552 25842 6604 25848
rect 6552 25764 6604 25770
rect 6552 25706 6604 25712
rect 6460 24948 6512 24954
rect 6460 24890 6512 24896
rect 5816 24812 5868 24818
rect 5816 24754 5868 24760
rect 6276 24812 6328 24818
rect 6276 24754 6328 24760
rect 6368 24812 6420 24818
rect 6368 24754 6420 24760
rect 5448 24744 5500 24750
rect 5448 24686 5500 24692
rect 4804 24676 4856 24682
rect 4804 24618 4856 24624
rect 5264 24676 5316 24682
rect 5264 24618 5316 24624
rect 3424 24608 3476 24614
rect 3424 24550 3476 24556
rect 3976 24608 4028 24614
rect 3976 24550 4028 24556
rect 3436 24410 3464 24550
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 3424 24404 3476 24410
rect 3424 24346 3476 24352
rect 3240 24200 3292 24206
rect 3240 24142 3292 24148
rect 3056 24064 3108 24070
rect 3056 24006 3108 24012
rect 1952 23724 2004 23730
rect 1952 23666 2004 23672
rect 2872 23724 2924 23730
rect 2872 23666 2924 23672
rect 2964 23724 3016 23730
rect 2964 23666 3016 23672
rect 1676 23520 1728 23526
rect 1676 23462 1728 23468
rect 1400 22636 1452 22642
rect 1400 22578 1452 22584
rect 1412 22098 1440 22578
rect 1400 22092 1452 22098
rect 1400 22034 1452 22040
rect 1688 22030 1716 23462
rect 1964 23225 1992 23666
rect 2884 23322 2912 23666
rect 2872 23316 2924 23322
rect 2872 23258 2924 23264
rect 1950 23216 2006 23225
rect 3068 23186 3096 24006
rect 3252 23866 3280 24142
rect 3240 23860 3292 23866
rect 3240 23802 3292 23808
rect 3436 23662 3464 24346
rect 5460 24342 5488 24686
rect 5828 24682 5856 24754
rect 5816 24676 5868 24682
rect 5816 24618 5868 24624
rect 5448 24336 5500 24342
rect 5448 24278 5500 24284
rect 3976 24064 4028 24070
rect 3976 24006 4028 24012
rect 3988 23730 4016 24006
rect 4874 23964 5182 23973
rect 4874 23962 4880 23964
rect 4936 23962 4960 23964
rect 5016 23962 5040 23964
rect 5096 23962 5120 23964
rect 5176 23962 5182 23964
rect 4936 23910 4938 23962
rect 5118 23910 5120 23962
rect 4874 23908 4880 23910
rect 4936 23908 4960 23910
rect 5016 23908 5040 23910
rect 5096 23908 5120 23910
rect 5176 23908 5182 23910
rect 4874 23899 5182 23908
rect 5828 23866 5856 24618
rect 6380 24274 6408 24754
rect 6472 24274 6500 24890
rect 6564 24818 6592 25706
rect 6748 25362 6776 25978
rect 6840 25362 6868 27338
rect 7196 26784 7248 26790
rect 7196 26726 7248 26732
rect 7012 26512 7064 26518
rect 7104 26512 7156 26518
rect 7012 26454 7064 26460
rect 7102 26480 7104 26489
rect 7156 26480 7158 26489
rect 6920 26444 6972 26450
rect 6920 26386 6972 26392
rect 6932 25820 6960 26386
rect 7024 25974 7052 26454
rect 7102 26415 7158 26424
rect 7208 26314 7236 26726
rect 7196 26308 7248 26314
rect 7196 26250 7248 26256
rect 7208 26042 7236 26250
rect 7196 26036 7248 26042
rect 7196 25978 7248 25984
rect 7012 25968 7064 25974
rect 7012 25910 7064 25916
rect 7196 25900 7248 25906
rect 7116 25860 7196 25888
rect 7116 25820 7144 25860
rect 7196 25842 7248 25848
rect 6932 25792 7144 25820
rect 6736 25356 6788 25362
rect 6736 25298 6788 25304
rect 6828 25356 6880 25362
rect 6828 25298 6880 25304
rect 6736 25152 6788 25158
rect 6736 25094 6788 25100
rect 6748 24818 6776 25094
rect 6840 24954 6868 25298
rect 6932 25294 6960 25792
rect 7300 25362 7328 28358
rect 7760 28014 7788 28426
rect 8484 28416 8536 28422
rect 8484 28358 8536 28364
rect 8496 28150 8524 28358
rect 9140 28218 9168 28494
rect 9692 28218 9720 28494
rect 9128 28212 9180 28218
rect 9128 28154 9180 28160
rect 9680 28212 9732 28218
rect 9680 28154 9732 28160
rect 8484 28144 8536 28150
rect 8484 28086 8536 28092
rect 7748 28008 7800 28014
rect 7748 27950 7800 27956
rect 7760 27402 7788 27950
rect 9692 27538 9720 28154
rect 10416 28076 10468 28082
rect 10416 28018 10468 28024
rect 10428 27606 10456 28018
rect 10876 28008 10928 28014
rect 10876 27950 10928 27956
rect 10416 27600 10468 27606
rect 10416 27542 10468 27548
rect 10888 27538 10916 27950
rect 10968 27940 11020 27946
rect 10968 27882 11020 27888
rect 9680 27532 9732 27538
rect 9680 27474 9732 27480
rect 10876 27532 10928 27538
rect 10876 27474 10928 27480
rect 8852 27464 8904 27470
rect 8852 27406 8904 27412
rect 7472 27396 7524 27402
rect 7472 27338 7524 27344
rect 7656 27396 7708 27402
rect 7656 27338 7708 27344
rect 7748 27396 7800 27402
rect 7748 27338 7800 27344
rect 7380 26784 7432 26790
rect 7380 26726 7432 26732
rect 7392 26586 7420 26726
rect 7484 26586 7512 27338
rect 7668 27130 7696 27338
rect 8760 27328 8812 27334
rect 8760 27270 8812 27276
rect 7656 27124 7708 27130
rect 7656 27066 7708 27072
rect 8116 27056 8168 27062
rect 8116 26998 8168 27004
rect 8300 27056 8352 27062
rect 8300 26998 8352 27004
rect 7840 26784 7892 26790
rect 7840 26726 7892 26732
rect 7380 26580 7432 26586
rect 7380 26522 7432 26528
rect 7472 26580 7524 26586
rect 7472 26522 7524 26528
rect 7472 26376 7524 26382
rect 7472 26318 7524 26324
rect 7484 25770 7512 26318
rect 7472 25764 7524 25770
rect 7472 25706 7524 25712
rect 7380 25696 7432 25702
rect 7380 25638 7432 25644
rect 7392 25430 7420 25638
rect 7380 25424 7432 25430
rect 7380 25366 7432 25372
rect 7564 25424 7616 25430
rect 7564 25366 7616 25372
rect 7288 25356 7340 25362
rect 7288 25298 7340 25304
rect 6920 25288 6972 25294
rect 6920 25230 6972 25236
rect 6828 24948 6880 24954
rect 6828 24890 6880 24896
rect 6932 24818 6960 25230
rect 7392 24818 7420 25366
rect 7472 25356 7524 25362
rect 7472 25298 7524 25304
rect 6552 24812 6604 24818
rect 6552 24754 6604 24760
rect 6736 24812 6788 24818
rect 6736 24754 6788 24760
rect 6828 24812 6880 24818
rect 6828 24754 6880 24760
rect 6920 24812 6972 24818
rect 6920 24754 6972 24760
rect 7380 24812 7432 24818
rect 7380 24754 7432 24760
rect 6564 24682 6592 24754
rect 6840 24682 6868 24754
rect 6552 24676 6604 24682
rect 6552 24618 6604 24624
rect 6828 24676 6880 24682
rect 6828 24618 6880 24624
rect 6368 24268 6420 24274
rect 6368 24210 6420 24216
rect 6460 24268 6512 24274
rect 6460 24210 6512 24216
rect 6932 24206 6960 24754
rect 7104 24608 7156 24614
rect 7104 24550 7156 24556
rect 6736 24200 6788 24206
rect 6736 24142 6788 24148
rect 6828 24200 6880 24206
rect 6828 24142 6880 24148
rect 6920 24200 6972 24206
rect 6920 24142 6972 24148
rect 6184 24064 6236 24070
rect 6184 24006 6236 24012
rect 5816 23860 5868 23866
rect 5816 23802 5868 23808
rect 3976 23724 4028 23730
rect 3976 23666 4028 23672
rect 3424 23656 3476 23662
rect 3424 23598 3476 23604
rect 1950 23151 2006 23160
rect 3056 23180 3108 23186
rect 3056 23122 3108 23128
rect 3436 23118 3464 23598
rect 3988 23322 4016 23666
rect 4804 23656 4856 23662
rect 4804 23598 4856 23604
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 3976 23316 4028 23322
rect 3976 23258 4028 23264
rect 4816 23118 4844 23598
rect 6196 23526 6224 24006
rect 6184 23520 6236 23526
rect 6184 23462 6236 23468
rect 3240 23112 3292 23118
rect 3240 23054 3292 23060
rect 3424 23112 3476 23118
rect 3424 23054 3476 23060
rect 4804 23112 4856 23118
rect 4804 23054 4856 23060
rect 2688 22976 2740 22982
rect 2688 22918 2740 22924
rect 2700 22710 2728 22918
rect 2688 22704 2740 22710
rect 2688 22646 2740 22652
rect 2320 22636 2372 22642
rect 2320 22578 2372 22584
rect 2332 22094 2360 22578
rect 3252 22234 3280 23054
rect 4816 22574 4844 23054
rect 4874 22876 5182 22885
rect 4874 22874 4880 22876
rect 4936 22874 4960 22876
rect 5016 22874 5040 22876
rect 5096 22874 5120 22876
rect 5176 22874 5182 22876
rect 4936 22822 4938 22874
rect 5118 22822 5120 22874
rect 4874 22820 4880 22822
rect 4936 22820 4960 22822
rect 5016 22820 5040 22822
rect 5096 22820 5120 22822
rect 5176 22820 5182 22822
rect 4874 22811 5182 22820
rect 5448 22636 5500 22642
rect 5448 22578 5500 22584
rect 4804 22568 4856 22574
rect 4804 22510 4856 22516
rect 4712 22500 4764 22506
rect 4712 22442 4764 22448
rect 3884 22432 3936 22438
rect 3884 22374 3936 22380
rect 3240 22228 3292 22234
rect 3240 22170 3292 22176
rect 2412 22094 2464 22098
rect 2332 22092 2464 22094
rect 2332 22066 2412 22092
rect 1676 22024 1728 22030
rect 1676 21966 1728 21972
rect 2332 21554 2360 22066
rect 2412 22034 2464 22040
rect 3896 22030 3924 22374
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4724 22094 4752 22442
rect 4816 22234 4844 22510
rect 4804 22228 4856 22234
rect 4804 22170 4856 22176
rect 4724 22066 4844 22094
rect 3884 22024 3936 22030
rect 3884 21966 3936 21972
rect 2320 21548 2372 21554
rect 2320 21490 2372 21496
rect 2872 21548 2924 21554
rect 2872 21490 2924 21496
rect 1584 21344 1636 21350
rect 1584 21286 1636 21292
rect 1596 20874 1624 21286
rect 2884 21146 2912 21490
rect 4816 21486 4844 22066
rect 5264 21888 5316 21894
rect 5264 21830 5316 21836
rect 4874 21788 5182 21797
rect 4874 21786 4880 21788
rect 4936 21786 4960 21788
rect 5016 21786 5040 21788
rect 5096 21786 5120 21788
rect 5176 21786 5182 21788
rect 4936 21734 4938 21786
rect 5118 21734 5120 21786
rect 4874 21732 4880 21734
rect 4936 21732 4960 21734
rect 5016 21732 5040 21734
rect 5096 21732 5120 21734
rect 5176 21732 5182 21734
rect 4874 21723 5182 21732
rect 5276 21622 5304 21830
rect 5460 21690 5488 22578
rect 6748 22574 6776 24142
rect 6840 23118 6868 24142
rect 7116 24138 7144 24550
rect 7104 24132 7156 24138
rect 7104 24074 7156 24080
rect 6920 23724 6972 23730
rect 6920 23666 6972 23672
rect 6828 23112 6880 23118
rect 6828 23054 6880 23060
rect 6840 22642 6868 23054
rect 6932 22778 6960 23666
rect 7116 23594 7144 24074
rect 7196 24064 7248 24070
rect 7196 24006 7248 24012
rect 7208 23866 7236 24006
rect 7196 23860 7248 23866
rect 7196 23802 7248 23808
rect 7380 23656 7432 23662
rect 7380 23598 7432 23604
rect 7104 23588 7156 23594
rect 7104 23530 7156 23536
rect 7288 23044 7340 23050
rect 7288 22986 7340 22992
rect 6920 22772 6972 22778
rect 6920 22714 6972 22720
rect 6828 22636 6880 22642
rect 6828 22578 6880 22584
rect 6736 22568 6788 22574
rect 6736 22510 6788 22516
rect 6736 21888 6788 21894
rect 6736 21830 6788 21836
rect 5448 21684 5500 21690
rect 5448 21626 5500 21632
rect 5264 21616 5316 21622
rect 5264 21558 5316 21564
rect 4804 21480 4856 21486
rect 4804 21422 4856 21428
rect 5264 21480 5316 21486
rect 5264 21422 5316 21428
rect 5724 21480 5776 21486
rect 6748 21434 6776 21830
rect 6840 21593 6868 22578
rect 7300 22574 7328 22986
rect 7392 22574 7420 23598
rect 7288 22568 7340 22574
rect 7288 22510 7340 22516
rect 7380 22568 7432 22574
rect 7380 22510 7432 22516
rect 6920 22228 6972 22234
rect 6920 22170 6972 22176
rect 6932 21622 6960 22170
rect 7012 22092 7064 22098
rect 7064 22052 7144 22080
rect 7012 22034 7064 22040
rect 7012 21956 7064 21962
rect 7012 21898 7064 21904
rect 6920 21616 6972 21622
rect 6826 21584 6882 21593
rect 6920 21558 6972 21564
rect 6826 21519 6882 21528
rect 5724 21422 5776 21428
rect 4620 21344 4672 21350
rect 4620 21286 4672 21292
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 2872 21140 2924 21146
rect 2872 21082 2924 21088
rect 4632 20874 4660 21286
rect 5276 20942 5304 21422
rect 5448 21412 5500 21418
rect 5448 21354 5500 21360
rect 5460 21010 5488 21354
rect 5736 21146 5764 21422
rect 6656 21418 6776 21434
rect 6644 21412 6776 21418
rect 6696 21406 6776 21412
rect 6644 21354 6696 21360
rect 5724 21140 5776 21146
rect 5724 21082 5776 21088
rect 5448 21004 5500 21010
rect 5448 20946 5500 20952
rect 5264 20936 5316 20942
rect 5264 20878 5316 20884
rect 5356 20936 5408 20942
rect 5356 20878 5408 20884
rect 1584 20868 1636 20874
rect 1584 20810 1636 20816
rect 4620 20868 4672 20874
rect 4620 20810 4672 20816
rect 2780 20800 2832 20806
rect 2780 20742 2832 20748
rect 5264 20800 5316 20806
rect 5264 20742 5316 20748
rect 2688 20256 2740 20262
rect 2688 20198 2740 20204
rect 1308 20052 1360 20058
rect 1308 19994 1360 20000
rect 846 19952 902 19961
rect 846 19887 902 19896
rect 860 19854 888 19887
rect 848 19848 900 19854
rect 848 19790 900 19796
rect 2700 19786 2728 20198
rect 2792 19854 2820 20742
rect 4874 20700 5182 20709
rect 4874 20698 4880 20700
rect 4936 20698 4960 20700
rect 5016 20698 5040 20700
rect 5096 20698 5120 20700
rect 5176 20698 5182 20700
rect 4936 20646 4938 20698
rect 5118 20646 5120 20698
rect 4874 20644 4880 20646
rect 4936 20644 4960 20646
rect 5016 20644 5040 20646
rect 5096 20644 5120 20646
rect 5176 20644 5182 20646
rect 4874 20635 5182 20644
rect 5276 20466 5304 20742
rect 5368 20602 5396 20878
rect 5356 20596 5408 20602
rect 5356 20538 5408 20544
rect 5736 20534 5764 21082
rect 6748 21078 6776 21406
rect 6840 21146 6868 21519
rect 6920 21480 6972 21486
rect 6920 21422 6972 21428
rect 6828 21140 6880 21146
rect 6828 21082 6880 21088
rect 6736 21072 6788 21078
rect 6736 21014 6788 21020
rect 6276 20800 6328 20806
rect 6276 20742 6328 20748
rect 6000 20596 6052 20602
rect 6000 20538 6052 20544
rect 5724 20528 5776 20534
rect 5724 20470 5776 20476
rect 3884 20460 3936 20466
rect 3884 20402 3936 20408
rect 5264 20460 5316 20466
rect 5264 20402 5316 20408
rect 3240 20392 3292 20398
rect 3240 20334 3292 20340
rect 2780 19848 2832 19854
rect 2780 19790 2832 19796
rect 2688 19780 2740 19786
rect 2688 19722 2740 19728
rect 1676 19712 1728 19718
rect 1676 19654 1728 19660
rect 1688 19378 1716 19654
rect 2792 19446 2820 19790
rect 2780 19440 2832 19446
rect 2780 19382 2832 19388
rect 1676 19372 1728 19378
rect 1676 19314 1728 19320
rect 2320 18284 2372 18290
rect 2372 18244 2452 18272
rect 2320 18226 2372 18232
rect 2320 17604 2372 17610
rect 2320 17546 2372 17552
rect 1952 17196 2004 17202
rect 1952 17138 2004 17144
rect 1964 16794 1992 17138
rect 1952 16788 2004 16794
rect 1952 16730 2004 16736
rect 2332 16522 2360 17546
rect 2424 16998 2452 18244
rect 2412 16992 2464 16998
rect 2412 16934 2464 16940
rect 2320 16516 2372 16522
rect 2320 16458 2372 16464
rect 2332 16402 2360 16458
rect 2056 16374 2360 16402
rect 2056 15026 2084 16374
rect 2320 16244 2372 16250
rect 2320 16186 2372 16192
rect 2332 15026 2360 16186
rect 1952 15020 2004 15026
rect 1952 14962 2004 14968
rect 2044 15020 2096 15026
rect 2044 14962 2096 14968
rect 2320 15020 2372 15026
rect 2320 14962 2372 14968
rect 1964 14618 1992 14962
rect 1952 14612 2004 14618
rect 1952 14554 2004 14560
rect 1860 14408 1912 14414
rect 1860 14350 1912 14356
rect 1400 14340 1452 14346
rect 1400 14282 1452 14288
rect 1412 13938 1440 14282
rect 1768 14272 1820 14278
rect 1768 14214 1820 14220
rect 1780 13938 1808 14214
rect 1400 13932 1452 13938
rect 1400 13874 1452 13880
rect 1492 13932 1544 13938
rect 1492 13874 1544 13880
rect 1676 13932 1728 13938
rect 1676 13874 1728 13880
rect 1768 13932 1820 13938
rect 1768 13874 1820 13880
rect 1412 13258 1440 13874
rect 1504 13326 1532 13874
rect 1688 13734 1716 13874
rect 1676 13728 1728 13734
rect 1676 13670 1728 13676
rect 1688 13530 1716 13670
rect 1676 13524 1728 13530
rect 1676 13466 1728 13472
rect 1872 13462 1900 14350
rect 2056 13870 2084 14962
rect 2136 14408 2188 14414
rect 2136 14350 2188 14356
rect 2148 14074 2176 14350
rect 2228 14272 2280 14278
rect 2228 14214 2280 14220
rect 2136 14068 2188 14074
rect 2136 14010 2188 14016
rect 2240 14006 2268 14214
rect 2228 14000 2280 14006
rect 2228 13942 2280 13948
rect 2332 13938 2360 14962
rect 2320 13932 2372 13938
rect 2320 13874 2372 13880
rect 2044 13864 2096 13870
rect 2044 13806 2096 13812
rect 1860 13456 1912 13462
rect 1860 13398 1912 13404
rect 1492 13320 1544 13326
rect 1492 13262 1544 13268
rect 1400 13252 1452 13258
rect 1400 13194 1452 13200
rect 2056 12220 2084 13806
rect 2332 12238 2360 13874
rect 2424 13870 2452 16934
rect 2596 16720 2648 16726
rect 2596 16662 2648 16668
rect 2608 16590 2636 16662
rect 2596 16584 2648 16590
rect 2596 16526 2648 16532
rect 2504 16516 2556 16522
rect 2504 16458 2556 16464
rect 2516 16250 2544 16458
rect 2504 16244 2556 16250
rect 2504 16186 2556 16192
rect 2792 15502 2820 19382
rect 3252 19378 3280 20334
rect 3896 19786 3924 20402
rect 4068 20256 4120 20262
rect 4068 20198 4120 20204
rect 5632 20256 5684 20262
rect 5632 20198 5684 20204
rect 3884 19780 3936 19786
rect 3884 19722 3936 19728
rect 3896 19378 3924 19722
rect 4080 19378 4108 20198
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4874 19612 5182 19621
rect 4874 19610 4880 19612
rect 4936 19610 4960 19612
rect 5016 19610 5040 19612
rect 5096 19610 5120 19612
rect 5176 19610 5182 19612
rect 4936 19558 4938 19610
rect 5118 19558 5120 19610
rect 4874 19556 4880 19558
rect 4936 19556 4960 19558
rect 5016 19556 5040 19558
rect 5096 19556 5120 19558
rect 5176 19556 5182 19558
rect 4874 19547 5182 19556
rect 5644 19378 5672 20198
rect 6012 19786 6040 20538
rect 6184 19916 6236 19922
rect 6184 19858 6236 19864
rect 6000 19780 6052 19786
rect 6000 19722 6052 19728
rect 6092 19780 6144 19786
rect 6092 19722 6144 19728
rect 5908 19712 5960 19718
rect 5908 19654 5960 19660
rect 5920 19378 5948 19654
rect 3240 19372 3292 19378
rect 3240 19314 3292 19320
rect 3884 19372 3936 19378
rect 3884 19314 3936 19320
rect 4068 19372 4120 19378
rect 4068 19314 4120 19320
rect 5632 19372 5684 19378
rect 5632 19314 5684 19320
rect 5908 19372 5960 19378
rect 5908 19314 5960 19320
rect 3896 18834 3924 19314
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 5264 18964 5316 18970
rect 5264 18906 5316 18912
rect 3884 18828 3936 18834
rect 3884 18770 3936 18776
rect 4804 18692 4856 18698
rect 4804 18634 4856 18640
rect 4816 18426 4844 18634
rect 4874 18524 5182 18533
rect 4874 18522 4880 18524
rect 4936 18522 4960 18524
rect 5016 18522 5040 18524
rect 5096 18522 5120 18524
rect 5176 18522 5182 18524
rect 4936 18470 4938 18522
rect 5118 18470 5120 18522
rect 4874 18468 4880 18470
rect 4936 18468 4960 18470
rect 5016 18468 5040 18470
rect 5096 18468 5120 18470
rect 5176 18468 5182 18470
rect 4874 18459 5182 18468
rect 4804 18420 4856 18426
rect 4804 18362 4856 18368
rect 4896 18420 4948 18426
rect 4896 18362 4948 18368
rect 4908 18290 4936 18362
rect 5276 18290 5304 18906
rect 6012 18766 6040 19722
rect 6104 19514 6132 19722
rect 6196 19514 6224 19858
rect 6092 19508 6144 19514
rect 6092 19450 6144 19456
rect 6184 19508 6236 19514
rect 6184 19450 6236 19456
rect 6196 19378 6224 19450
rect 6288 19378 6316 20742
rect 6840 20534 6868 21082
rect 6828 20528 6880 20534
rect 6828 20470 6880 20476
rect 6552 20460 6604 20466
rect 6552 20402 6604 20408
rect 6368 20392 6420 20398
rect 6368 20334 6420 20340
rect 6380 19990 6408 20334
rect 6564 19990 6592 20402
rect 6828 20256 6880 20262
rect 6828 20198 6880 20204
rect 6368 19984 6420 19990
rect 6368 19926 6420 19932
rect 6552 19984 6604 19990
rect 6552 19926 6604 19932
rect 6460 19712 6512 19718
rect 6460 19654 6512 19660
rect 6472 19378 6500 19654
rect 6736 19508 6788 19514
rect 6736 19450 6788 19456
rect 6748 19378 6776 19450
rect 6840 19378 6868 20198
rect 6932 19446 6960 21422
rect 7024 20602 7052 21898
rect 7116 21690 7144 22052
rect 7196 22024 7248 22030
rect 7196 21966 7248 21972
rect 7208 21690 7236 21966
rect 7104 21684 7156 21690
rect 7104 21626 7156 21632
rect 7196 21684 7248 21690
rect 7196 21626 7248 21632
rect 7102 21584 7158 21593
rect 7102 21519 7104 21528
rect 7156 21519 7158 21528
rect 7196 21548 7248 21554
rect 7104 21490 7156 21496
rect 7300 21536 7328 22510
rect 7392 21570 7420 22510
rect 7484 21690 7512 25298
rect 7576 24818 7604 25366
rect 7748 25356 7800 25362
rect 7748 25298 7800 25304
rect 7760 24818 7788 25298
rect 7564 24812 7616 24818
rect 7564 24754 7616 24760
rect 7748 24812 7800 24818
rect 7748 24754 7800 24760
rect 7760 23526 7788 24754
rect 7852 24410 7880 26726
rect 8128 26586 8156 26998
rect 8116 26580 8168 26586
rect 8116 26522 8168 26528
rect 8208 26308 8260 26314
rect 8208 26250 8260 26256
rect 8220 25906 8248 26250
rect 8208 25900 8260 25906
rect 8208 25842 8260 25848
rect 8024 25696 8076 25702
rect 8024 25638 8076 25644
rect 7932 25152 7984 25158
rect 7932 25094 7984 25100
rect 7840 24404 7892 24410
rect 7840 24346 7892 24352
rect 7748 23520 7800 23526
rect 7748 23462 7800 23468
rect 7656 22636 7708 22642
rect 7656 22578 7708 22584
rect 7668 22234 7696 22578
rect 7656 22228 7708 22234
rect 7656 22170 7708 22176
rect 7748 21956 7800 21962
rect 7748 21898 7800 21904
rect 7760 21706 7788 21898
rect 7760 21690 7880 21706
rect 7472 21684 7524 21690
rect 7472 21626 7524 21632
rect 7760 21684 7892 21690
rect 7760 21678 7840 21684
rect 7392 21554 7512 21570
rect 7392 21548 7524 21554
rect 7392 21542 7472 21548
rect 7248 21508 7328 21536
rect 7196 21490 7248 21496
rect 7472 21490 7524 21496
rect 7104 21412 7156 21418
rect 7104 21354 7156 21360
rect 7116 20874 7144 21354
rect 7208 21010 7236 21490
rect 7196 21004 7248 21010
rect 7196 20946 7248 20952
rect 7104 20868 7156 20874
rect 7104 20810 7156 20816
rect 7012 20596 7064 20602
rect 7012 20538 7064 20544
rect 7208 20330 7236 20946
rect 7564 20936 7616 20942
rect 7564 20878 7616 20884
rect 7576 20806 7604 20878
rect 7564 20800 7616 20806
rect 7564 20742 7616 20748
rect 7196 20324 7248 20330
rect 7196 20266 7248 20272
rect 7012 19780 7064 19786
rect 7012 19722 7064 19728
rect 7564 19780 7616 19786
rect 7564 19722 7616 19728
rect 7024 19514 7052 19722
rect 7012 19508 7064 19514
rect 7012 19450 7064 19456
rect 6920 19440 6972 19446
rect 6920 19382 6972 19388
rect 7576 19378 7604 19722
rect 7656 19508 7708 19514
rect 7656 19450 7708 19456
rect 6184 19372 6236 19378
rect 6184 19314 6236 19320
rect 6276 19372 6328 19378
rect 6276 19314 6328 19320
rect 6460 19372 6512 19378
rect 6460 19314 6512 19320
rect 6736 19372 6788 19378
rect 6736 19314 6788 19320
rect 6828 19372 6880 19378
rect 6828 19314 6880 19320
rect 7564 19372 7616 19378
rect 7564 19314 7616 19320
rect 7104 19304 7156 19310
rect 7104 19246 7156 19252
rect 7012 19236 7064 19242
rect 7012 19178 7064 19184
rect 6000 18760 6052 18766
rect 6000 18702 6052 18708
rect 7024 18630 7052 19178
rect 7116 18630 7144 19246
rect 5724 18624 5776 18630
rect 5724 18566 5776 18572
rect 6644 18624 6696 18630
rect 6644 18566 6696 18572
rect 7012 18624 7064 18630
rect 7012 18566 7064 18572
rect 7104 18624 7156 18630
rect 7104 18566 7156 18572
rect 2872 18284 2924 18290
rect 2872 18226 2924 18232
rect 3056 18284 3108 18290
rect 3976 18284 4028 18290
rect 3056 18226 3108 18232
rect 3896 18244 3976 18272
rect 2884 17882 2912 18226
rect 2872 17876 2924 17882
rect 2872 17818 2924 17824
rect 3068 17678 3096 18226
rect 3896 18154 3924 18244
rect 3976 18226 4028 18232
rect 4896 18284 4948 18290
rect 4896 18226 4948 18232
rect 5172 18284 5224 18290
rect 5172 18226 5224 18232
rect 5264 18284 5316 18290
rect 5264 18226 5316 18232
rect 3884 18148 3936 18154
rect 3884 18090 3936 18096
rect 3608 18080 3660 18086
rect 3608 18022 3660 18028
rect 3620 17678 3648 18022
rect 3056 17672 3108 17678
rect 3056 17614 3108 17620
rect 3608 17672 3660 17678
rect 3608 17614 3660 17620
rect 3240 17128 3292 17134
rect 3240 17070 3292 17076
rect 3896 17082 3924 18090
rect 4160 18080 4212 18086
rect 4080 18040 4160 18068
rect 4080 17746 4108 18040
rect 4160 18022 4212 18028
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 5184 17746 5212 18226
rect 5276 17882 5304 18226
rect 5736 18222 5764 18566
rect 6000 18420 6052 18426
rect 6000 18362 6052 18368
rect 6184 18420 6236 18426
rect 6184 18362 6236 18368
rect 5724 18216 5776 18222
rect 5724 18158 5776 18164
rect 5540 18148 5592 18154
rect 5540 18090 5592 18096
rect 5552 17882 5580 18090
rect 5264 17876 5316 17882
rect 5264 17818 5316 17824
rect 5540 17876 5592 17882
rect 5540 17818 5592 17824
rect 4068 17740 4120 17746
rect 4068 17682 4120 17688
rect 5172 17740 5224 17746
rect 5172 17682 5224 17688
rect 4160 17672 4212 17678
rect 4160 17614 4212 17620
rect 4804 17672 4856 17678
rect 4804 17614 4856 17620
rect 4172 17338 4200 17614
rect 4712 17536 4764 17542
rect 4712 17478 4764 17484
rect 4160 17332 4212 17338
rect 4160 17274 4212 17280
rect 4068 17196 4120 17202
rect 4068 17138 4120 17144
rect 4080 17082 4108 17138
rect 2872 16992 2924 16998
rect 2872 16934 2924 16940
rect 2884 16726 2912 16934
rect 2872 16720 2924 16726
rect 2872 16662 2924 16668
rect 2964 16720 3016 16726
rect 2964 16662 3016 16668
rect 2976 16572 3004 16662
rect 2884 16544 3004 16572
rect 2780 15496 2832 15502
rect 2780 15438 2832 15444
rect 2504 15428 2556 15434
rect 2504 15370 2556 15376
rect 2516 15162 2544 15370
rect 2780 15360 2832 15366
rect 2780 15302 2832 15308
rect 2504 15156 2556 15162
rect 2504 15098 2556 15104
rect 2792 15094 2820 15302
rect 2780 15088 2832 15094
rect 2780 15030 2832 15036
rect 2792 14550 2820 15030
rect 2780 14544 2832 14550
rect 2780 14486 2832 14492
rect 2884 14346 2912 16544
rect 3252 15026 3280 17070
rect 3896 17054 4108 17082
rect 3608 16992 3660 16998
rect 3608 16934 3660 16940
rect 3620 16522 3648 16934
rect 3896 16590 3924 17054
rect 3976 16992 4028 16998
rect 3976 16934 4028 16940
rect 4068 16992 4120 16998
rect 4172 16980 4200 17274
rect 4724 17202 4752 17478
rect 4816 17338 4844 17614
rect 5736 17610 5764 18158
rect 6012 18154 6040 18362
rect 6000 18148 6052 18154
rect 6000 18090 6052 18096
rect 6092 18080 6144 18086
rect 6092 18022 6144 18028
rect 6104 17882 6132 18022
rect 6092 17876 6144 17882
rect 6092 17818 6144 17824
rect 6196 17678 6224 18362
rect 6656 18358 6684 18566
rect 6644 18352 6696 18358
rect 6644 18294 6696 18300
rect 7024 18222 7052 18566
rect 7012 18216 7064 18222
rect 7012 18158 7064 18164
rect 6644 18148 6696 18154
rect 6644 18090 6696 18096
rect 6552 18080 6604 18086
rect 6552 18022 6604 18028
rect 6184 17672 6236 17678
rect 6184 17614 6236 17620
rect 5264 17604 5316 17610
rect 5264 17546 5316 17552
rect 5724 17604 5776 17610
rect 5724 17546 5776 17552
rect 4874 17436 5182 17445
rect 4874 17434 4880 17436
rect 4936 17434 4960 17436
rect 5016 17434 5040 17436
rect 5096 17434 5120 17436
rect 5176 17434 5182 17436
rect 4936 17382 4938 17434
rect 5118 17382 5120 17434
rect 4874 17380 4880 17382
rect 4936 17380 4960 17382
rect 5016 17380 5040 17382
rect 5096 17380 5120 17382
rect 5176 17380 5182 17382
rect 4874 17371 5182 17380
rect 4804 17332 4856 17338
rect 4804 17274 4856 17280
rect 5276 17202 5304 17546
rect 4712 17196 4764 17202
rect 4712 17138 4764 17144
rect 4804 17196 4856 17202
rect 4804 17138 4856 17144
rect 5264 17196 5316 17202
rect 5264 17138 5316 17144
rect 5448 17196 5500 17202
rect 5448 17138 5500 17144
rect 4620 17128 4672 17134
rect 4620 17070 4672 17076
rect 4120 16952 4200 16980
rect 4068 16934 4120 16940
rect 3988 16590 4016 16934
rect 3884 16584 3936 16590
rect 3884 16526 3936 16532
rect 3976 16584 4028 16590
rect 3976 16526 4028 16532
rect 3608 16516 3660 16522
rect 3608 16458 3660 16464
rect 3988 16182 4016 16526
rect 3976 16176 4028 16182
rect 3976 16118 4028 16124
rect 3988 15502 4016 16118
rect 3976 15496 4028 15502
rect 3976 15438 4028 15444
rect 3884 15156 3936 15162
rect 3884 15098 3936 15104
rect 3896 15026 3924 15098
rect 4080 15026 4108 16934
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4436 16720 4488 16726
rect 4436 16662 4488 16668
rect 4448 16590 4476 16662
rect 4632 16590 4660 17070
rect 4816 16794 4844 17138
rect 4804 16788 4856 16794
rect 4804 16730 4856 16736
rect 4436 16584 4488 16590
rect 4436 16526 4488 16532
rect 4620 16584 4672 16590
rect 4620 16526 4672 16532
rect 4252 16448 4304 16454
rect 4252 16390 4304 16396
rect 4528 16448 4580 16454
rect 4528 16390 4580 16396
rect 4264 16114 4292 16390
rect 4540 16114 4568 16390
rect 4816 16182 4844 16730
rect 5276 16726 5304 17138
rect 5460 16998 5488 17138
rect 5736 17066 5764 17546
rect 6564 17202 6592 18022
rect 6656 17678 6684 18090
rect 6920 18080 6972 18086
rect 6920 18022 6972 18028
rect 6736 17876 6788 17882
rect 6736 17818 6788 17824
rect 6644 17672 6696 17678
rect 6644 17614 6696 17620
rect 6184 17196 6236 17202
rect 6184 17138 6236 17144
rect 6552 17196 6604 17202
rect 6552 17138 6604 17144
rect 5724 17060 5776 17066
rect 5724 17002 5776 17008
rect 5448 16992 5500 16998
rect 5448 16934 5500 16940
rect 5264 16720 5316 16726
rect 5264 16662 5316 16668
rect 4874 16348 5182 16357
rect 4874 16346 4880 16348
rect 4936 16346 4960 16348
rect 5016 16346 5040 16348
rect 5096 16346 5120 16348
rect 5176 16346 5182 16348
rect 4936 16294 4938 16346
rect 5118 16294 5120 16346
rect 4874 16292 4880 16294
rect 4936 16292 4960 16294
rect 5016 16292 5040 16294
rect 5096 16292 5120 16294
rect 5176 16292 5182 16294
rect 4874 16283 5182 16292
rect 4804 16176 4856 16182
rect 4804 16118 4856 16124
rect 4252 16108 4304 16114
rect 4252 16050 4304 16056
rect 4528 16108 4580 16114
rect 4528 16050 4580 16056
rect 4712 16108 4764 16114
rect 4712 16050 4764 16056
rect 4620 16040 4672 16046
rect 4620 15982 4672 15988
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4632 15570 4660 15982
rect 4620 15564 4672 15570
rect 4620 15506 4672 15512
rect 4724 15502 4752 16050
rect 4712 15496 4764 15502
rect 4712 15438 4764 15444
rect 4816 15366 4844 16118
rect 4804 15360 4856 15366
rect 4804 15302 4856 15308
rect 4816 15042 4844 15302
rect 4874 15260 5182 15269
rect 4874 15258 4880 15260
rect 4936 15258 4960 15260
rect 5016 15258 5040 15260
rect 5096 15258 5120 15260
rect 5176 15258 5182 15260
rect 4936 15206 4938 15258
rect 5118 15206 5120 15258
rect 4874 15204 4880 15206
rect 4936 15204 4960 15206
rect 5016 15204 5040 15206
rect 5096 15204 5120 15206
rect 5176 15204 5182 15206
rect 4874 15195 5182 15204
rect 3240 15020 3292 15026
rect 3240 14962 3292 14968
rect 3884 15020 3936 15026
rect 3884 14962 3936 14968
rect 4068 15020 4120 15026
rect 4068 14962 4120 14968
rect 4724 15014 4844 15042
rect 4988 15020 5040 15026
rect 3252 14482 3280 14962
rect 4724 14958 4752 15014
rect 4988 14962 5040 14968
rect 4712 14952 4764 14958
rect 4712 14894 4764 14900
rect 5000 14890 5028 14962
rect 4160 14884 4212 14890
rect 4080 14844 4160 14872
rect 3976 14816 4028 14822
rect 3976 14758 4028 14764
rect 3988 14550 4016 14758
rect 3700 14544 3752 14550
rect 3700 14486 3752 14492
rect 3976 14544 4028 14550
rect 3976 14486 4028 14492
rect 3240 14476 3292 14482
rect 3240 14418 3292 14424
rect 3608 14408 3660 14414
rect 3608 14350 3660 14356
rect 2872 14340 2924 14346
rect 2872 14282 2924 14288
rect 2412 13864 2464 13870
rect 2412 13806 2464 13812
rect 2136 12232 2188 12238
rect 2056 12192 2136 12220
rect 2136 12174 2188 12180
rect 2320 12232 2372 12238
rect 2320 12174 2372 12180
rect 1676 12096 1728 12102
rect 1676 12038 1728 12044
rect 1688 11762 1716 12038
rect 2424 11830 2452 13806
rect 2688 13252 2740 13258
rect 2688 13194 2740 13200
rect 2700 12850 2728 13194
rect 2688 12844 2740 12850
rect 2688 12786 2740 12792
rect 2700 12434 2728 12786
rect 2516 12406 2728 12434
rect 2516 12238 2544 12406
rect 2884 12238 2912 14282
rect 3620 13734 3648 14350
rect 3608 13728 3660 13734
rect 3608 13670 3660 13676
rect 3712 12374 3740 14486
rect 3884 14272 3936 14278
rect 3884 14214 3936 14220
rect 3792 12844 3844 12850
rect 3792 12786 3844 12792
rect 3804 12714 3832 12786
rect 3792 12708 3844 12714
rect 3792 12650 3844 12656
rect 3700 12368 3752 12374
rect 3700 12310 3752 12316
rect 3804 12238 3832 12650
rect 2504 12232 2556 12238
rect 2504 12174 2556 12180
rect 2872 12232 2924 12238
rect 2872 12174 2924 12180
rect 3792 12232 3844 12238
rect 3792 12174 3844 12180
rect 2516 11898 2544 12174
rect 3240 12096 3292 12102
rect 3240 12038 3292 12044
rect 2504 11892 2556 11898
rect 2504 11834 2556 11840
rect 2412 11824 2464 11830
rect 2412 11766 2464 11772
rect 1676 11756 1728 11762
rect 1676 11698 1728 11704
rect 3252 11694 3280 12038
rect 3896 11762 3924 14214
rect 3988 13818 4016 14486
rect 4080 14414 4108 14844
rect 4160 14826 4212 14832
rect 4988 14884 5040 14890
rect 4988 14826 5040 14832
rect 4620 14816 4672 14822
rect 4620 14758 4672 14764
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4068 14408 4120 14414
rect 4068 14350 4120 14356
rect 4080 14006 4108 14350
rect 4068 14000 4120 14006
rect 4068 13942 4120 13948
rect 4632 13870 4660 14758
rect 5000 14618 5028 14826
rect 4988 14612 5040 14618
rect 4988 14554 5040 14560
rect 5000 14414 5028 14554
rect 4988 14408 5040 14414
rect 4988 14350 5040 14356
rect 4804 14272 4856 14278
rect 4804 14214 4856 14220
rect 4712 14068 4764 14074
rect 4712 14010 4764 14016
rect 4620 13864 4672 13870
rect 3988 13790 4108 13818
rect 4620 13806 4672 13812
rect 3976 13728 4028 13734
rect 3976 13670 4028 13676
rect 3988 13190 4016 13670
rect 3976 13184 4028 13190
rect 3976 13126 4028 13132
rect 3988 12850 4016 13126
rect 3976 12844 4028 12850
rect 3976 12786 4028 12792
rect 4080 12782 4108 13790
rect 4632 13734 4660 13806
rect 4620 13728 4672 13734
rect 4620 13670 4672 13676
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4068 12776 4120 12782
rect 4068 12718 4120 12724
rect 4080 12306 4108 12718
rect 4620 12640 4672 12646
rect 4620 12582 4672 12588
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4252 12436 4304 12442
rect 4632 12434 4660 12582
rect 4304 12406 4660 12434
rect 4252 12378 4304 12384
rect 4068 12300 4120 12306
rect 4068 12242 4120 12248
rect 4632 12238 4660 12406
rect 4724 12306 4752 14010
rect 4816 14006 4844 14214
rect 4874 14172 5182 14181
rect 4874 14170 4880 14172
rect 4936 14170 4960 14172
rect 5016 14170 5040 14172
rect 5096 14170 5120 14172
rect 5176 14170 5182 14172
rect 4936 14118 4938 14170
rect 5118 14118 5120 14170
rect 4874 14116 4880 14118
rect 4936 14116 4960 14118
rect 5016 14116 5040 14118
rect 5096 14116 5120 14118
rect 5176 14116 5182 14118
rect 4874 14107 5182 14116
rect 4804 14000 4856 14006
rect 4804 13942 4856 13948
rect 5276 13530 5304 16662
rect 5460 16658 5488 16934
rect 5448 16652 5500 16658
rect 5448 16594 5500 16600
rect 5632 16448 5684 16454
rect 5632 16390 5684 16396
rect 5736 16402 5764 17002
rect 5816 16992 5868 16998
rect 5816 16934 5868 16940
rect 5828 16590 5856 16934
rect 5816 16584 5868 16590
rect 6000 16584 6052 16590
rect 5868 16544 5948 16572
rect 5816 16526 5868 16532
rect 5448 15972 5500 15978
rect 5448 15914 5500 15920
rect 5356 15360 5408 15366
rect 5356 15302 5408 15308
rect 5368 14618 5396 15302
rect 5356 14612 5408 14618
rect 5356 14554 5408 14560
rect 5460 14498 5488 15914
rect 5540 15360 5592 15366
rect 5540 15302 5592 15308
rect 5368 14470 5488 14498
rect 5264 13524 5316 13530
rect 5264 13466 5316 13472
rect 5264 13184 5316 13190
rect 5264 13126 5316 13132
rect 4874 13084 5182 13093
rect 4874 13082 4880 13084
rect 4936 13082 4960 13084
rect 5016 13082 5040 13084
rect 5096 13082 5120 13084
rect 5176 13082 5182 13084
rect 4936 13030 4938 13082
rect 5118 13030 5120 13082
rect 4874 13028 4880 13030
rect 4936 13028 4960 13030
rect 5016 13028 5040 13030
rect 5096 13028 5120 13030
rect 5176 13028 5182 13030
rect 4874 13019 5182 13028
rect 4712 12300 4764 12306
rect 4712 12242 4764 12248
rect 4620 12232 4672 12238
rect 4620 12174 4672 12180
rect 4160 12164 4212 12170
rect 4160 12106 4212 12112
rect 4172 11762 4200 12106
rect 3884 11756 3936 11762
rect 3884 11698 3936 11704
rect 4160 11756 4212 11762
rect 4160 11698 4212 11704
rect 3240 11688 3292 11694
rect 3240 11630 3292 11636
rect 3516 11620 3568 11626
rect 3516 11562 3568 11568
rect 3528 10810 3556 11562
rect 3516 10804 3568 10810
rect 3516 10746 3568 10752
rect 3424 9376 3476 9382
rect 3424 9318 3476 9324
rect 3436 9042 3464 9318
rect 3424 9036 3476 9042
rect 3424 8978 3476 8984
rect 3436 8430 3464 8978
rect 3528 8498 3556 10746
rect 3896 10742 3924 11698
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4632 11150 4660 12174
rect 4344 11144 4396 11150
rect 4344 11086 4396 11092
rect 4620 11144 4672 11150
rect 4724 11132 4752 12242
rect 4804 12096 4856 12102
rect 4804 12038 4856 12044
rect 4816 11778 4844 12038
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 4816 11750 4936 11778
rect 4804 11688 4856 11694
rect 4804 11630 4856 11636
rect 4816 11354 4844 11630
rect 4804 11348 4856 11354
rect 4804 11290 4856 11296
rect 4804 11144 4856 11150
rect 4724 11104 4804 11132
rect 4620 11086 4672 11092
rect 4804 11086 4856 11092
rect 3884 10736 3936 10742
rect 3884 10678 3936 10684
rect 3896 9586 3924 10678
rect 4160 10600 4212 10606
rect 4080 10548 4160 10554
rect 4080 10542 4212 10548
rect 4080 10526 4200 10542
rect 4356 10538 4384 11086
rect 4712 11008 4764 11014
rect 4712 10950 4764 10956
rect 4344 10532 4396 10538
rect 4080 10146 4108 10526
rect 4344 10474 4396 10480
rect 4620 10464 4672 10470
rect 4620 10406 4672 10412
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4080 10118 4200 10146
rect 3884 9580 3936 9586
rect 3884 9522 3936 9528
rect 4172 9466 4200 10118
rect 4632 9518 4660 10406
rect 4724 10062 4752 10950
rect 4816 10674 4844 11086
rect 4908 11014 4936 11750
rect 5172 11756 5224 11762
rect 5276 11744 5304 13126
rect 5368 12714 5396 14470
rect 5448 14272 5500 14278
rect 5448 14214 5500 14220
rect 5356 12708 5408 12714
rect 5356 12650 5408 12656
rect 5368 12374 5396 12650
rect 5356 12368 5408 12374
rect 5356 12310 5408 12316
rect 5356 12232 5408 12238
rect 5356 12174 5408 12180
rect 5368 11830 5396 12174
rect 5356 11824 5408 11830
rect 5356 11766 5408 11772
rect 5224 11716 5304 11744
rect 5172 11698 5224 11704
rect 5184 11150 5212 11698
rect 5172 11144 5224 11150
rect 5172 11086 5224 11092
rect 4896 11008 4948 11014
rect 5356 11008 5408 11014
rect 4896 10950 4948 10956
rect 5276 10968 5356 10996
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 5276 10674 5304 10968
rect 5356 10950 5408 10956
rect 4804 10668 4856 10674
rect 4804 10610 4856 10616
rect 5264 10668 5316 10674
rect 5264 10610 5316 10616
rect 4712 10056 4764 10062
rect 4712 9998 4764 10004
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 4712 9716 4764 9722
rect 4712 9658 4764 9664
rect 4724 9518 4752 9658
rect 4080 9438 4200 9466
rect 4620 9512 4672 9518
rect 4620 9454 4672 9460
rect 4712 9512 4764 9518
rect 4712 9454 4764 9460
rect 4988 9512 5040 9518
rect 4988 9454 5040 9460
rect 3792 9376 3844 9382
rect 3792 9318 3844 9324
rect 3804 8974 3832 9318
rect 4080 9160 4108 9438
rect 4712 9376 4764 9382
rect 4712 9318 4764 9324
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4080 9132 4200 9160
rect 3792 8968 3844 8974
rect 3792 8910 3844 8916
rect 3516 8492 3568 8498
rect 3516 8434 3568 8440
rect 3424 8424 3476 8430
rect 4172 8378 4200 9132
rect 4724 8498 4752 9318
rect 5000 9110 5028 9454
rect 5276 9110 5304 10610
rect 5356 10600 5408 10606
rect 5356 10542 5408 10548
rect 5368 9926 5396 10542
rect 5356 9920 5408 9926
rect 5356 9862 5408 9868
rect 5368 9722 5396 9862
rect 5356 9716 5408 9722
rect 5356 9658 5408 9664
rect 5356 9580 5408 9586
rect 5460 9568 5488 14214
rect 5552 13802 5580 15302
rect 5644 14278 5672 16390
rect 5736 16374 5856 16402
rect 5724 16108 5776 16114
rect 5724 16050 5776 16056
rect 5736 15434 5764 16050
rect 5724 15428 5776 15434
rect 5724 15370 5776 15376
rect 5736 15026 5764 15370
rect 5724 15020 5776 15026
rect 5724 14962 5776 14968
rect 5632 14272 5684 14278
rect 5632 14214 5684 14220
rect 5632 13864 5684 13870
rect 5828 13852 5856 16374
rect 5920 16114 5948 16544
rect 6000 16526 6052 16532
rect 5908 16108 5960 16114
rect 5908 16050 5960 16056
rect 5920 14822 5948 16050
rect 6012 15094 6040 16526
rect 6196 16522 6224 17138
rect 6748 17082 6776 17818
rect 6932 17678 6960 18022
rect 7116 17882 7144 18566
rect 7472 18284 7524 18290
rect 7472 18226 7524 18232
rect 7484 17882 7512 18226
rect 7104 17876 7156 17882
rect 7104 17818 7156 17824
rect 7472 17876 7524 17882
rect 7472 17818 7524 17824
rect 6920 17672 6972 17678
rect 6920 17614 6972 17620
rect 7576 17490 7604 19314
rect 7668 17678 7696 19450
rect 7760 19378 7788 21678
rect 7840 21626 7892 21632
rect 7944 21622 7972 25094
rect 8036 24818 8064 25638
rect 8220 25294 8248 25842
rect 8312 25770 8340 26998
rect 8392 26444 8444 26450
rect 8392 26386 8444 26392
rect 8404 25906 8432 26386
rect 8576 26376 8628 26382
rect 8576 26318 8628 26324
rect 8588 25906 8616 26318
rect 8772 25906 8800 27270
rect 8392 25900 8444 25906
rect 8392 25842 8444 25848
rect 8576 25900 8628 25906
rect 8576 25842 8628 25848
rect 8760 25900 8812 25906
rect 8760 25842 8812 25848
rect 8300 25764 8352 25770
rect 8300 25706 8352 25712
rect 8312 25362 8340 25706
rect 8300 25356 8352 25362
rect 8300 25298 8352 25304
rect 8208 25288 8260 25294
rect 8208 25230 8260 25236
rect 8300 25152 8352 25158
rect 8300 25094 8352 25100
rect 8484 25152 8536 25158
rect 8484 25094 8536 25100
rect 8116 24880 8168 24886
rect 8116 24822 8168 24828
rect 8024 24812 8076 24818
rect 8024 24754 8076 24760
rect 8128 24274 8156 24822
rect 8312 24410 8340 25094
rect 8392 24812 8444 24818
rect 8392 24754 8444 24760
rect 8404 24614 8432 24754
rect 8392 24608 8444 24614
rect 8392 24550 8444 24556
rect 8300 24404 8352 24410
rect 8300 24346 8352 24352
rect 8116 24268 8168 24274
rect 8116 24210 8168 24216
rect 8300 24200 8352 24206
rect 8404 24188 8432 24550
rect 8352 24160 8432 24188
rect 8300 24142 8352 24148
rect 8312 22964 8340 24142
rect 8392 23588 8444 23594
rect 8392 23530 8444 23536
rect 8404 23118 8432 23530
rect 8392 23112 8444 23118
rect 8392 23054 8444 23060
rect 8312 22936 8432 22964
rect 8300 22432 8352 22438
rect 8300 22374 8352 22380
rect 8312 22094 8340 22374
rect 8220 22066 8340 22094
rect 8220 22030 8248 22066
rect 8404 22030 8432 22936
rect 8496 22030 8524 25094
rect 8588 22778 8616 25842
rect 8772 25430 8800 25842
rect 8760 25424 8812 25430
rect 8760 25366 8812 25372
rect 8864 24206 8892 27406
rect 9312 26988 9364 26994
rect 9312 26930 9364 26936
rect 9496 26988 9548 26994
rect 9496 26930 9548 26936
rect 9324 25158 9352 26930
rect 9404 26920 9456 26926
rect 9404 26862 9456 26868
rect 9416 26450 9444 26862
rect 9404 26444 9456 26450
rect 9404 26386 9456 26392
rect 9416 26246 9444 26386
rect 9404 26240 9456 26246
rect 9404 26182 9456 26188
rect 9416 25906 9444 26182
rect 9508 26042 9536 26930
rect 10600 26784 10652 26790
rect 10600 26726 10652 26732
rect 10612 26382 10640 26726
rect 10888 26382 10916 27474
rect 10600 26376 10652 26382
rect 10600 26318 10652 26324
rect 10876 26376 10928 26382
rect 10876 26318 10928 26324
rect 9496 26036 9548 26042
rect 9496 25978 9548 25984
rect 10980 25906 11008 27882
rect 11336 27872 11388 27878
rect 11336 27814 11388 27820
rect 11348 27470 11376 27814
rect 12544 27674 12572 28494
rect 13176 28484 13228 28490
rect 13176 28426 13228 28432
rect 16856 28484 16908 28490
rect 16856 28426 16908 28432
rect 12716 28416 12768 28422
rect 12716 28358 12768 28364
rect 12728 28082 12756 28358
rect 12716 28076 12768 28082
rect 12716 28018 12768 28024
rect 12624 27940 12676 27946
rect 12624 27882 12676 27888
rect 12532 27668 12584 27674
rect 12532 27610 12584 27616
rect 11336 27464 11388 27470
rect 11336 27406 11388 27412
rect 12636 27334 12664 27882
rect 12624 27328 12676 27334
rect 12624 27270 12676 27276
rect 12440 26988 12492 26994
rect 12440 26930 12492 26936
rect 11612 26376 11664 26382
rect 11612 26318 11664 26324
rect 11244 26308 11296 26314
rect 11244 26250 11296 26256
rect 11256 26042 11284 26250
rect 11244 26036 11296 26042
rect 11244 25978 11296 25984
rect 9404 25900 9456 25906
rect 9404 25842 9456 25848
rect 9588 25900 9640 25906
rect 9588 25842 9640 25848
rect 10968 25900 11020 25906
rect 10968 25842 11020 25848
rect 9600 25362 9628 25842
rect 11624 25362 11652 26318
rect 12452 26246 12480 26930
rect 12636 26790 12664 27270
rect 12992 26920 13044 26926
rect 12992 26862 13044 26868
rect 12624 26784 12676 26790
rect 12624 26726 12676 26732
rect 12716 26512 12768 26518
rect 12716 26454 12768 26460
rect 12440 26240 12492 26246
rect 12440 26182 12492 26188
rect 12728 25906 12756 26454
rect 13004 26314 13032 26862
rect 13188 26790 13216 28426
rect 16580 28212 16632 28218
rect 16580 28154 16632 28160
rect 14096 28144 14148 28150
rect 14096 28086 14148 28092
rect 14004 27872 14056 27878
rect 14004 27814 14056 27820
rect 14016 27538 14044 27814
rect 14004 27532 14056 27538
rect 14004 27474 14056 27480
rect 13636 27464 13688 27470
rect 13636 27406 13688 27412
rect 13360 27396 13412 27402
rect 13360 27338 13412 27344
rect 13544 27396 13596 27402
rect 13544 27338 13596 27344
rect 13176 26784 13228 26790
rect 13176 26726 13228 26732
rect 13188 26330 13216 26726
rect 13268 26376 13320 26382
rect 13188 26324 13268 26330
rect 13188 26318 13320 26324
rect 12992 26308 13044 26314
rect 12992 26250 13044 26256
rect 13188 26302 13308 26318
rect 12716 25900 12768 25906
rect 12716 25842 12768 25848
rect 13004 25702 13032 26250
rect 13188 26234 13216 26302
rect 13372 26296 13400 27338
rect 13556 27062 13584 27338
rect 13544 27056 13596 27062
rect 13544 26998 13596 27004
rect 13648 26994 13676 27406
rect 14016 27146 14044 27474
rect 13924 27130 14044 27146
rect 13912 27124 14044 27130
rect 13964 27118 14044 27124
rect 13912 27066 13964 27072
rect 13820 27056 13872 27062
rect 13820 26998 13872 27004
rect 13636 26988 13688 26994
rect 13636 26930 13688 26936
rect 13648 26790 13676 26930
rect 13636 26784 13688 26790
rect 13636 26726 13688 26732
rect 13544 26308 13596 26314
rect 13372 26268 13544 26296
rect 13096 26206 13216 26234
rect 13268 26240 13320 26246
rect 13096 26042 13124 26206
rect 13268 26182 13320 26188
rect 13084 26036 13136 26042
rect 13084 25978 13136 25984
rect 13280 25974 13308 26182
rect 13268 25968 13320 25974
rect 13268 25910 13320 25916
rect 13084 25832 13136 25838
rect 13084 25774 13136 25780
rect 12992 25696 13044 25702
rect 12992 25638 13044 25644
rect 9588 25356 9640 25362
rect 9588 25298 9640 25304
rect 11612 25356 11664 25362
rect 11612 25298 11664 25304
rect 10048 25288 10100 25294
rect 10048 25230 10100 25236
rect 9312 25152 9364 25158
rect 9312 25094 9364 25100
rect 9956 24812 10008 24818
rect 9956 24754 10008 24760
rect 8852 24200 8904 24206
rect 8852 24142 8904 24148
rect 8944 24132 8996 24138
rect 8944 24074 8996 24080
rect 8668 23112 8720 23118
rect 8668 23054 8720 23060
rect 8576 22772 8628 22778
rect 8576 22714 8628 22720
rect 8208 22024 8260 22030
rect 8208 21966 8260 21972
rect 8392 22024 8444 22030
rect 8392 21966 8444 21972
rect 8484 22024 8536 22030
rect 8484 21966 8536 21972
rect 7932 21616 7984 21622
rect 7932 21558 7984 21564
rect 8024 21548 8076 21554
rect 8024 21490 8076 21496
rect 7840 21344 7892 21350
rect 7840 21286 7892 21292
rect 7852 20942 7880 21286
rect 8036 21010 8064 21490
rect 8024 21004 8076 21010
rect 8024 20946 8076 20952
rect 7840 20936 7892 20942
rect 7840 20878 7892 20884
rect 8024 20528 8076 20534
rect 8024 20470 8076 20476
rect 8036 19990 8064 20470
rect 8116 20324 8168 20330
rect 8116 20266 8168 20272
rect 8024 19984 8076 19990
rect 8024 19926 8076 19932
rect 8128 19922 8156 20266
rect 8116 19916 8168 19922
rect 8116 19858 8168 19864
rect 8220 19854 8248 21966
rect 8680 21146 8708 23054
rect 8956 21894 8984 24074
rect 9404 24064 9456 24070
rect 9404 24006 9456 24012
rect 9312 23112 9364 23118
rect 9312 23054 9364 23060
rect 9036 22976 9088 22982
rect 9036 22918 9088 22924
rect 9220 22976 9272 22982
rect 9220 22918 9272 22924
rect 9048 22438 9076 22918
rect 9232 22506 9260 22918
rect 9220 22500 9272 22506
rect 9220 22442 9272 22448
rect 9036 22432 9088 22438
rect 9036 22374 9088 22380
rect 8944 21888 8996 21894
rect 8944 21830 8996 21836
rect 8956 21418 8984 21830
rect 8944 21412 8996 21418
rect 8944 21354 8996 21360
rect 8668 21140 8720 21146
rect 8668 21082 8720 21088
rect 8208 19848 8260 19854
rect 8208 19790 8260 19796
rect 7748 19372 7800 19378
rect 7800 19332 8340 19360
rect 7748 19314 7800 19320
rect 8312 18698 8340 19332
rect 8680 18970 8708 21082
rect 9324 20942 9352 23054
rect 9416 22642 9444 24006
rect 9968 23798 9996 24754
rect 10060 24750 10088 25230
rect 10968 25220 11020 25226
rect 10968 25162 11020 25168
rect 10508 25152 10560 25158
rect 10508 25094 10560 25100
rect 10520 24818 10548 25094
rect 10324 24812 10376 24818
rect 10324 24754 10376 24760
rect 10508 24812 10560 24818
rect 10508 24754 10560 24760
rect 10048 24744 10100 24750
rect 10048 24686 10100 24692
rect 10060 24070 10088 24686
rect 10048 24064 10100 24070
rect 10048 24006 10100 24012
rect 9956 23792 10008 23798
rect 9956 23734 10008 23740
rect 9772 23112 9824 23118
rect 9772 23054 9824 23060
rect 9404 22636 9456 22642
rect 9404 22578 9456 22584
rect 9416 21010 9444 22578
rect 9784 22166 9812 23054
rect 9968 22642 9996 23734
rect 10336 23730 10364 24754
rect 10784 24744 10836 24750
rect 10784 24686 10836 24692
rect 10416 24608 10468 24614
rect 10416 24550 10468 24556
rect 10428 23866 10456 24550
rect 10416 23860 10468 23866
rect 10416 23802 10468 23808
rect 10324 23724 10376 23730
rect 10324 23666 10376 23672
rect 10140 23180 10192 23186
rect 10140 23122 10192 23128
rect 9956 22636 10008 22642
rect 9956 22578 10008 22584
rect 9772 22160 9824 22166
rect 9772 22102 9824 22108
rect 9968 22030 9996 22578
rect 9956 22024 10008 22030
rect 9956 21966 10008 21972
rect 9772 21956 9824 21962
rect 9772 21898 9824 21904
rect 9404 21004 9456 21010
rect 9404 20946 9456 20952
rect 9312 20936 9364 20942
rect 9312 20878 9364 20884
rect 9036 20800 9088 20806
rect 9036 20742 9088 20748
rect 9048 20398 9076 20742
rect 9036 20392 9088 20398
rect 9036 20334 9088 20340
rect 9324 19990 9352 20878
rect 9680 20868 9732 20874
rect 9680 20810 9732 20816
rect 9692 20602 9720 20810
rect 9680 20596 9732 20602
rect 9680 20538 9732 20544
rect 9312 19984 9364 19990
rect 9312 19926 9364 19932
rect 9324 19514 9352 19926
rect 9784 19854 9812 21898
rect 10152 21894 10180 23122
rect 10336 22710 10364 23666
rect 10428 23662 10456 23802
rect 10416 23656 10468 23662
rect 10416 23598 10468 23604
rect 10796 23526 10824 24686
rect 10980 23730 11008 25162
rect 11624 24750 11652 25298
rect 12440 25220 12492 25226
rect 12440 25162 12492 25168
rect 11612 24744 11664 24750
rect 11612 24686 11664 24692
rect 12348 24744 12400 24750
rect 12348 24686 12400 24692
rect 12072 24608 12124 24614
rect 12072 24550 12124 24556
rect 12084 24206 12112 24550
rect 12360 24274 12388 24686
rect 12452 24410 12480 25162
rect 12624 25152 12676 25158
rect 12624 25094 12676 25100
rect 12440 24404 12492 24410
rect 12440 24346 12492 24352
rect 12348 24268 12400 24274
rect 12348 24210 12400 24216
rect 12636 24206 12664 25094
rect 13096 24206 13124 25774
rect 13176 25696 13228 25702
rect 13176 25638 13228 25644
rect 12072 24200 12124 24206
rect 12072 24142 12124 24148
rect 12624 24200 12676 24206
rect 12624 24142 12676 24148
rect 12808 24200 12860 24206
rect 12808 24142 12860 24148
rect 12992 24200 13044 24206
rect 12992 24142 13044 24148
rect 13084 24200 13136 24206
rect 13084 24142 13136 24148
rect 12072 24064 12124 24070
rect 12072 24006 12124 24012
rect 12084 23730 12112 24006
rect 10968 23724 11020 23730
rect 10968 23666 11020 23672
rect 12072 23724 12124 23730
rect 12072 23666 12124 23672
rect 10784 23520 10836 23526
rect 10784 23462 10836 23468
rect 10784 23112 10836 23118
rect 10784 23054 10836 23060
rect 10796 22778 10824 23054
rect 12084 22778 12112 23666
rect 12440 23656 12492 23662
rect 12440 23598 12492 23604
rect 10784 22772 10836 22778
rect 10784 22714 10836 22720
rect 12072 22772 12124 22778
rect 12072 22714 12124 22720
rect 10324 22704 10376 22710
rect 10324 22646 10376 22652
rect 10416 22500 10468 22506
rect 10416 22442 10468 22448
rect 10428 21962 10456 22442
rect 10796 22438 10824 22714
rect 10968 22704 11020 22710
rect 11020 22652 11284 22658
rect 10968 22646 11284 22652
rect 10980 22642 11284 22646
rect 10980 22636 11296 22642
rect 10980 22630 11244 22636
rect 11244 22578 11296 22584
rect 10968 22568 11020 22574
rect 10968 22510 11020 22516
rect 10784 22432 10836 22438
rect 10784 22374 10836 22380
rect 10796 22030 10824 22374
rect 10980 22166 11008 22510
rect 12072 22432 12124 22438
rect 12072 22374 12124 22380
rect 12164 22432 12216 22438
rect 12164 22374 12216 22380
rect 12084 22166 12112 22374
rect 10968 22160 11020 22166
rect 10968 22102 11020 22108
rect 12072 22160 12124 22166
rect 12072 22102 12124 22108
rect 10784 22024 10836 22030
rect 10784 21966 10836 21972
rect 10416 21956 10468 21962
rect 10416 21898 10468 21904
rect 10140 21888 10192 21894
rect 10140 21830 10192 21836
rect 10152 20806 10180 21830
rect 10980 21146 11008 22102
rect 12176 22094 12204 22374
rect 12176 22066 12388 22094
rect 12176 22030 12204 22066
rect 12164 22024 12216 22030
rect 12164 21966 12216 21972
rect 12360 21962 12388 22066
rect 11704 21956 11756 21962
rect 12072 21956 12124 21962
rect 11756 21916 12072 21944
rect 11704 21898 11756 21904
rect 12072 21898 12124 21904
rect 12348 21956 12400 21962
rect 12348 21898 12400 21904
rect 11520 21888 11572 21894
rect 11520 21830 11572 21836
rect 11532 21554 11560 21830
rect 12162 21720 12218 21729
rect 12162 21655 12218 21664
rect 12176 21622 12204 21655
rect 12164 21616 12216 21622
rect 12164 21558 12216 21564
rect 12254 21584 12310 21593
rect 11520 21548 11572 21554
rect 12254 21519 12256 21528
rect 11520 21490 11572 21496
rect 12308 21519 12310 21528
rect 12256 21490 12308 21496
rect 11888 21412 11940 21418
rect 11888 21354 11940 21360
rect 10600 21140 10652 21146
rect 10600 21082 10652 21088
rect 10968 21140 11020 21146
rect 10968 21082 11020 21088
rect 10140 20800 10192 20806
rect 10140 20742 10192 20748
rect 10612 20466 10640 21082
rect 10784 20800 10836 20806
rect 10784 20742 10836 20748
rect 10796 20534 10824 20742
rect 10784 20528 10836 20534
rect 10782 20496 10784 20505
rect 10836 20496 10838 20505
rect 10600 20460 10652 20466
rect 10782 20431 10838 20440
rect 11428 20460 11480 20466
rect 10600 20402 10652 20408
rect 11428 20402 11480 20408
rect 10324 20392 10376 20398
rect 10324 20334 10376 20340
rect 10336 19854 10364 20334
rect 10784 20256 10836 20262
rect 10784 20198 10836 20204
rect 9772 19848 9824 19854
rect 10324 19848 10376 19854
rect 9824 19808 9904 19836
rect 9772 19790 9824 19796
rect 9680 19712 9732 19718
rect 9680 19654 9732 19660
rect 9312 19508 9364 19514
rect 9312 19450 9364 19456
rect 8944 19168 8996 19174
rect 8944 19110 8996 19116
rect 9496 19168 9548 19174
rect 9496 19110 9548 19116
rect 8668 18964 8720 18970
rect 8668 18906 8720 18912
rect 8300 18692 8352 18698
rect 8300 18634 8352 18640
rect 8956 18630 8984 19110
rect 8944 18624 8996 18630
rect 8944 18566 8996 18572
rect 9036 18624 9088 18630
rect 9036 18566 9088 18572
rect 8668 18080 8720 18086
rect 8668 18022 8720 18028
rect 8680 17746 8708 18022
rect 8668 17740 8720 17746
rect 8668 17682 8720 17688
rect 8956 17678 8984 18566
rect 7656 17672 7708 17678
rect 7656 17614 7708 17620
rect 8944 17672 8996 17678
rect 8944 17614 8996 17620
rect 7840 17604 7892 17610
rect 7840 17546 7892 17552
rect 7852 17490 7880 17546
rect 7576 17462 7880 17490
rect 6564 17066 6776 17082
rect 6552 17060 6776 17066
rect 6604 17054 6776 17060
rect 6552 17002 6604 17008
rect 6368 16992 6420 16998
rect 6368 16934 6420 16940
rect 6460 16992 6512 16998
rect 6460 16934 6512 16940
rect 6380 16794 6408 16934
rect 6368 16788 6420 16794
rect 6368 16730 6420 16736
rect 6472 16590 6500 16934
rect 6564 16590 6592 17002
rect 7656 16992 7708 16998
rect 7656 16934 7708 16940
rect 7668 16590 7696 16934
rect 6460 16584 6512 16590
rect 6460 16526 6512 16532
rect 6552 16584 6604 16590
rect 6552 16526 6604 16532
rect 6828 16584 6880 16590
rect 6828 16526 6880 16532
rect 7656 16584 7708 16590
rect 7656 16526 7708 16532
rect 6184 16516 6236 16522
rect 6184 16458 6236 16464
rect 6184 15904 6236 15910
rect 6184 15846 6236 15852
rect 6196 15570 6224 15846
rect 6184 15564 6236 15570
rect 6184 15506 6236 15512
rect 6564 15502 6592 16526
rect 6840 16114 6868 16526
rect 7852 16250 7880 17462
rect 8116 17332 8168 17338
rect 8116 17274 8168 17280
rect 8128 17202 8156 17274
rect 8116 17196 8168 17202
rect 8116 17138 8168 17144
rect 8484 17196 8536 17202
rect 8484 17138 8536 17144
rect 7840 16244 7892 16250
rect 7840 16186 7892 16192
rect 8128 16114 8156 17138
rect 8496 16810 8524 17138
rect 8496 16782 8616 16810
rect 8588 16726 8616 16782
rect 8576 16720 8628 16726
rect 8576 16662 8628 16668
rect 6828 16108 6880 16114
rect 6828 16050 6880 16056
rect 7656 16108 7708 16114
rect 7656 16050 7708 16056
rect 7748 16108 7800 16114
rect 8116 16108 8168 16114
rect 7748 16050 7800 16056
rect 8036 16068 8116 16096
rect 7196 15904 7248 15910
rect 7196 15846 7248 15852
rect 6092 15496 6144 15502
rect 6092 15438 6144 15444
rect 6552 15496 6604 15502
rect 6552 15438 6604 15444
rect 6000 15088 6052 15094
rect 6000 15030 6052 15036
rect 6104 15026 6132 15438
rect 7208 15026 7236 15846
rect 7668 15638 7696 16050
rect 7760 15706 7788 16050
rect 7748 15700 7800 15706
rect 7748 15642 7800 15648
rect 7656 15632 7708 15638
rect 7656 15574 7708 15580
rect 7656 15428 7708 15434
rect 7656 15370 7708 15376
rect 7668 15094 7696 15370
rect 7656 15088 7708 15094
rect 7656 15030 7708 15036
rect 6092 15020 6144 15026
rect 6092 14962 6144 14968
rect 7196 15020 7248 15026
rect 7196 14962 7248 14968
rect 7288 15020 7340 15026
rect 7288 14962 7340 14968
rect 5908 14816 5960 14822
rect 5908 14758 5960 14764
rect 6368 14816 6420 14822
rect 6368 14758 6420 14764
rect 6552 14816 6604 14822
rect 6552 14758 6604 14764
rect 6380 14074 6408 14758
rect 5908 14068 5960 14074
rect 5908 14010 5960 14016
rect 6368 14068 6420 14074
rect 6368 14010 6420 14016
rect 5684 13824 5856 13852
rect 5632 13806 5684 13812
rect 5540 13796 5592 13802
rect 5540 13738 5592 13744
rect 5552 13462 5580 13738
rect 5540 13456 5592 13462
rect 5540 13398 5592 13404
rect 5552 12850 5580 13398
rect 5644 13326 5672 13806
rect 5632 13320 5684 13326
rect 5632 13262 5684 13268
rect 5540 12844 5592 12850
rect 5540 12786 5592 12792
rect 5540 11756 5592 11762
rect 5540 11698 5592 11704
rect 5724 11756 5776 11762
rect 5724 11698 5776 11704
rect 5552 11150 5580 11698
rect 5736 11150 5764 11698
rect 5540 11144 5592 11150
rect 5540 11086 5592 11092
rect 5724 11144 5776 11150
rect 5724 11086 5776 11092
rect 5540 10124 5592 10130
rect 5540 10066 5592 10072
rect 5552 9674 5580 10066
rect 5920 10062 5948 14010
rect 6092 13864 6144 13870
rect 6092 13806 6144 13812
rect 5908 10056 5960 10062
rect 5908 9998 5960 10004
rect 5816 9920 5868 9926
rect 5816 9862 5868 9868
rect 5552 9646 5672 9674
rect 5644 9586 5672 9646
rect 5408 9540 5488 9568
rect 5356 9522 5408 9528
rect 4988 9104 5040 9110
rect 4988 9046 5040 9052
rect 5264 9104 5316 9110
rect 5264 9046 5316 9052
rect 5460 8974 5488 9540
rect 5540 9580 5592 9586
rect 5540 9522 5592 9528
rect 5632 9580 5684 9586
rect 5632 9522 5684 9528
rect 5552 9489 5580 9522
rect 5538 9480 5594 9489
rect 5828 9450 5856 9862
rect 5538 9415 5594 9424
rect 5816 9444 5868 9450
rect 5816 9386 5868 9392
rect 5540 9376 5592 9382
rect 5540 9318 5592 9324
rect 5552 8974 5580 9318
rect 5448 8968 5500 8974
rect 5448 8910 5500 8916
rect 5540 8968 5592 8974
rect 5540 8910 5592 8916
rect 4804 8832 4856 8838
rect 4804 8774 4856 8780
rect 4620 8492 4672 8498
rect 4620 8434 4672 8440
rect 4712 8492 4764 8498
rect 4712 8434 4764 8440
rect 3424 8366 3476 8372
rect 4080 8350 4200 8378
rect 4080 8004 4108 8350
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4080 7976 4200 8004
rect 4172 7478 4200 7976
rect 4632 7954 4660 8434
rect 4712 8356 4764 8362
rect 4712 8298 4764 8304
rect 4724 8022 4752 8298
rect 4712 8016 4764 8022
rect 4712 7958 4764 7964
rect 4620 7948 4672 7954
rect 4620 7890 4672 7896
rect 4436 7744 4488 7750
rect 4436 7686 4488 7692
rect 4160 7472 4212 7478
rect 4160 7414 4212 7420
rect 4448 7410 4476 7686
rect 4632 7546 4660 7890
rect 4620 7540 4672 7546
rect 4620 7482 4672 7488
rect 4816 7426 4844 8774
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 4896 8628 4948 8634
rect 4896 8570 4948 8576
rect 4908 7818 4936 8570
rect 5080 8492 5132 8498
rect 5080 8434 5132 8440
rect 4988 8424 5040 8430
rect 4988 8366 5040 8372
rect 4896 7812 4948 7818
rect 4896 7754 4948 7760
rect 5000 7750 5028 8366
rect 5092 7750 5120 8434
rect 5264 8288 5316 8294
rect 5264 8230 5316 8236
rect 5276 7886 5304 8230
rect 5448 8016 5500 8022
rect 5448 7958 5500 7964
rect 5264 7880 5316 7886
rect 5460 7857 5488 7958
rect 5264 7822 5316 7828
rect 5446 7848 5502 7857
rect 5356 7812 5408 7818
rect 5446 7783 5502 7792
rect 5632 7812 5684 7818
rect 5356 7754 5408 7760
rect 5632 7754 5684 7760
rect 4988 7744 5040 7750
rect 4988 7686 5040 7692
rect 5080 7744 5132 7750
rect 5080 7686 5132 7692
rect 5264 7744 5316 7750
rect 5264 7686 5316 7692
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 5276 7546 5304 7686
rect 5264 7540 5316 7546
rect 5264 7482 5316 7488
rect 4632 7410 4844 7426
rect 4436 7404 4488 7410
rect 4436 7346 4488 7352
rect 4620 7404 4844 7410
rect 4672 7398 4844 7404
rect 4620 7346 4672 7352
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4632 4622 4660 7346
rect 4712 7268 4764 7274
rect 4712 7210 4764 7216
rect 4724 5234 4752 7210
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 5276 6338 5304 7482
rect 5368 7274 5396 7754
rect 5356 7268 5408 7274
rect 5356 7210 5408 7216
rect 5644 6458 5672 7754
rect 5724 7404 5776 7410
rect 5724 7346 5776 7352
rect 5632 6452 5684 6458
rect 5632 6394 5684 6400
rect 5276 6322 5488 6338
rect 5736 6322 5764 7346
rect 5828 7342 5856 9386
rect 5908 8832 5960 8838
rect 5908 8774 5960 8780
rect 5816 7336 5868 7342
rect 5816 7278 5868 7284
rect 5264 6316 5488 6322
rect 5316 6310 5488 6316
rect 5460 6304 5488 6310
rect 5540 6316 5592 6322
rect 5460 6276 5540 6304
rect 5264 6258 5316 6264
rect 5540 6258 5592 6264
rect 5724 6316 5776 6322
rect 5724 6258 5776 6264
rect 5724 6180 5776 6186
rect 5724 6122 5776 6128
rect 4804 6112 4856 6118
rect 4804 6054 4856 6060
rect 4816 5302 4844 6054
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 4804 5296 4856 5302
rect 4804 5238 4856 5244
rect 4712 5228 4764 5234
rect 4712 5170 4764 5176
rect 4816 5098 4844 5238
rect 5736 5234 5764 6122
rect 5920 5710 5948 8774
rect 6000 6248 6052 6254
rect 6000 6190 6052 6196
rect 5908 5704 5960 5710
rect 5908 5646 5960 5652
rect 5920 5234 5948 5646
rect 6012 5574 6040 6190
rect 6104 5710 6132 13806
rect 6368 12776 6420 12782
rect 6368 12718 6420 12724
rect 6184 11552 6236 11558
rect 6184 11494 6236 11500
rect 6196 9994 6224 11494
rect 6276 10600 6328 10606
rect 6276 10542 6328 10548
rect 6288 10266 6316 10542
rect 6276 10260 6328 10266
rect 6276 10202 6328 10208
rect 6184 9988 6236 9994
rect 6184 9930 6236 9936
rect 6276 7268 6328 7274
rect 6276 7210 6328 7216
rect 6380 7256 6408 12718
rect 6564 11744 6592 14758
rect 7208 14550 7236 14962
rect 7196 14544 7248 14550
rect 7196 14486 7248 14492
rect 7300 14414 7328 14962
rect 7380 14476 7432 14482
rect 7380 14418 7432 14424
rect 7288 14408 7340 14414
rect 7288 14350 7340 14356
rect 6920 13864 6972 13870
rect 6920 13806 6972 13812
rect 6932 12782 6960 13806
rect 7196 13796 7248 13802
rect 7196 13738 7248 13744
rect 7208 13462 7236 13738
rect 7196 13456 7248 13462
rect 7196 13398 7248 13404
rect 7288 13184 7340 13190
rect 7288 13126 7340 13132
rect 6920 12776 6972 12782
rect 6920 12718 6972 12724
rect 6736 12436 6788 12442
rect 6736 12378 6788 12384
rect 6644 11756 6696 11762
rect 6564 11716 6644 11744
rect 6644 11698 6696 11704
rect 6552 11620 6604 11626
rect 6552 11562 6604 11568
rect 6564 11082 6592 11562
rect 6552 11076 6604 11082
rect 6552 11018 6604 11024
rect 6564 10554 6592 11018
rect 6656 10674 6684 11698
rect 6644 10668 6696 10674
rect 6644 10610 6696 10616
rect 6564 10526 6684 10554
rect 6656 9994 6684 10526
rect 6552 9988 6604 9994
rect 6552 9930 6604 9936
rect 6644 9988 6696 9994
rect 6644 9930 6696 9936
rect 6564 9654 6592 9930
rect 6552 9648 6604 9654
rect 6552 9590 6604 9596
rect 6564 9489 6592 9590
rect 6656 9586 6684 9930
rect 6644 9580 6696 9586
rect 6644 9522 6696 9528
rect 6550 9480 6606 9489
rect 6550 9415 6606 9424
rect 6552 9376 6604 9382
rect 6552 9318 6604 9324
rect 6564 9042 6592 9318
rect 6552 9036 6604 9042
rect 6552 8978 6604 8984
rect 6748 8974 6776 12378
rect 6828 12096 6880 12102
rect 6828 12038 6880 12044
rect 6840 11694 6868 12038
rect 6932 11762 6960 12718
rect 7300 12306 7328 13126
rect 7288 12300 7340 12306
rect 7288 12242 7340 12248
rect 7392 12238 7420 14418
rect 7668 14074 7696 15030
rect 7760 14482 7788 15642
rect 8036 15502 8064 16068
rect 8116 16050 8168 16056
rect 8392 16108 8444 16114
rect 8392 16050 8444 16056
rect 8484 16108 8536 16114
rect 8484 16050 8536 16056
rect 8116 15904 8168 15910
rect 8116 15846 8168 15852
rect 8300 15904 8352 15910
rect 8300 15846 8352 15852
rect 8128 15570 8156 15846
rect 8116 15564 8168 15570
rect 8116 15506 8168 15512
rect 8024 15496 8076 15502
rect 8024 15438 8076 15444
rect 7748 14476 7800 14482
rect 7748 14418 7800 14424
rect 7656 14068 7708 14074
rect 7656 14010 7708 14016
rect 7656 13932 7708 13938
rect 7760 13920 7788 14418
rect 8208 14272 8260 14278
rect 8208 14214 8260 14220
rect 8312 14226 8340 15846
rect 8404 15502 8432 16050
rect 8496 15502 8524 16050
rect 8588 16046 8616 16662
rect 8852 16584 8904 16590
rect 8852 16526 8904 16532
rect 8864 16046 8892 16526
rect 8956 16454 8984 17614
rect 9048 17542 9076 18566
rect 9312 18284 9364 18290
rect 9312 18226 9364 18232
rect 9324 17678 9352 18226
rect 9508 18222 9536 19110
rect 9692 18766 9720 19654
rect 9772 19372 9824 19378
rect 9772 19314 9824 19320
rect 9680 18760 9732 18766
rect 9680 18702 9732 18708
rect 9680 18624 9732 18630
rect 9680 18566 9732 18572
rect 9496 18216 9548 18222
rect 9496 18158 9548 18164
rect 9588 17740 9640 17746
rect 9588 17682 9640 17688
rect 9312 17672 9364 17678
rect 9312 17614 9364 17620
rect 9036 17536 9088 17542
rect 9036 17478 9088 17484
rect 9048 17338 9076 17478
rect 9036 17332 9088 17338
rect 9036 17274 9088 17280
rect 9324 17270 9352 17614
rect 9496 17604 9548 17610
rect 9496 17546 9548 17552
rect 9404 17536 9456 17542
rect 9404 17478 9456 17484
rect 9312 17264 9364 17270
rect 9312 17206 9364 17212
rect 9416 17202 9444 17478
rect 9404 17196 9456 17202
rect 9404 17138 9456 17144
rect 9416 16590 9444 17138
rect 9508 16726 9536 17546
rect 9600 17134 9628 17682
rect 9692 17678 9720 18566
rect 9784 18426 9812 19314
rect 9876 18970 9904 19808
rect 10324 19790 10376 19796
rect 10140 19712 10192 19718
rect 10140 19654 10192 19660
rect 10048 19304 10100 19310
rect 10048 19246 10100 19252
rect 9864 18964 9916 18970
rect 9864 18906 9916 18912
rect 10060 18766 10088 19246
rect 10152 18902 10180 19654
rect 10336 19446 10364 19790
rect 10796 19514 10824 20198
rect 11440 19514 11468 20402
rect 11900 20058 11928 21354
rect 12360 20806 12388 21898
rect 12452 21536 12480 23598
rect 12820 23322 12848 24142
rect 12900 24064 12952 24070
rect 12900 24006 12952 24012
rect 12912 23798 12940 24006
rect 12900 23792 12952 23798
rect 12900 23734 12952 23740
rect 13004 23322 13032 24142
rect 13096 23730 13124 24142
rect 13188 24138 13216 25638
rect 13280 25498 13308 25910
rect 13372 25838 13400 26268
rect 13544 26250 13596 26256
rect 13452 26036 13504 26042
rect 13452 25978 13504 25984
rect 13360 25832 13412 25838
rect 13360 25774 13412 25780
rect 13464 25702 13492 25978
rect 13648 25906 13676 26726
rect 13728 26240 13780 26246
rect 13728 26182 13780 26188
rect 13740 26042 13768 26182
rect 13728 26036 13780 26042
rect 13728 25978 13780 25984
rect 13832 25974 13860 26998
rect 14016 26858 14044 27118
rect 14004 26852 14056 26858
rect 14004 26794 14056 26800
rect 14004 26580 14056 26586
rect 14004 26522 14056 26528
rect 14016 26234 14044 26522
rect 14108 26450 14136 28086
rect 14740 28076 14792 28082
rect 14740 28018 14792 28024
rect 14280 27328 14332 27334
rect 14280 27270 14332 27276
rect 14188 27124 14240 27130
rect 14188 27066 14240 27072
rect 14096 26444 14148 26450
rect 14096 26386 14148 26392
rect 14200 26382 14228 27066
rect 14292 26994 14320 27270
rect 14280 26988 14332 26994
rect 14280 26930 14332 26936
rect 14372 26988 14424 26994
rect 14372 26930 14424 26936
rect 14384 26874 14412 26930
rect 14752 26926 14780 28018
rect 15752 27872 15804 27878
rect 15752 27814 15804 27820
rect 16120 27872 16172 27878
rect 16120 27814 16172 27820
rect 15764 27470 15792 27814
rect 15752 27464 15804 27470
rect 15752 27406 15804 27412
rect 15660 27396 15712 27402
rect 15660 27338 15712 27344
rect 15672 27130 15700 27338
rect 15660 27124 15712 27130
rect 15660 27066 15712 27072
rect 15476 26988 15528 26994
rect 15476 26930 15528 26936
rect 14292 26846 14412 26874
rect 14740 26920 14792 26926
rect 14740 26862 14792 26868
rect 14292 26790 14320 26846
rect 14280 26784 14332 26790
rect 14280 26726 14332 26732
rect 14372 26784 14424 26790
rect 14372 26726 14424 26732
rect 14188 26376 14240 26382
rect 14188 26318 14240 26324
rect 14016 26206 14136 26234
rect 14108 26042 14136 26206
rect 14200 26042 14228 26318
rect 14096 26036 14148 26042
rect 14096 25978 14148 25984
rect 14188 26036 14240 26042
rect 14188 25978 14240 25984
rect 13820 25968 13872 25974
rect 13820 25910 13872 25916
rect 13544 25900 13596 25906
rect 13544 25842 13596 25848
rect 13636 25900 13688 25906
rect 13636 25842 13688 25848
rect 13452 25696 13504 25702
rect 13452 25638 13504 25644
rect 13268 25492 13320 25498
rect 13268 25434 13320 25440
rect 13464 24274 13492 25638
rect 13556 25158 13584 25842
rect 13544 25152 13596 25158
rect 13544 25094 13596 25100
rect 13452 24268 13504 24274
rect 13452 24210 13504 24216
rect 13832 24206 13860 25910
rect 14384 25906 14412 26726
rect 15488 26586 15516 26930
rect 15476 26580 15528 26586
rect 15476 26522 15528 26528
rect 15108 26376 15160 26382
rect 15108 26318 15160 26324
rect 14372 25900 14424 25906
rect 14372 25842 14424 25848
rect 14556 25900 14608 25906
rect 14556 25842 14608 25848
rect 14568 25294 14596 25842
rect 14556 25288 14608 25294
rect 14556 25230 14608 25236
rect 14924 25288 14976 25294
rect 14924 25230 14976 25236
rect 13820 24200 13872 24206
rect 13820 24142 13872 24148
rect 13176 24132 13228 24138
rect 13176 24074 13228 24080
rect 14648 24132 14700 24138
rect 14648 24074 14700 24080
rect 13360 24064 13412 24070
rect 13360 24006 13412 24012
rect 13372 23798 13400 24006
rect 14660 23866 14688 24074
rect 14648 23860 14700 23866
rect 14648 23802 14700 23808
rect 13360 23792 13412 23798
rect 13360 23734 13412 23740
rect 14936 23730 14964 25230
rect 15016 24812 15068 24818
rect 15016 24754 15068 24760
rect 13084 23724 13136 23730
rect 13084 23666 13136 23672
rect 14924 23724 14976 23730
rect 14924 23666 14976 23672
rect 13820 23588 13872 23594
rect 13820 23530 13872 23536
rect 12808 23316 12860 23322
rect 12808 23258 12860 23264
rect 12992 23316 13044 23322
rect 12992 23258 13044 23264
rect 13004 23202 13032 23258
rect 13004 23186 13216 23202
rect 13004 23180 13228 23186
rect 13004 23174 13176 23180
rect 13176 23122 13228 23128
rect 12624 23112 12676 23118
rect 12624 23054 12676 23060
rect 12532 22228 12584 22234
rect 12532 22170 12584 22176
rect 12544 22098 12572 22170
rect 12532 22092 12584 22098
rect 12532 22034 12584 22040
rect 12636 21894 12664 23054
rect 13832 23050 13860 23530
rect 14004 23520 14056 23526
rect 14004 23462 14056 23468
rect 13912 23180 13964 23186
rect 13912 23122 13964 23128
rect 13820 23044 13872 23050
rect 13820 22986 13872 22992
rect 12716 22976 12768 22982
rect 12716 22918 12768 22924
rect 12624 21888 12676 21894
rect 12624 21830 12676 21836
rect 12532 21548 12584 21554
rect 12452 21508 12532 21536
rect 12584 21508 12664 21536
rect 12532 21490 12584 21496
rect 12348 20800 12400 20806
rect 12348 20742 12400 20748
rect 12636 20466 12664 21508
rect 12728 21350 12756 22918
rect 13636 22568 13688 22574
rect 13636 22510 13688 22516
rect 12900 22432 12952 22438
rect 12900 22374 12952 22380
rect 13084 22432 13136 22438
rect 13084 22374 13136 22380
rect 12912 22166 12940 22374
rect 12900 22160 12952 22166
rect 12900 22102 12952 22108
rect 12992 22092 13044 22098
rect 12992 22034 13044 22040
rect 12808 21956 12860 21962
rect 12808 21898 12860 21904
rect 12716 21344 12768 21350
rect 12716 21286 12768 21292
rect 12820 21078 12848 21898
rect 13004 21593 13032 22034
rect 13096 21729 13124 22374
rect 13648 22234 13676 22510
rect 13636 22228 13688 22234
rect 13636 22170 13688 22176
rect 13728 22228 13780 22234
rect 13728 22170 13780 22176
rect 13360 22024 13412 22030
rect 13360 21966 13412 21972
rect 13176 21888 13228 21894
rect 13176 21830 13228 21836
rect 13082 21720 13138 21729
rect 13082 21655 13138 21664
rect 12990 21584 13046 21593
rect 12990 21519 13046 21528
rect 12808 21072 12860 21078
rect 12808 21014 12860 21020
rect 12808 20596 12860 20602
rect 12808 20538 12860 20544
rect 12624 20460 12676 20466
rect 12624 20402 12676 20408
rect 11888 20052 11940 20058
rect 11888 19994 11940 20000
rect 12636 19854 12664 20402
rect 12624 19848 12676 19854
rect 12676 19796 12756 19802
rect 12624 19790 12756 19796
rect 12636 19774 12756 19790
rect 10784 19508 10836 19514
rect 10784 19450 10836 19456
rect 11428 19508 11480 19514
rect 11428 19450 11480 19456
rect 10232 19440 10284 19446
rect 10232 19382 10284 19388
rect 10324 19440 10376 19446
rect 10324 19382 10376 19388
rect 10140 18896 10192 18902
rect 10140 18838 10192 18844
rect 9956 18760 10008 18766
rect 9956 18702 10008 18708
rect 10048 18760 10100 18766
rect 10048 18702 10100 18708
rect 9772 18420 9824 18426
rect 9772 18362 9824 18368
rect 9968 17882 9996 18702
rect 10048 18284 10100 18290
rect 10048 18226 10100 18232
rect 9956 17876 10008 17882
rect 9956 17818 10008 17824
rect 10060 17814 10088 18226
rect 10244 17814 10272 19382
rect 11796 19372 11848 19378
rect 11796 19314 11848 19320
rect 11704 19304 11756 19310
rect 11704 19246 11756 19252
rect 10416 19236 10468 19242
rect 10416 19178 10468 19184
rect 11244 19236 11296 19242
rect 11244 19178 11296 19184
rect 10428 18970 10456 19178
rect 11152 19168 11204 19174
rect 11152 19110 11204 19116
rect 10416 18964 10468 18970
rect 10416 18906 10468 18912
rect 10692 18896 10744 18902
rect 10692 18838 10744 18844
rect 10324 18692 10376 18698
rect 10324 18634 10376 18640
rect 10336 18426 10364 18634
rect 10324 18420 10376 18426
rect 10324 18362 10376 18368
rect 10508 18080 10560 18086
rect 10508 18022 10560 18028
rect 10048 17808 10100 17814
rect 10048 17750 10100 17756
rect 10232 17808 10284 17814
rect 10232 17750 10284 17756
rect 10520 17678 10548 18022
rect 10704 17882 10732 18838
rect 11164 18834 11192 19110
rect 11256 18970 11284 19178
rect 11244 18964 11296 18970
rect 11244 18906 11296 18912
rect 11152 18828 11204 18834
rect 11152 18770 11204 18776
rect 11716 18766 11744 19246
rect 11612 18760 11664 18766
rect 11612 18702 11664 18708
rect 11704 18760 11756 18766
rect 11704 18702 11756 18708
rect 10968 18624 11020 18630
rect 11020 18584 11100 18612
rect 10968 18566 11020 18572
rect 10692 17876 10744 17882
rect 10692 17818 10744 17824
rect 9680 17672 9732 17678
rect 9680 17614 9732 17620
rect 10508 17672 10560 17678
rect 10508 17614 10560 17620
rect 10704 17338 10732 17818
rect 10876 17536 10928 17542
rect 10876 17478 10928 17484
rect 10140 17332 10192 17338
rect 10140 17274 10192 17280
rect 10692 17332 10744 17338
rect 10692 17274 10744 17280
rect 10048 17196 10100 17202
rect 10048 17138 10100 17144
rect 9588 17128 9640 17134
rect 9588 17070 9640 17076
rect 9600 16794 9628 17070
rect 9956 16992 10008 16998
rect 9956 16934 10008 16940
rect 9588 16788 9640 16794
rect 9588 16730 9640 16736
rect 9496 16720 9548 16726
rect 9496 16662 9548 16668
rect 9968 16658 9996 16934
rect 10060 16794 10088 17138
rect 10048 16788 10100 16794
rect 10048 16730 10100 16736
rect 9956 16652 10008 16658
rect 9956 16594 10008 16600
rect 9404 16584 9456 16590
rect 9404 16526 9456 16532
rect 9680 16516 9732 16522
rect 9680 16458 9732 16464
rect 8944 16448 8996 16454
rect 8944 16390 8996 16396
rect 8576 16040 8628 16046
rect 8576 15982 8628 15988
rect 8852 16040 8904 16046
rect 8852 15982 8904 15988
rect 8392 15496 8444 15502
rect 8392 15438 8444 15444
rect 8484 15496 8536 15502
rect 8484 15438 8536 15444
rect 8864 15434 8892 15982
rect 8852 15428 8904 15434
rect 8852 15370 8904 15376
rect 8392 15360 8444 15366
rect 8392 15302 8444 15308
rect 8404 15162 8432 15302
rect 8392 15156 8444 15162
rect 8392 15098 8444 15104
rect 8864 14958 8892 15370
rect 9692 15162 9720 16458
rect 9956 16108 10008 16114
rect 9956 16050 10008 16056
rect 9864 15904 9916 15910
rect 9864 15846 9916 15852
rect 9680 15156 9732 15162
rect 9680 15098 9732 15104
rect 9036 15088 9088 15094
rect 9036 15030 9088 15036
rect 8852 14952 8904 14958
rect 8852 14894 8904 14900
rect 8760 14884 8812 14890
rect 8760 14826 8812 14832
rect 8668 14816 8720 14822
rect 8668 14758 8720 14764
rect 8680 14482 8708 14758
rect 8668 14476 8720 14482
rect 8668 14418 8720 14424
rect 8576 14408 8628 14414
rect 8576 14350 8628 14356
rect 7708 13892 7788 13920
rect 7656 13874 7708 13880
rect 7840 13796 7892 13802
rect 7840 13738 7892 13744
rect 7656 13184 7708 13190
rect 7656 13126 7708 13132
rect 7012 12232 7064 12238
rect 7012 12174 7064 12180
rect 7380 12232 7432 12238
rect 7380 12174 7432 12180
rect 7564 12232 7616 12238
rect 7564 12174 7616 12180
rect 7024 12102 7052 12174
rect 7012 12096 7064 12102
rect 7012 12038 7064 12044
rect 6920 11756 6972 11762
rect 6920 11698 6972 11704
rect 6828 11688 6880 11694
rect 6828 11630 6880 11636
rect 7472 11688 7524 11694
rect 7472 11630 7524 11636
rect 6840 10062 6868 11630
rect 7484 10674 7512 11630
rect 7576 11218 7604 12174
rect 7564 11212 7616 11218
rect 7564 11154 7616 11160
rect 7472 10668 7524 10674
rect 7472 10610 7524 10616
rect 7196 10464 7248 10470
rect 7196 10406 7248 10412
rect 6828 10056 6880 10062
rect 6828 9998 6880 10004
rect 7208 9586 7236 10406
rect 7484 10130 7512 10610
rect 7472 10124 7524 10130
rect 7472 10066 7524 10072
rect 7472 9920 7524 9926
rect 7472 9862 7524 9868
rect 7484 9654 7512 9862
rect 7472 9648 7524 9654
rect 7472 9590 7524 9596
rect 7196 9580 7248 9586
rect 7196 9522 7248 9528
rect 7208 9382 7236 9522
rect 7196 9376 7248 9382
rect 7196 9318 7248 9324
rect 6736 8968 6788 8974
rect 6736 8910 6788 8916
rect 7472 8832 7524 8838
rect 7472 8774 7524 8780
rect 6828 8560 6880 8566
rect 6828 8502 6880 8508
rect 6736 8424 6788 8430
rect 6736 8366 6788 8372
rect 6748 7818 6776 8366
rect 6736 7812 6788 7818
rect 6736 7754 6788 7760
rect 6552 7744 6604 7750
rect 6552 7686 6604 7692
rect 6564 7410 6592 7686
rect 6644 7540 6696 7546
rect 6644 7482 6696 7488
rect 6552 7404 6604 7410
rect 6552 7346 6604 7352
rect 6552 7268 6604 7274
rect 6380 7228 6552 7256
rect 6288 6934 6316 7210
rect 6276 6928 6328 6934
rect 6276 6870 6328 6876
rect 6380 6798 6408 7228
rect 6552 7210 6604 7216
rect 6368 6792 6420 6798
rect 6368 6734 6420 6740
rect 6184 6656 6236 6662
rect 6184 6598 6236 6604
rect 6196 6322 6224 6598
rect 6656 6390 6684 7482
rect 6748 7410 6776 7754
rect 6736 7404 6788 7410
rect 6736 7346 6788 7352
rect 6736 6656 6788 6662
rect 6736 6598 6788 6604
rect 6748 6458 6776 6598
rect 6736 6452 6788 6458
rect 6736 6394 6788 6400
rect 6644 6384 6696 6390
rect 6644 6326 6696 6332
rect 6184 6316 6236 6322
rect 6184 6258 6236 6264
rect 6092 5704 6144 5710
rect 6092 5646 6144 5652
rect 6000 5568 6052 5574
rect 6000 5510 6052 5516
rect 6104 5370 6132 5646
rect 6644 5568 6696 5574
rect 6644 5510 6696 5516
rect 6092 5364 6144 5370
rect 6092 5306 6144 5312
rect 6104 5250 6132 5306
rect 5724 5228 5776 5234
rect 5724 5170 5776 5176
rect 5908 5228 5960 5234
rect 6104 5222 6224 5250
rect 6656 5234 6684 5510
rect 6748 5234 6776 6394
rect 6840 6322 6868 8502
rect 7484 7410 7512 8774
rect 7668 7886 7696 13126
rect 7852 9518 7880 13738
rect 7932 13728 7984 13734
rect 7932 13670 7984 13676
rect 8024 13728 8076 13734
rect 8024 13670 8076 13676
rect 7944 13530 7972 13670
rect 7932 13524 7984 13530
rect 7932 13466 7984 13472
rect 8036 13462 8064 13670
rect 8024 13456 8076 13462
rect 8024 13398 8076 13404
rect 8116 13184 8168 13190
rect 8116 13126 8168 13132
rect 8024 12844 8076 12850
rect 8024 12786 8076 12792
rect 7932 12640 7984 12646
rect 7932 12582 7984 12588
rect 7944 11558 7972 12582
rect 8036 12442 8064 12786
rect 8128 12646 8156 13126
rect 8116 12640 8168 12646
rect 8116 12582 8168 12588
rect 8024 12436 8076 12442
rect 8024 12378 8076 12384
rect 8220 12306 8248 14214
rect 8312 14198 8524 14226
rect 8392 12844 8444 12850
rect 8312 12804 8392 12832
rect 8208 12300 8260 12306
rect 8208 12242 8260 12248
rect 8220 12186 8248 12242
rect 8036 12158 8248 12186
rect 8036 12102 8064 12158
rect 8024 12096 8076 12102
rect 8024 12038 8076 12044
rect 8116 12096 8168 12102
rect 8116 12038 8168 12044
rect 8128 11830 8156 12038
rect 8116 11824 8168 11830
rect 8116 11766 8168 11772
rect 7932 11552 7984 11558
rect 7932 11494 7984 11500
rect 8208 11552 8260 11558
rect 8208 11494 8260 11500
rect 8220 11286 8248 11494
rect 8312 11354 8340 12804
rect 8392 12786 8444 12792
rect 8392 12708 8444 12714
rect 8392 12650 8444 12656
rect 8404 12442 8432 12650
rect 8392 12436 8444 12442
rect 8392 12378 8444 12384
rect 8392 12232 8444 12238
rect 8496 12220 8524 14198
rect 8588 14074 8616 14350
rect 8576 14068 8628 14074
rect 8576 14010 8628 14016
rect 8772 13802 8800 14826
rect 8864 14550 8892 14894
rect 8944 14884 8996 14890
rect 8944 14826 8996 14832
rect 8852 14544 8904 14550
rect 8852 14486 8904 14492
rect 8760 13796 8812 13802
rect 8760 13738 8812 13744
rect 8772 13530 8800 13738
rect 8760 13524 8812 13530
rect 8760 13466 8812 13472
rect 8956 13326 8984 14826
rect 9048 14482 9076 15030
rect 9680 15020 9732 15026
rect 9680 14962 9732 14968
rect 9036 14476 9088 14482
rect 9036 14418 9088 14424
rect 9692 14414 9720 14962
rect 9680 14408 9732 14414
rect 9680 14350 9732 14356
rect 9772 14340 9824 14346
rect 9772 14282 9824 14288
rect 9496 14272 9548 14278
rect 9496 14214 9548 14220
rect 9128 13728 9180 13734
rect 9128 13670 9180 13676
rect 9140 13326 9168 13670
rect 8944 13320 8996 13326
rect 8944 13262 8996 13268
rect 9128 13320 9180 13326
rect 9128 13262 9180 13268
rect 9036 13184 9088 13190
rect 9036 13126 9088 13132
rect 8576 12436 8628 12442
rect 8576 12378 8628 12384
rect 8444 12192 8524 12220
rect 8392 12174 8444 12180
rect 8588 11354 8616 12378
rect 8668 12232 8720 12238
rect 8668 12174 8720 12180
rect 8680 11762 8708 12174
rect 9048 12170 9076 13126
rect 9128 12368 9180 12374
rect 9128 12310 9180 12316
rect 9036 12164 9088 12170
rect 9036 12106 9088 12112
rect 8668 11756 8720 11762
rect 8668 11698 8720 11704
rect 8300 11348 8352 11354
rect 8300 11290 8352 11296
rect 8392 11348 8444 11354
rect 8392 11290 8444 11296
rect 8576 11348 8628 11354
rect 8576 11290 8628 11296
rect 8208 11280 8260 11286
rect 8208 11222 8260 11228
rect 8220 10062 8248 11222
rect 8404 11150 8432 11290
rect 9048 11218 9076 12106
rect 9140 11762 9168 12310
rect 9508 12238 9536 14214
rect 9784 14006 9812 14282
rect 9772 14000 9824 14006
rect 9772 13942 9824 13948
rect 9876 13870 9904 15846
rect 9968 14958 9996 16050
rect 10152 14958 10180 17274
rect 10232 17128 10284 17134
rect 10284 17088 10364 17116
rect 10232 17070 10284 17076
rect 10232 16992 10284 16998
rect 10232 16934 10284 16940
rect 10244 16182 10272 16934
rect 10232 16176 10284 16182
rect 10232 16118 10284 16124
rect 10336 16096 10364 17088
rect 10600 16788 10652 16794
rect 10600 16730 10652 16736
rect 10612 16114 10640 16730
rect 10692 16516 10744 16522
rect 10692 16458 10744 16464
rect 10704 16114 10732 16458
rect 10888 16182 10916 17478
rect 11072 16794 11100 18584
rect 11520 18420 11572 18426
rect 11520 18362 11572 18368
rect 11152 18284 11204 18290
rect 11152 18226 11204 18232
rect 11164 17202 11192 18226
rect 11244 17740 11296 17746
rect 11244 17682 11296 17688
rect 11152 17196 11204 17202
rect 11152 17138 11204 17144
rect 11060 16788 11112 16794
rect 11060 16730 11112 16736
rect 10784 16176 10836 16182
rect 10784 16118 10836 16124
rect 10876 16176 10928 16182
rect 10876 16118 10928 16124
rect 11060 16176 11112 16182
rect 11060 16118 11112 16124
rect 10416 16108 10468 16114
rect 10336 16068 10416 16096
rect 10600 16108 10652 16114
rect 10416 16050 10468 16056
rect 10520 16068 10600 16096
rect 10428 15910 10456 16050
rect 10416 15904 10468 15910
rect 10416 15846 10468 15852
rect 10520 15042 10548 16068
rect 10600 16050 10652 16056
rect 10692 16108 10744 16114
rect 10692 16050 10744 16056
rect 10600 15904 10652 15910
rect 10600 15846 10652 15852
rect 10244 15014 10548 15042
rect 10612 15026 10640 15846
rect 10704 15094 10732 16050
rect 10692 15088 10744 15094
rect 10692 15030 10744 15036
rect 10600 15020 10652 15026
rect 9956 14952 10008 14958
rect 9956 14894 10008 14900
rect 10140 14952 10192 14958
rect 10140 14894 10192 14900
rect 10048 14884 10100 14890
rect 10048 14826 10100 14832
rect 10060 14346 10088 14826
rect 10140 14816 10192 14822
rect 10140 14758 10192 14764
rect 10152 14618 10180 14758
rect 10140 14612 10192 14618
rect 10140 14554 10192 14560
rect 10048 14340 10100 14346
rect 10048 14282 10100 14288
rect 9864 13864 9916 13870
rect 9864 13806 9916 13812
rect 10152 13802 10180 14554
rect 10140 13796 10192 13802
rect 10140 13738 10192 13744
rect 10152 13326 10180 13738
rect 9772 13320 9824 13326
rect 9772 13262 9824 13268
rect 10140 13320 10192 13326
rect 10140 13262 10192 13268
rect 9784 12442 9812 13262
rect 10140 13184 10192 13190
rect 10140 13126 10192 13132
rect 10152 12850 10180 13126
rect 10140 12844 10192 12850
rect 10140 12786 10192 12792
rect 9772 12436 9824 12442
rect 9772 12378 9824 12384
rect 9784 12238 9812 12378
rect 10244 12238 10272 15014
rect 10600 14962 10652 14968
rect 10508 14952 10560 14958
rect 10508 14894 10560 14900
rect 10416 14272 10468 14278
rect 10416 14214 10468 14220
rect 10324 13728 10376 13734
rect 10324 13670 10376 13676
rect 10336 13326 10364 13670
rect 10324 13320 10376 13326
rect 10324 13262 10376 13268
rect 10324 12980 10376 12986
rect 10324 12922 10376 12928
rect 10336 12850 10364 12922
rect 10428 12850 10456 14214
rect 10520 13938 10548 14894
rect 10508 13932 10560 13938
rect 10508 13874 10560 13880
rect 10520 13326 10548 13874
rect 10612 13870 10640 14962
rect 10796 14906 10824 16118
rect 10888 14958 10916 16118
rect 11072 15586 11100 16118
rect 11152 15904 11204 15910
rect 11256 15892 11284 17682
rect 11336 17264 11388 17270
rect 11336 17206 11388 17212
rect 11348 16017 11376 17206
rect 11532 16658 11560 18362
rect 11624 17882 11652 18702
rect 11612 17876 11664 17882
rect 11612 17818 11664 17824
rect 11704 17604 11756 17610
rect 11704 17546 11756 17552
rect 11612 17060 11664 17066
rect 11612 17002 11664 17008
rect 11520 16652 11572 16658
rect 11520 16594 11572 16600
rect 11334 16008 11390 16017
rect 11334 15943 11336 15952
rect 11388 15943 11390 15952
rect 11336 15914 11388 15920
rect 11204 15864 11284 15892
rect 11152 15846 11204 15852
rect 10980 15558 11100 15586
rect 10980 15162 11008 15558
rect 11164 15434 11192 15846
rect 11152 15428 11204 15434
rect 11204 15388 11284 15416
rect 11152 15370 11204 15376
rect 10968 15156 11020 15162
rect 10968 15098 11020 15104
rect 10980 15008 11008 15098
rect 11150 15056 11206 15065
rect 11060 15020 11112 15026
rect 10980 14980 11060 15008
rect 10704 14878 10824 14906
rect 10876 14952 10928 14958
rect 10876 14894 10928 14900
rect 10704 14278 10732 14878
rect 10980 14618 11008 14980
rect 11150 14991 11152 15000
rect 11060 14962 11112 14968
rect 11204 14991 11206 15000
rect 11152 14962 11204 14968
rect 10968 14612 11020 14618
rect 10968 14554 11020 14560
rect 10784 14544 10836 14550
rect 10784 14486 10836 14492
rect 10692 14272 10744 14278
rect 10692 14214 10744 14220
rect 10704 14006 10732 14214
rect 10692 14000 10744 14006
rect 10692 13942 10744 13948
rect 10600 13864 10652 13870
rect 10600 13806 10652 13812
rect 10612 13394 10640 13806
rect 10600 13388 10652 13394
rect 10600 13330 10652 13336
rect 10508 13320 10560 13326
rect 10508 13262 10560 13268
rect 10692 13184 10744 13190
rect 10692 13126 10744 13132
rect 10704 12850 10732 13126
rect 10796 12918 10824 14486
rect 11256 14414 11284 15388
rect 11244 14408 11296 14414
rect 11244 14350 11296 14356
rect 11060 13864 11112 13870
rect 11060 13806 11112 13812
rect 11072 13530 11100 13806
rect 11060 13524 11112 13530
rect 11060 13466 11112 13472
rect 10784 12912 10836 12918
rect 10784 12854 10836 12860
rect 10324 12844 10376 12850
rect 10324 12786 10376 12792
rect 10416 12844 10468 12850
rect 10416 12786 10468 12792
rect 10692 12844 10744 12850
rect 10692 12786 10744 12792
rect 10876 12640 10928 12646
rect 10876 12582 10928 12588
rect 11244 12640 11296 12646
rect 11244 12582 11296 12588
rect 9496 12232 9548 12238
rect 9496 12174 9548 12180
rect 9772 12232 9824 12238
rect 9772 12174 9824 12180
rect 10232 12232 10284 12238
rect 10232 12174 10284 12180
rect 10784 12232 10836 12238
rect 10784 12174 10836 12180
rect 10796 11762 10824 12174
rect 9128 11756 9180 11762
rect 9128 11698 9180 11704
rect 9404 11756 9456 11762
rect 9404 11698 9456 11704
rect 10324 11756 10376 11762
rect 10324 11698 10376 11704
rect 10784 11756 10836 11762
rect 10784 11698 10836 11704
rect 9036 11212 9088 11218
rect 9036 11154 9088 11160
rect 8392 11144 8444 11150
rect 8392 11086 8444 11092
rect 9048 11082 9076 11154
rect 9416 11150 9444 11698
rect 9404 11144 9456 11150
rect 9404 11086 9456 11092
rect 9036 11076 9088 11082
rect 9036 11018 9088 11024
rect 8300 11008 8352 11014
rect 8300 10950 8352 10956
rect 8208 10056 8260 10062
rect 8208 9998 8260 10004
rect 8312 9994 8340 10950
rect 9048 10742 9076 11018
rect 9128 11008 9180 11014
rect 9128 10950 9180 10956
rect 9036 10736 9088 10742
rect 9036 10678 9088 10684
rect 9140 10674 9168 10950
rect 9128 10668 9180 10674
rect 9128 10610 9180 10616
rect 9312 10668 9364 10674
rect 9312 10610 9364 10616
rect 8392 10600 8444 10606
rect 8392 10542 8444 10548
rect 8300 9988 8352 9994
rect 8300 9930 8352 9936
rect 8116 9920 8168 9926
rect 8116 9862 8168 9868
rect 8208 9920 8260 9926
rect 8208 9862 8260 9868
rect 7840 9512 7892 9518
rect 7840 9454 7892 9460
rect 7852 8974 7880 9454
rect 8128 8974 8156 9862
rect 8220 9722 8248 9862
rect 8208 9716 8260 9722
rect 8208 9658 8260 9664
rect 8220 9178 8248 9658
rect 8208 9172 8260 9178
rect 8208 9114 8260 9120
rect 7840 8968 7892 8974
rect 7840 8910 7892 8916
rect 8116 8968 8168 8974
rect 8116 8910 8168 8916
rect 7748 8832 7800 8838
rect 7748 8774 7800 8780
rect 7656 7880 7708 7886
rect 7576 7828 7656 7834
rect 7576 7822 7708 7828
rect 7576 7806 7696 7822
rect 7472 7404 7524 7410
rect 7472 7346 7524 7352
rect 6828 6316 6880 6322
rect 6828 6258 6880 6264
rect 5908 5170 5960 5176
rect 4804 5092 4856 5098
rect 4804 5034 4856 5040
rect 4896 5024 4948 5030
rect 4896 4966 4948 4972
rect 5448 5024 5500 5030
rect 5448 4966 5500 4972
rect 4908 4622 4936 4966
rect 5460 4622 5488 4966
rect 5736 4690 5764 5170
rect 5724 4684 5776 4690
rect 5724 4626 5776 4632
rect 6196 4622 6224 5222
rect 6644 5228 6696 5234
rect 6644 5170 6696 5176
rect 6736 5228 6788 5234
rect 6736 5170 6788 5176
rect 6840 5166 6868 6258
rect 6828 5160 6880 5166
rect 6828 5102 6880 5108
rect 6552 4752 6604 4758
rect 6552 4694 6604 4700
rect 4620 4616 4672 4622
rect 4620 4558 4672 4564
rect 4896 4616 4948 4622
rect 4896 4558 4948 4564
rect 5448 4616 5500 4622
rect 5448 4558 5500 4564
rect 6184 4616 6236 4622
rect 6184 4558 6236 4564
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 6564 4282 6592 4694
rect 7484 4622 7512 7346
rect 7576 6322 7604 7806
rect 7656 7336 7708 7342
rect 7656 7278 7708 7284
rect 7668 6730 7696 7278
rect 7656 6724 7708 6730
rect 7656 6666 7708 6672
rect 7668 6458 7696 6666
rect 7656 6452 7708 6458
rect 7656 6394 7708 6400
rect 7760 6322 7788 8774
rect 8300 8288 8352 8294
rect 8300 8230 8352 8236
rect 7840 8084 7892 8090
rect 7840 8026 7892 8032
rect 7852 7886 7880 8026
rect 7840 7880 7892 7886
rect 7840 7822 7892 7828
rect 8116 7880 8168 7886
rect 8116 7822 8168 7828
rect 8128 7342 8156 7822
rect 8312 7410 8340 8230
rect 8404 7834 8432 10542
rect 9324 10130 9352 10610
rect 9312 10124 9364 10130
rect 9312 10066 9364 10072
rect 8760 9988 8812 9994
rect 8760 9930 8812 9936
rect 8772 9654 8800 9930
rect 9324 9722 9352 10066
rect 9312 9716 9364 9722
rect 9312 9658 9364 9664
rect 8760 9648 8812 9654
rect 8760 9590 8812 9596
rect 9416 9518 9444 11086
rect 9772 11076 9824 11082
rect 9772 11018 9824 11024
rect 9496 10668 9548 10674
rect 9496 10610 9548 10616
rect 9508 10062 9536 10610
rect 9496 10056 9548 10062
rect 9496 9998 9548 10004
rect 8576 9512 8628 9518
rect 8576 9454 8628 9460
rect 9404 9512 9456 9518
rect 9404 9454 9456 9460
rect 8588 7886 8616 9454
rect 9784 9042 9812 11018
rect 10336 11014 10364 11698
rect 10324 11008 10376 11014
rect 10324 10950 10376 10956
rect 9864 10464 9916 10470
rect 9864 10406 9916 10412
rect 9772 9036 9824 9042
rect 9772 8978 9824 8984
rect 9784 8430 9812 8978
rect 9876 8430 9904 10406
rect 10048 9920 10100 9926
rect 10048 9862 10100 9868
rect 9772 8424 9824 8430
rect 9772 8366 9824 8372
rect 9864 8424 9916 8430
rect 9864 8366 9916 8372
rect 9220 8356 9272 8362
rect 9220 8298 9272 8304
rect 8944 8084 8996 8090
rect 8944 8026 8996 8032
rect 8956 7886 8984 8026
rect 9232 7954 9260 8298
rect 9772 8288 9824 8294
rect 9772 8230 9824 8236
rect 9220 7948 9272 7954
rect 9220 7890 9272 7896
rect 9784 7886 9812 8230
rect 9876 7886 9904 8366
rect 10060 8294 10088 9862
rect 10336 9586 10364 10950
rect 10796 10062 10824 11698
rect 10888 11150 10916 12582
rect 10968 11688 11020 11694
rect 10968 11630 11020 11636
rect 10980 11150 11008 11630
rect 10876 11144 10928 11150
rect 10876 11086 10928 11092
rect 10968 11144 11020 11150
rect 10968 11086 11020 11092
rect 10784 10056 10836 10062
rect 10784 9998 10836 10004
rect 10324 9580 10376 9586
rect 10324 9522 10376 9528
rect 11256 9042 11284 12582
rect 11336 12096 11388 12102
rect 11336 12038 11388 12044
rect 11348 11150 11376 12038
rect 11532 11694 11560 16594
rect 11624 12238 11652 17002
rect 11716 16674 11744 17546
rect 11808 17338 11836 19314
rect 12440 19304 12492 19310
rect 12440 19246 12492 19252
rect 12348 19236 12400 19242
rect 12348 19178 12400 19184
rect 12360 18970 12388 19178
rect 12348 18964 12400 18970
rect 12348 18906 12400 18912
rect 12164 18760 12216 18766
rect 12084 18720 12164 18748
rect 11980 18692 12032 18698
rect 11980 18634 12032 18640
rect 11992 18290 12020 18634
rect 12084 18290 12112 18720
rect 12164 18702 12216 18708
rect 12360 18426 12388 18906
rect 12452 18698 12480 19246
rect 12440 18692 12492 18698
rect 12440 18634 12492 18640
rect 12624 18624 12676 18630
rect 12624 18566 12676 18572
rect 12348 18420 12400 18426
rect 12348 18362 12400 18368
rect 11980 18284 12032 18290
rect 11980 18226 12032 18232
rect 12072 18284 12124 18290
rect 12072 18226 12124 18232
rect 11796 17332 11848 17338
rect 11796 17274 11848 17280
rect 12084 17066 12112 18226
rect 12636 17814 12664 18566
rect 12728 18086 12756 19774
rect 12820 19378 12848 20538
rect 13084 19848 13136 19854
rect 13084 19790 13136 19796
rect 13096 19378 13124 19790
rect 13188 19378 13216 21830
rect 13372 21622 13400 21966
rect 13648 21894 13676 22170
rect 13740 22098 13768 22170
rect 13728 22092 13780 22098
rect 13728 22034 13780 22040
rect 13832 22030 13860 22986
rect 13924 22710 13952 23122
rect 14016 22982 14044 23462
rect 15028 23118 15056 24754
rect 15120 24070 15148 26318
rect 15488 25974 15516 26522
rect 15476 25968 15528 25974
rect 15476 25910 15528 25916
rect 15764 25906 15792 27406
rect 16132 27402 16160 27814
rect 16120 27396 16172 27402
rect 16120 27338 16172 27344
rect 16028 26988 16080 26994
rect 16028 26930 16080 26936
rect 16488 26988 16540 26994
rect 16488 26930 16540 26936
rect 15936 26376 15988 26382
rect 15936 26318 15988 26324
rect 15752 25900 15804 25906
rect 15752 25842 15804 25848
rect 15948 25498 15976 26318
rect 16040 25974 16068 26930
rect 16120 26920 16172 26926
rect 16120 26862 16172 26868
rect 16132 26042 16160 26862
rect 16500 26586 16528 26930
rect 16488 26580 16540 26586
rect 16488 26522 16540 26528
rect 16592 26518 16620 28154
rect 16764 28076 16816 28082
rect 16764 28018 16816 28024
rect 16776 27606 16804 28018
rect 16868 27878 16896 28426
rect 17052 28218 17080 28494
rect 17132 28416 17184 28422
rect 17132 28358 17184 28364
rect 17040 28212 17092 28218
rect 17040 28154 17092 28160
rect 16856 27872 16908 27878
rect 16856 27814 16908 27820
rect 16764 27600 16816 27606
rect 16764 27542 16816 27548
rect 16868 26994 16896 27814
rect 17144 27674 17172 28358
rect 18604 28144 18656 28150
rect 18604 28086 18656 28092
rect 18144 27872 18196 27878
rect 18144 27814 18196 27820
rect 18236 27872 18288 27878
rect 18236 27814 18288 27820
rect 17132 27668 17184 27674
rect 17132 27610 17184 27616
rect 17144 27538 17172 27610
rect 18156 27538 18184 27814
rect 18248 27606 18276 27814
rect 18236 27600 18288 27606
rect 18236 27542 18288 27548
rect 17132 27532 17184 27538
rect 17132 27474 17184 27480
rect 18144 27532 18196 27538
rect 18144 27474 18196 27480
rect 16856 26988 16908 26994
rect 16856 26930 16908 26936
rect 17316 26988 17368 26994
rect 17316 26930 17368 26936
rect 16672 26580 16724 26586
rect 16672 26522 16724 26528
rect 16580 26512 16632 26518
rect 16580 26454 16632 26460
rect 16592 26246 16620 26454
rect 16580 26240 16632 26246
rect 16580 26182 16632 26188
rect 16120 26036 16172 26042
rect 16120 25978 16172 25984
rect 16028 25968 16080 25974
rect 16028 25910 16080 25916
rect 16488 25832 16540 25838
rect 16488 25774 16540 25780
rect 15936 25492 15988 25498
rect 15936 25434 15988 25440
rect 15476 25152 15528 25158
rect 15476 25094 15528 25100
rect 15384 24812 15436 24818
rect 15384 24754 15436 24760
rect 15200 24200 15252 24206
rect 15200 24142 15252 24148
rect 15108 24064 15160 24070
rect 15108 24006 15160 24012
rect 14648 23112 14700 23118
rect 14648 23054 14700 23060
rect 15016 23112 15068 23118
rect 15016 23054 15068 23060
rect 14004 22976 14056 22982
rect 14004 22918 14056 22924
rect 14660 22778 14688 23054
rect 14648 22772 14700 22778
rect 14648 22714 14700 22720
rect 13912 22704 13964 22710
rect 13912 22646 13964 22652
rect 14372 22500 14424 22506
rect 14372 22442 14424 22448
rect 13820 22024 13872 22030
rect 13820 21966 13872 21972
rect 13636 21888 13688 21894
rect 13636 21830 13688 21836
rect 13648 21690 13676 21830
rect 13636 21684 13688 21690
rect 13636 21626 13688 21632
rect 13360 21616 13412 21622
rect 13360 21558 13412 21564
rect 13372 20602 13400 21558
rect 13912 21344 13964 21350
rect 13912 21286 13964 21292
rect 13820 21004 13872 21010
rect 13820 20946 13872 20952
rect 13360 20596 13412 20602
rect 13360 20538 13412 20544
rect 13832 20482 13860 20946
rect 13740 20466 13860 20482
rect 13728 20460 13860 20466
rect 13780 20454 13860 20460
rect 13728 20402 13780 20408
rect 13452 20256 13504 20262
rect 13452 20198 13504 20204
rect 12808 19372 12860 19378
rect 12808 19314 12860 19320
rect 12900 19372 12952 19378
rect 12900 19314 12952 19320
rect 13084 19372 13136 19378
rect 13084 19314 13136 19320
rect 13176 19372 13228 19378
rect 13176 19314 13228 19320
rect 13360 19372 13412 19378
rect 13360 19314 13412 19320
rect 12716 18080 12768 18086
rect 12716 18022 12768 18028
rect 12624 17808 12676 17814
rect 12624 17750 12676 17756
rect 12728 17678 12756 18022
rect 12912 17746 12940 19314
rect 12992 18216 13044 18222
rect 12992 18158 13044 18164
rect 13004 17882 13032 18158
rect 12992 17876 13044 17882
rect 12992 17818 13044 17824
rect 12900 17740 12952 17746
rect 12900 17682 12952 17688
rect 12164 17672 12216 17678
rect 12164 17614 12216 17620
rect 12716 17672 12768 17678
rect 12716 17614 12768 17620
rect 12072 17060 12124 17066
rect 12072 17002 12124 17008
rect 11716 16646 11836 16674
rect 11704 16516 11756 16522
rect 11704 16458 11756 16464
rect 11716 16250 11744 16458
rect 11704 16244 11756 16250
rect 11704 16186 11756 16192
rect 11716 15706 11744 16186
rect 11808 15910 11836 16646
rect 11980 16652 12032 16658
rect 11980 16594 12032 16600
rect 11888 16584 11940 16590
rect 11888 16526 11940 16532
rect 11900 16114 11928 16526
rect 11888 16108 11940 16114
rect 11888 16050 11940 16056
rect 11796 15904 11848 15910
rect 11796 15846 11848 15852
rect 11704 15700 11756 15706
rect 11704 15642 11756 15648
rect 11808 15638 11836 15846
rect 11796 15632 11848 15638
rect 11796 15574 11848 15580
rect 11900 15162 11928 16050
rect 11992 15570 12020 16594
rect 12176 16590 12204 17614
rect 12440 16992 12492 16998
rect 12440 16934 12492 16940
rect 12164 16584 12216 16590
rect 12164 16526 12216 16532
rect 12452 16266 12480 16934
rect 12452 16250 12572 16266
rect 12452 16244 12584 16250
rect 12452 16238 12532 16244
rect 12532 16186 12584 16192
rect 11980 15564 12032 15570
rect 11980 15506 12032 15512
rect 12544 15502 12572 16186
rect 12532 15496 12584 15502
rect 12532 15438 12584 15444
rect 11888 15156 11940 15162
rect 11888 15098 11940 15104
rect 12348 15156 12400 15162
rect 12348 15098 12400 15104
rect 12360 14346 12388 15098
rect 12728 14890 12756 17614
rect 13096 17610 13124 19314
rect 13174 19000 13230 19009
rect 13174 18935 13176 18944
rect 13228 18935 13230 18944
rect 13176 18906 13228 18912
rect 13188 17678 13216 18906
rect 13372 18834 13400 19314
rect 13464 19310 13492 20198
rect 13820 19780 13872 19786
rect 13820 19722 13872 19728
rect 13832 19514 13860 19722
rect 13820 19508 13872 19514
rect 13820 19450 13872 19456
rect 13924 19378 13952 21286
rect 14384 21185 14412 22442
rect 14660 22030 14688 22714
rect 14648 22024 14700 22030
rect 14648 21966 14700 21972
rect 14924 21888 14976 21894
rect 14924 21830 14976 21836
rect 14648 21684 14700 21690
rect 14648 21626 14700 21632
rect 14556 21412 14608 21418
rect 14556 21354 14608 21360
rect 14370 21176 14426 21185
rect 14370 21111 14426 21120
rect 14096 21072 14148 21078
rect 14096 21014 14148 21020
rect 14004 20868 14056 20874
rect 14004 20810 14056 20816
rect 14016 19514 14044 20810
rect 14108 19854 14136 21014
rect 14186 20496 14242 20505
rect 14186 20431 14188 20440
rect 14240 20431 14242 20440
rect 14188 20402 14240 20408
rect 14188 20256 14240 20262
rect 14188 20198 14240 20204
rect 14096 19848 14148 19854
rect 14096 19790 14148 19796
rect 14004 19508 14056 19514
rect 14004 19450 14056 19456
rect 14200 19378 14228 20198
rect 14280 19712 14332 19718
rect 14280 19654 14332 19660
rect 14292 19446 14320 19654
rect 14280 19440 14332 19446
rect 14280 19382 14332 19388
rect 13912 19372 13964 19378
rect 13912 19314 13964 19320
rect 14188 19372 14240 19378
rect 14188 19314 14240 19320
rect 13452 19304 13504 19310
rect 14200 19281 14228 19314
rect 13452 19246 13504 19252
rect 14186 19272 14242 19281
rect 14186 19207 14242 19216
rect 13544 19168 13596 19174
rect 13544 19110 13596 19116
rect 13360 18828 13412 18834
rect 13360 18770 13412 18776
rect 13268 18760 13320 18766
rect 13268 18702 13320 18708
rect 13176 17672 13228 17678
rect 13176 17614 13228 17620
rect 13084 17604 13136 17610
rect 13084 17546 13136 17552
rect 12808 16992 12860 16998
rect 12808 16934 12860 16940
rect 12820 16590 12848 16934
rect 13096 16794 13124 17546
rect 13280 17542 13308 18702
rect 13556 17882 13584 19110
rect 13544 17876 13596 17882
rect 13544 17818 13596 17824
rect 14292 17746 14320 19382
rect 14280 17740 14332 17746
rect 14280 17682 14332 17688
rect 13912 17672 13964 17678
rect 13912 17614 13964 17620
rect 13268 17536 13320 17542
rect 13268 17478 13320 17484
rect 13820 17196 13872 17202
rect 13820 17138 13872 17144
rect 13084 16788 13136 16794
rect 13084 16730 13136 16736
rect 13452 16652 13504 16658
rect 13452 16594 13504 16600
rect 12808 16584 12860 16590
rect 12808 16526 12860 16532
rect 12820 16114 12848 16526
rect 13268 16448 13320 16454
rect 13268 16390 13320 16396
rect 13280 16114 13308 16390
rect 13464 16182 13492 16594
rect 13832 16250 13860 17138
rect 13924 17134 13952 17614
rect 13912 17128 13964 17134
rect 13912 17070 13964 17076
rect 13924 16794 13952 17070
rect 13912 16788 13964 16794
rect 13912 16730 13964 16736
rect 14292 16658 14320 17682
rect 14280 16652 14332 16658
rect 14280 16594 14332 16600
rect 14384 16590 14412 21111
rect 14568 20466 14596 21354
rect 14660 21350 14688 21626
rect 14936 21554 14964 21830
rect 14924 21548 14976 21554
rect 14924 21490 14976 21496
rect 14648 21344 14700 21350
rect 14648 21286 14700 21292
rect 14936 21010 14964 21490
rect 14924 21004 14976 21010
rect 14924 20946 14976 20952
rect 14740 20800 14792 20806
rect 14740 20742 14792 20748
rect 14556 20460 14608 20466
rect 14556 20402 14608 20408
rect 14648 19984 14700 19990
rect 14648 19926 14700 19932
rect 14556 19780 14608 19786
rect 14556 19722 14608 19728
rect 14568 18698 14596 19722
rect 14660 19718 14688 19926
rect 14648 19712 14700 19718
rect 14648 19654 14700 19660
rect 14660 19310 14688 19654
rect 14752 19310 14780 20742
rect 15028 20058 15056 23054
rect 15108 21344 15160 21350
rect 15108 21286 15160 21292
rect 15120 20874 15148 21286
rect 15108 20868 15160 20874
rect 15108 20810 15160 20816
rect 15016 20052 15068 20058
rect 15016 19994 15068 20000
rect 14924 19712 14976 19718
rect 14924 19654 14976 19660
rect 14936 19378 14964 19654
rect 14924 19372 14976 19378
rect 14924 19314 14976 19320
rect 14648 19304 14700 19310
rect 14648 19246 14700 19252
rect 14740 19304 14792 19310
rect 14740 19246 14792 19252
rect 14752 19122 14780 19246
rect 14660 19094 14780 19122
rect 14832 19168 14884 19174
rect 14832 19110 14884 19116
rect 14660 18834 14688 19094
rect 14648 18828 14700 18834
rect 14648 18770 14700 18776
rect 14740 18760 14792 18766
rect 14844 18748 14872 19110
rect 14792 18720 14872 18748
rect 14740 18702 14792 18708
rect 14556 18692 14608 18698
rect 14556 18634 14608 18640
rect 14740 17672 14792 17678
rect 14740 17614 14792 17620
rect 14752 17338 14780 17614
rect 14740 17332 14792 17338
rect 14740 17274 14792 17280
rect 14372 16584 14424 16590
rect 14372 16526 14424 16532
rect 14740 16516 14792 16522
rect 14740 16458 14792 16464
rect 14280 16448 14332 16454
rect 14280 16390 14332 16396
rect 13820 16244 13872 16250
rect 13820 16186 13872 16192
rect 13452 16176 13504 16182
rect 13452 16118 13504 16124
rect 12808 16108 12860 16114
rect 12808 16050 12860 16056
rect 13268 16108 13320 16114
rect 13268 16050 13320 16056
rect 12716 14884 12768 14890
rect 12716 14826 12768 14832
rect 12820 14414 12848 16050
rect 12900 16040 12952 16046
rect 12900 15982 12952 15988
rect 12912 14482 12940 15982
rect 13464 15366 13492 16118
rect 14292 16114 14320 16390
rect 13544 16108 13596 16114
rect 13544 16050 13596 16056
rect 14280 16108 14332 16114
rect 14280 16050 14332 16056
rect 13268 15360 13320 15366
rect 13268 15302 13320 15308
rect 13452 15360 13504 15366
rect 13452 15302 13504 15308
rect 13280 15026 13308 15302
rect 13464 15065 13492 15302
rect 13556 15201 13584 16050
rect 13728 15972 13780 15978
rect 13728 15914 13780 15920
rect 13542 15192 13598 15201
rect 13542 15127 13598 15136
rect 13450 15056 13506 15065
rect 13268 15020 13320 15026
rect 13450 14991 13506 15000
rect 13268 14962 13320 14968
rect 13176 14952 13228 14958
rect 13176 14894 13228 14900
rect 12992 14816 13044 14822
rect 12992 14758 13044 14764
rect 13004 14618 13032 14758
rect 13188 14618 13216 14894
rect 13360 14884 13412 14890
rect 13360 14826 13412 14832
rect 12992 14612 13044 14618
rect 12992 14554 13044 14560
rect 13176 14612 13228 14618
rect 13176 14554 13228 14560
rect 12900 14476 12952 14482
rect 12900 14418 12952 14424
rect 13004 14414 13032 14554
rect 12808 14408 12860 14414
rect 12808 14350 12860 14356
rect 12992 14408 13044 14414
rect 12992 14350 13044 14356
rect 12348 14340 12400 14346
rect 12348 14282 12400 14288
rect 12360 13938 12388 14282
rect 12348 13932 12400 13938
rect 12348 13874 12400 13880
rect 13372 13920 13400 14826
rect 13556 13988 13584 15127
rect 13740 15094 13768 15914
rect 13820 15564 13872 15570
rect 13820 15506 13872 15512
rect 13832 15094 13860 15506
rect 14096 15360 14148 15366
rect 14096 15302 14148 15308
rect 13728 15088 13780 15094
rect 13728 15030 13780 15036
rect 13820 15088 13872 15094
rect 13820 15030 13872 15036
rect 13728 14952 13780 14958
rect 13728 14894 13780 14900
rect 13740 14550 13768 14894
rect 13832 14890 13860 15030
rect 14004 15020 14056 15026
rect 14004 14962 14056 14968
rect 13820 14884 13872 14890
rect 13820 14826 13872 14832
rect 14016 14618 14044 14962
rect 14004 14612 14056 14618
rect 14004 14554 14056 14560
rect 13728 14544 13780 14550
rect 13728 14486 13780 14492
rect 13728 14000 13780 14006
rect 13556 13960 13728 13988
rect 13452 13932 13504 13938
rect 13372 13892 13452 13920
rect 11796 13184 11848 13190
rect 11796 13126 11848 13132
rect 11808 12238 11836 13126
rect 13176 12640 13228 12646
rect 13176 12582 13228 12588
rect 11612 12232 11664 12238
rect 11612 12174 11664 12180
rect 11796 12232 11848 12238
rect 11796 12174 11848 12180
rect 12164 12232 12216 12238
rect 12164 12174 12216 12180
rect 12176 11898 12204 12174
rect 12440 12096 12492 12102
rect 12440 12038 12492 12044
rect 12624 12096 12676 12102
rect 12624 12038 12676 12044
rect 12164 11892 12216 11898
rect 12164 11834 12216 11840
rect 12452 11762 12480 12038
rect 12636 11762 12664 12038
rect 13188 11830 13216 12582
rect 13176 11824 13228 11830
rect 13176 11766 13228 11772
rect 13372 11762 13400 13892
rect 13452 13874 13504 13880
rect 13556 12889 13584 13960
rect 13728 13942 13780 13948
rect 13820 13932 13872 13938
rect 13820 13874 13872 13880
rect 13912 13932 13964 13938
rect 13912 13874 13964 13880
rect 13832 13530 13860 13874
rect 13924 13734 13952 13874
rect 13912 13728 13964 13734
rect 13912 13670 13964 13676
rect 13820 13524 13872 13530
rect 13820 13466 13872 13472
rect 13542 12880 13598 12889
rect 13542 12815 13544 12824
rect 13596 12815 13598 12824
rect 13544 12786 13596 12792
rect 14016 12782 14044 14554
rect 14108 14006 14136 15302
rect 14752 15162 14780 16458
rect 14844 16130 14872 18720
rect 14936 17338 14964 19314
rect 15028 18358 15056 19994
rect 15212 18766 15240 24142
rect 15396 23882 15424 24754
rect 15304 23866 15424 23882
rect 15488 23866 15516 25094
rect 15948 24954 15976 25434
rect 16500 25226 16528 25774
rect 16488 25220 16540 25226
rect 16488 25162 16540 25168
rect 15936 24948 15988 24954
rect 15936 24890 15988 24896
rect 15568 24064 15620 24070
rect 15568 24006 15620 24012
rect 15292 23860 15424 23866
rect 15344 23854 15424 23860
rect 15476 23860 15528 23866
rect 15292 23802 15344 23808
rect 15476 23802 15528 23808
rect 15580 23730 15608 24006
rect 15948 23730 15976 24890
rect 16500 24682 16528 25162
rect 16684 25158 16712 26522
rect 16868 26314 16896 26930
rect 17132 26920 17184 26926
rect 17132 26862 17184 26868
rect 17144 26586 17172 26862
rect 17132 26580 17184 26586
rect 17132 26522 17184 26528
rect 16856 26308 16908 26314
rect 16856 26250 16908 26256
rect 16948 26308 17000 26314
rect 16948 26250 17000 26256
rect 17224 26308 17276 26314
rect 17224 26250 17276 26256
rect 16868 25906 16896 26250
rect 16856 25900 16908 25906
rect 16856 25842 16908 25848
rect 16960 25702 16988 26250
rect 17040 26240 17092 26246
rect 17040 26182 17092 26188
rect 17052 25820 17080 26182
rect 17236 25974 17264 26250
rect 17224 25968 17276 25974
rect 17224 25910 17276 25916
rect 17328 25906 17356 26930
rect 17500 26852 17552 26858
rect 17500 26794 17552 26800
rect 17512 26042 17540 26794
rect 17592 26784 17644 26790
rect 17592 26726 17644 26732
rect 17604 26382 17632 26726
rect 17592 26376 17644 26382
rect 17592 26318 17644 26324
rect 18156 26314 18184 27474
rect 18616 26994 18644 28086
rect 18512 26988 18564 26994
rect 18512 26930 18564 26936
rect 18604 26988 18656 26994
rect 18604 26930 18656 26936
rect 20996 26988 21048 26994
rect 20996 26930 21048 26936
rect 18524 26586 18552 26930
rect 18512 26580 18564 26586
rect 18512 26522 18564 26528
rect 18616 26382 18644 26930
rect 20076 26784 20128 26790
rect 20076 26726 20128 26732
rect 20088 26382 20116 26726
rect 21008 26450 21036 26930
rect 20996 26444 21048 26450
rect 20996 26386 21048 26392
rect 18604 26376 18656 26382
rect 18604 26318 18656 26324
rect 20076 26376 20128 26382
rect 20076 26318 20128 26324
rect 18144 26308 18196 26314
rect 18144 26250 18196 26256
rect 17500 26036 17552 26042
rect 17500 25978 17552 25984
rect 17316 25900 17368 25906
rect 17316 25842 17368 25848
rect 17224 25832 17276 25838
rect 17052 25792 17224 25820
rect 17224 25774 17276 25780
rect 16948 25696 17000 25702
rect 16948 25638 17000 25644
rect 18616 25362 18644 26318
rect 21008 26024 21036 26386
rect 21088 26036 21140 26042
rect 21008 25996 21088 26024
rect 21088 25978 21140 25984
rect 20536 25968 20588 25974
rect 20536 25910 20588 25916
rect 20904 25968 20956 25974
rect 20904 25910 20956 25916
rect 19984 25832 20036 25838
rect 19984 25774 20036 25780
rect 19340 25696 19392 25702
rect 19340 25638 19392 25644
rect 18604 25356 18656 25362
rect 18604 25298 18656 25304
rect 16672 25152 16724 25158
rect 16672 25094 16724 25100
rect 16488 24676 16540 24682
rect 16488 24618 16540 24624
rect 16500 24342 16528 24618
rect 16488 24336 16540 24342
rect 16488 24278 16540 24284
rect 16500 23866 16528 24278
rect 16684 24274 16712 25094
rect 18616 24818 18644 25298
rect 19352 25294 19380 25638
rect 19996 25498 20024 25774
rect 19984 25492 20036 25498
rect 19984 25434 20036 25440
rect 19340 25288 19392 25294
rect 19340 25230 19392 25236
rect 20548 25158 20576 25910
rect 20812 25696 20864 25702
rect 20812 25638 20864 25644
rect 20536 25152 20588 25158
rect 20536 25094 20588 25100
rect 20548 24954 20576 25094
rect 20536 24948 20588 24954
rect 20536 24890 20588 24896
rect 20548 24818 20576 24890
rect 16856 24812 16908 24818
rect 16856 24754 16908 24760
rect 18604 24812 18656 24818
rect 18604 24754 18656 24760
rect 18696 24812 18748 24818
rect 18696 24754 18748 24760
rect 20536 24812 20588 24818
rect 20536 24754 20588 24760
rect 16868 24410 16896 24754
rect 16856 24404 16908 24410
rect 16856 24346 16908 24352
rect 18616 24274 18644 24754
rect 18708 24410 18736 24754
rect 20076 24608 20128 24614
rect 20076 24550 20128 24556
rect 18696 24404 18748 24410
rect 18696 24346 18748 24352
rect 16672 24268 16724 24274
rect 16672 24210 16724 24216
rect 18604 24268 18656 24274
rect 18604 24210 18656 24216
rect 19248 24268 19300 24274
rect 19248 24210 19300 24216
rect 16488 23860 16540 23866
rect 16488 23802 16540 23808
rect 16684 23730 16712 24210
rect 15568 23724 15620 23730
rect 15568 23666 15620 23672
rect 15936 23724 15988 23730
rect 15936 23666 15988 23672
rect 16672 23724 16724 23730
rect 16672 23666 16724 23672
rect 19260 23186 19288 24210
rect 20088 24138 20116 24550
rect 20824 24410 20852 25638
rect 20916 25498 20944 25910
rect 20996 25696 21048 25702
rect 20996 25638 21048 25644
rect 20904 25492 20956 25498
rect 20904 25434 20956 25440
rect 21008 25226 21036 25638
rect 20996 25220 21048 25226
rect 20996 25162 21048 25168
rect 20812 24404 20864 24410
rect 20812 24346 20864 24352
rect 19800 24132 19852 24138
rect 19800 24074 19852 24080
rect 20076 24132 20128 24138
rect 20076 24074 20128 24080
rect 19812 23662 19840 24074
rect 20088 23798 20116 24074
rect 21180 24064 21232 24070
rect 21180 24006 21232 24012
rect 20076 23792 20128 23798
rect 20076 23734 20128 23740
rect 21192 23730 21220 24006
rect 21180 23724 21232 23730
rect 21180 23666 21232 23672
rect 19800 23656 19852 23662
rect 19800 23598 19852 23604
rect 20904 23316 20956 23322
rect 20904 23258 20956 23264
rect 20260 23248 20312 23254
rect 20260 23190 20312 23196
rect 19248 23180 19300 23186
rect 19248 23122 19300 23128
rect 16672 23112 16724 23118
rect 16672 23054 16724 23060
rect 16212 22772 16264 22778
rect 16212 22714 16264 22720
rect 15844 22636 15896 22642
rect 16120 22636 16172 22642
rect 15844 22578 15896 22584
rect 16040 22596 16120 22624
rect 15476 22092 15528 22098
rect 15476 22034 15528 22040
rect 15292 21616 15344 21622
rect 15290 21584 15292 21593
rect 15344 21584 15346 21593
rect 15290 21519 15346 21528
rect 15384 21548 15436 21554
rect 15384 21490 15436 21496
rect 15396 21332 15424 21490
rect 15304 21304 15424 21332
rect 15304 21010 15332 21304
rect 15488 21146 15516 22034
rect 15568 22024 15620 22030
rect 15568 21966 15620 21972
rect 15580 21690 15608 21966
rect 15660 21888 15712 21894
rect 15660 21830 15712 21836
rect 15568 21684 15620 21690
rect 15568 21626 15620 21632
rect 15672 21554 15700 21830
rect 15856 21690 15884 22578
rect 16040 22438 16068 22596
rect 16120 22578 16172 22584
rect 16028 22432 16080 22438
rect 16028 22374 16080 22380
rect 15934 21856 15990 21865
rect 15934 21791 15990 21800
rect 15844 21684 15896 21690
rect 15844 21626 15896 21632
rect 15660 21548 15712 21554
rect 15660 21490 15712 21496
rect 15844 21548 15896 21554
rect 15844 21490 15896 21496
rect 15660 21344 15712 21350
rect 15660 21286 15712 21292
rect 15476 21140 15528 21146
rect 15476 21082 15528 21088
rect 15568 21140 15620 21146
rect 15568 21082 15620 21088
rect 15292 21004 15344 21010
rect 15292 20946 15344 20952
rect 15304 20330 15332 20946
rect 15580 20890 15608 21082
rect 15488 20862 15608 20890
rect 15384 20460 15436 20466
rect 15384 20402 15436 20408
rect 15292 20324 15344 20330
rect 15292 20266 15344 20272
rect 15292 20052 15344 20058
rect 15292 19994 15344 20000
rect 15304 19310 15332 19994
rect 15396 19786 15424 20402
rect 15488 19922 15516 20862
rect 15568 20800 15620 20806
rect 15568 20742 15620 20748
rect 15476 19916 15528 19922
rect 15476 19858 15528 19864
rect 15580 19786 15608 20742
rect 15672 19922 15700 21286
rect 15856 20942 15884 21490
rect 15948 21146 15976 21791
rect 16040 21622 16068 22374
rect 16120 22024 16172 22030
rect 16120 21966 16172 21972
rect 16028 21616 16080 21622
rect 16028 21558 16080 21564
rect 16132 21554 16160 21966
rect 16224 21962 16252 22714
rect 16684 22642 16712 23054
rect 17316 23044 17368 23050
rect 17316 22986 17368 22992
rect 18972 23044 19024 23050
rect 18972 22986 19024 22992
rect 17040 22704 17092 22710
rect 17040 22646 17092 22652
rect 16304 22636 16356 22642
rect 16304 22578 16356 22584
rect 16672 22636 16724 22642
rect 16672 22578 16724 22584
rect 16316 22234 16344 22578
rect 16304 22228 16356 22234
rect 16304 22170 16356 22176
rect 16212 21956 16264 21962
rect 16212 21898 16264 21904
rect 16120 21548 16172 21554
rect 16120 21490 16172 21496
rect 16028 21480 16080 21486
rect 16028 21422 16080 21428
rect 16040 21146 16068 21422
rect 15936 21140 15988 21146
rect 15936 21082 15988 21088
rect 16028 21140 16080 21146
rect 16028 21082 16080 21088
rect 16132 21078 16160 21490
rect 16120 21072 16172 21078
rect 16026 21040 16082 21049
rect 16120 21014 16172 21020
rect 16026 20975 16082 20984
rect 15752 20936 15804 20942
rect 15752 20878 15804 20884
rect 15844 20936 15896 20942
rect 15844 20878 15896 20884
rect 15764 20788 15792 20878
rect 16040 20874 16068 20975
rect 16028 20868 16080 20874
rect 15948 20828 16028 20856
rect 15948 20788 15976 20828
rect 16028 20810 16080 20816
rect 15764 20760 15976 20788
rect 15844 20392 15896 20398
rect 15844 20334 15896 20340
rect 15752 20256 15804 20262
rect 15752 20198 15804 20204
rect 15764 20058 15792 20198
rect 15752 20052 15804 20058
rect 15752 19994 15804 20000
rect 15660 19916 15712 19922
rect 15660 19858 15712 19864
rect 15384 19780 15436 19786
rect 15384 19722 15436 19728
rect 15568 19780 15620 19786
rect 15568 19722 15620 19728
rect 15476 19712 15528 19718
rect 15476 19654 15528 19660
rect 15488 19394 15516 19654
rect 15396 19378 15516 19394
rect 15672 19378 15700 19858
rect 15384 19372 15516 19378
rect 15436 19366 15516 19372
rect 15660 19372 15712 19378
rect 15384 19314 15436 19320
rect 15660 19314 15712 19320
rect 15752 19372 15804 19378
rect 15752 19314 15804 19320
rect 15292 19304 15344 19310
rect 15292 19246 15344 19252
rect 15292 18896 15344 18902
rect 15292 18838 15344 18844
rect 15200 18760 15252 18766
rect 15200 18702 15252 18708
rect 15016 18352 15068 18358
rect 15016 18294 15068 18300
rect 15304 17814 15332 18838
rect 15396 18698 15424 19314
rect 15476 18760 15528 18766
rect 15764 18714 15792 19314
rect 15476 18702 15528 18708
rect 15384 18692 15436 18698
rect 15384 18634 15436 18640
rect 15488 18086 15516 18702
rect 15672 18686 15792 18714
rect 15476 18080 15528 18086
rect 15476 18022 15528 18028
rect 15292 17808 15344 17814
rect 15292 17750 15344 17756
rect 15200 17672 15252 17678
rect 15200 17614 15252 17620
rect 15212 17354 15240 17614
rect 14924 17332 14976 17338
rect 14924 17274 14976 17280
rect 15120 17326 15240 17354
rect 14936 16250 14964 17274
rect 15120 17202 15148 17326
rect 15108 17196 15160 17202
rect 15108 17138 15160 17144
rect 15304 17116 15332 17750
rect 15384 17128 15436 17134
rect 15304 17088 15384 17116
rect 15304 16538 15332 17088
rect 15384 17070 15436 17076
rect 15488 16794 15516 18022
rect 15568 17536 15620 17542
rect 15568 17478 15620 17484
rect 15580 17134 15608 17478
rect 15672 17202 15700 18686
rect 15752 18624 15804 18630
rect 15752 18566 15804 18572
rect 15764 17202 15792 18566
rect 15856 17746 15884 20334
rect 16120 20052 16172 20058
rect 16120 19994 16172 20000
rect 15936 19848 15988 19854
rect 15936 19790 15988 19796
rect 15948 19514 15976 19790
rect 15936 19508 15988 19514
rect 15936 19450 15988 19456
rect 16132 18834 16160 19994
rect 16120 18828 16172 18834
rect 16120 18770 16172 18776
rect 16028 17876 16080 17882
rect 16028 17818 16080 17824
rect 15844 17740 15896 17746
rect 15844 17682 15896 17688
rect 16040 17202 16068 17818
rect 16132 17542 16160 18770
rect 16224 17678 16252 21898
rect 16316 21894 16344 22170
rect 16948 22160 17000 22166
rect 16948 22102 17000 22108
rect 16672 22024 16724 22030
rect 16672 21966 16724 21972
rect 16304 21888 16356 21894
rect 16304 21830 16356 21836
rect 16684 21690 16712 21966
rect 16960 21962 16988 22102
rect 17052 22030 17080 22646
rect 17328 22234 17356 22986
rect 18788 22976 18840 22982
rect 18788 22918 18840 22924
rect 18696 22636 18748 22642
rect 18696 22578 18748 22584
rect 18144 22568 18196 22574
rect 18144 22510 18196 22516
rect 17316 22228 17368 22234
rect 17316 22170 17368 22176
rect 18156 22098 18184 22510
rect 18144 22092 18196 22098
rect 18144 22034 18196 22040
rect 18708 22030 18736 22578
rect 18800 22574 18828 22918
rect 18984 22778 19012 22986
rect 18972 22772 19024 22778
rect 18972 22714 19024 22720
rect 18788 22568 18840 22574
rect 18788 22510 18840 22516
rect 19260 22098 19288 23122
rect 19340 22636 19392 22642
rect 19340 22578 19392 22584
rect 19248 22092 19300 22098
rect 19248 22034 19300 22040
rect 19352 22030 19380 22578
rect 20272 22574 20300 23190
rect 20812 23180 20864 23186
rect 20812 23122 20864 23128
rect 20720 23112 20772 23118
rect 20720 23054 20772 23060
rect 20260 22568 20312 22574
rect 20260 22510 20312 22516
rect 17040 22024 17092 22030
rect 17040 21966 17092 21972
rect 17592 22024 17644 22030
rect 17868 22024 17920 22030
rect 17592 21966 17644 21972
rect 17774 21992 17830 22001
rect 16948 21956 17000 21962
rect 16948 21898 17000 21904
rect 16764 21888 16816 21894
rect 16764 21830 16816 21836
rect 17316 21888 17368 21894
rect 17604 21865 17632 21966
rect 17868 21966 17920 21972
rect 18420 22024 18472 22030
rect 18420 21966 18472 21972
rect 18696 22024 18748 22030
rect 18696 21966 18748 21972
rect 19340 22024 19392 22030
rect 19340 21966 19392 21972
rect 17774 21927 17830 21936
rect 17788 21894 17816 21927
rect 17776 21888 17828 21894
rect 17316 21830 17368 21836
rect 17590 21856 17646 21865
rect 16672 21684 16724 21690
rect 16672 21626 16724 21632
rect 16396 21616 16448 21622
rect 16396 21558 16448 21564
rect 16408 21486 16436 21558
rect 16396 21480 16448 21486
rect 16396 21422 16448 21428
rect 16302 20904 16358 20913
rect 16302 20839 16358 20848
rect 16316 20806 16344 20839
rect 16304 20800 16356 20806
rect 16304 20742 16356 20748
rect 16304 19848 16356 19854
rect 16304 19790 16356 19796
rect 16316 18222 16344 19790
rect 16408 19786 16436 21422
rect 16396 19780 16448 19786
rect 16396 19722 16448 19728
rect 16672 19780 16724 19786
rect 16672 19722 16724 19728
rect 16408 19009 16436 19722
rect 16684 19514 16712 19722
rect 16672 19508 16724 19514
rect 16672 19450 16724 19456
rect 16776 19378 16804 21830
rect 17328 21622 17356 21830
rect 17776 21830 17828 21836
rect 17590 21791 17646 21800
rect 17316 21616 17368 21622
rect 17316 21558 17368 21564
rect 17500 21616 17552 21622
rect 17500 21558 17552 21564
rect 17040 21548 17092 21554
rect 17040 21490 17092 21496
rect 17224 21548 17276 21554
rect 17224 21490 17276 21496
rect 17052 21457 17080 21490
rect 17038 21448 17094 21457
rect 17236 21434 17264 21490
rect 17512 21434 17540 21558
rect 17236 21406 17540 21434
rect 17592 21480 17644 21486
rect 17592 21422 17644 21428
rect 17038 21383 17094 21392
rect 16948 20800 17000 20806
rect 16948 20742 17000 20748
rect 16960 20534 16988 20742
rect 16948 20528 17000 20534
rect 16948 20470 17000 20476
rect 17052 19854 17080 21383
rect 17604 21146 17632 21422
rect 17500 21140 17552 21146
rect 17500 21082 17552 21088
rect 17592 21140 17644 21146
rect 17592 21082 17644 21088
rect 17512 21010 17540 21082
rect 17788 21049 17816 21830
rect 17880 21350 17908 21966
rect 18052 21888 18104 21894
rect 18050 21856 18052 21865
rect 18104 21856 18106 21865
rect 18050 21791 18106 21800
rect 18432 21690 18460 21966
rect 18604 21956 18656 21962
rect 18604 21898 18656 21904
rect 18616 21690 18644 21898
rect 20732 21894 20760 23054
rect 20168 21888 20220 21894
rect 19706 21856 19762 21865
rect 20168 21830 20220 21836
rect 20720 21888 20772 21894
rect 20720 21830 20772 21836
rect 19706 21791 19762 21800
rect 18420 21684 18472 21690
rect 18420 21626 18472 21632
rect 18604 21684 18656 21690
rect 18604 21626 18656 21632
rect 18696 21548 18748 21554
rect 18696 21490 18748 21496
rect 18052 21480 18104 21486
rect 18052 21422 18104 21428
rect 17868 21344 17920 21350
rect 17868 21286 17920 21292
rect 17774 21040 17830 21049
rect 17500 21004 17552 21010
rect 17774 20975 17830 20984
rect 17500 20946 17552 20952
rect 17880 20913 17908 21286
rect 18064 20942 18092 21422
rect 18512 21412 18564 21418
rect 18512 21354 18564 21360
rect 18524 20942 18552 21354
rect 18604 21344 18656 21350
rect 18604 21286 18656 21292
rect 18616 21146 18644 21286
rect 18708 21146 18736 21490
rect 18970 21176 19026 21185
rect 18604 21140 18656 21146
rect 18604 21082 18656 21088
rect 18696 21140 18748 21146
rect 18970 21111 19026 21120
rect 18696 21082 18748 21088
rect 18984 20942 19012 21111
rect 18052 20936 18104 20942
rect 17866 20904 17922 20913
rect 18052 20878 18104 20884
rect 18512 20936 18564 20942
rect 18512 20878 18564 20884
rect 18604 20936 18656 20942
rect 18604 20878 18656 20884
rect 18972 20936 19024 20942
rect 18972 20878 19024 20884
rect 17866 20839 17922 20848
rect 17684 20460 17736 20466
rect 17684 20402 17736 20408
rect 17696 20058 17724 20402
rect 17684 20052 17736 20058
rect 17684 19994 17736 20000
rect 17040 19848 17092 19854
rect 17040 19790 17092 19796
rect 16856 19712 16908 19718
rect 16856 19654 16908 19660
rect 17776 19712 17828 19718
rect 17776 19654 17828 19660
rect 16868 19378 16896 19654
rect 17788 19378 17816 19654
rect 18064 19378 18092 20878
rect 18616 19854 18644 20878
rect 18788 20528 18840 20534
rect 18788 20470 18840 20476
rect 18800 20058 18828 20470
rect 18788 20052 18840 20058
rect 18788 19994 18840 20000
rect 18696 19916 18748 19922
rect 18696 19858 18748 19864
rect 18604 19848 18656 19854
rect 18604 19790 18656 19796
rect 18328 19780 18380 19786
rect 18328 19722 18380 19728
rect 16764 19372 16816 19378
rect 16764 19314 16816 19320
rect 16856 19372 16908 19378
rect 16856 19314 16908 19320
rect 17040 19372 17092 19378
rect 17040 19314 17092 19320
rect 17776 19372 17828 19378
rect 17776 19314 17828 19320
rect 18052 19372 18104 19378
rect 18052 19314 18104 19320
rect 17052 19281 17080 19314
rect 17038 19272 17094 19281
rect 17038 19207 17094 19216
rect 16394 19000 16450 19009
rect 16394 18935 16450 18944
rect 16304 18216 16356 18222
rect 16304 18158 16356 18164
rect 16212 17672 16264 17678
rect 16212 17614 16264 17620
rect 16304 17604 16356 17610
rect 16304 17546 16356 17552
rect 16120 17536 16172 17542
rect 16120 17478 16172 17484
rect 16316 17202 16344 17546
rect 15660 17196 15712 17202
rect 15660 17138 15712 17144
rect 15752 17196 15804 17202
rect 15752 17138 15804 17144
rect 16028 17196 16080 17202
rect 16028 17138 16080 17144
rect 16304 17196 16356 17202
rect 16304 17138 16356 17144
rect 15568 17128 15620 17134
rect 15568 17070 15620 17076
rect 16316 17066 16344 17138
rect 16304 17060 16356 17066
rect 16304 17002 16356 17008
rect 15476 16788 15528 16794
rect 15476 16730 15528 16736
rect 15212 16510 15332 16538
rect 15212 16250 15240 16510
rect 14924 16244 14976 16250
rect 14924 16186 14976 16192
rect 15200 16244 15252 16250
rect 15200 16186 15252 16192
rect 14844 16102 14964 16130
rect 14740 15156 14792 15162
rect 14740 15098 14792 15104
rect 14188 15020 14240 15026
rect 14188 14962 14240 14968
rect 14200 14618 14228 14962
rect 14740 14952 14792 14958
rect 14740 14894 14792 14900
rect 14372 14816 14424 14822
rect 14372 14758 14424 14764
rect 14188 14612 14240 14618
rect 14188 14554 14240 14560
rect 14384 14482 14412 14758
rect 14752 14482 14780 14894
rect 14372 14476 14424 14482
rect 14372 14418 14424 14424
rect 14740 14476 14792 14482
rect 14740 14418 14792 14424
rect 14280 14272 14332 14278
rect 14280 14214 14332 14220
rect 14096 14000 14148 14006
rect 14096 13942 14148 13948
rect 14004 12776 14056 12782
rect 14004 12718 14056 12724
rect 14108 12714 14136 13942
rect 14292 13938 14320 14214
rect 14280 13932 14332 13938
rect 14280 13874 14332 13880
rect 14384 13818 14412 14418
rect 14556 13932 14608 13938
rect 14556 13874 14608 13880
rect 14292 13790 14412 13818
rect 14292 13530 14320 13790
rect 14372 13728 14424 13734
rect 14372 13670 14424 13676
rect 14280 13524 14332 13530
rect 14280 13466 14332 13472
rect 14384 13326 14412 13670
rect 14568 13326 14596 13874
rect 14372 13320 14424 13326
rect 14372 13262 14424 13268
rect 14556 13320 14608 13326
rect 14556 13262 14608 13268
rect 14832 13252 14884 13258
rect 14832 13194 14884 13200
rect 14556 13184 14608 13190
rect 14556 13126 14608 13132
rect 14568 12850 14596 13126
rect 14844 12986 14872 13194
rect 14832 12980 14884 12986
rect 14832 12922 14884 12928
rect 14556 12844 14608 12850
rect 14556 12786 14608 12792
rect 14648 12776 14700 12782
rect 14648 12718 14700 12724
rect 14096 12708 14148 12714
rect 14096 12650 14148 12656
rect 14660 11898 14688 12718
rect 14936 12434 14964 16102
rect 15108 16108 15160 16114
rect 15108 16050 15160 16056
rect 15016 16040 15068 16046
rect 15120 16017 15148 16050
rect 15016 15982 15068 15988
rect 15106 16008 15162 16017
rect 15028 15502 15056 15982
rect 15106 15943 15162 15952
rect 15488 15502 15516 16730
rect 15568 16584 15620 16590
rect 15568 16526 15620 16532
rect 15016 15496 15068 15502
rect 15016 15438 15068 15444
rect 15384 15496 15436 15502
rect 15384 15438 15436 15444
rect 15476 15496 15528 15502
rect 15476 15438 15528 15444
rect 15028 14414 15056 15438
rect 15396 15366 15424 15438
rect 15200 15360 15252 15366
rect 15200 15302 15252 15308
rect 15384 15360 15436 15366
rect 15384 15302 15436 15308
rect 15106 15192 15162 15201
rect 15106 15127 15162 15136
rect 15120 15094 15148 15127
rect 15212 15094 15240 15302
rect 15108 15088 15160 15094
rect 15108 15030 15160 15036
rect 15200 15088 15252 15094
rect 15200 15030 15252 15036
rect 15396 14958 15424 15302
rect 15384 14952 15436 14958
rect 15384 14894 15436 14900
rect 15384 14816 15436 14822
rect 15384 14758 15436 14764
rect 15016 14408 15068 14414
rect 15016 14350 15068 14356
rect 15396 13462 15424 14758
rect 15384 13456 15436 13462
rect 15384 13398 15436 13404
rect 15292 13320 15344 13326
rect 15292 13262 15344 13268
rect 15108 13252 15160 13258
rect 15108 13194 15160 13200
rect 15120 12714 15148 13194
rect 15304 12850 15332 13262
rect 15396 12918 15424 13398
rect 15384 12912 15436 12918
rect 15384 12854 15436 12860
rect 15292 12844 15344 12850
rect 15292 12786 15344 12792
rect 15108 12708 15160 12714
rect 15108 12650 15160 12656
rect 15292 12640 15344 12646
rect 15292 12582 15344 12588
rect 14844 12406 14964 12434
rect 14648 11892 14700 11898
rect 14648 11834 14700 11840
rect 11704 11756 11756 11762
rect 11704 11698 11756 11704
rect 11796 11756 11848 11762
rect 11796 11698 11848 11704
rect 12440 11756 12492 11762
rect 12440 11698 12492 11704
rect 12624 11756 12676 11762
rect 12624 11698 12676 11704
rect 13360 11756 13412 11762
rect 13360 11698 13412 11704
rect 11520 11688 11572 11694
rect 11520 11630 11572 11636
rect 11612 11552 11664 11558
rect 11612 11494 11664 11500
rect 11336 11144 11388 11150
rect 11336 11086 11388 11092
rect 11428 9104 11480 9110
rect 11428 9046 11480 9052
rect 10140 9036 10192 9042
rect 10140 8978 10192 8984
rect 11244 9036 11296 9042
rect 11244 8978 11296 8984
rect 10152 8634 10180 8978
rect 11060 8968 11112 8974
rect 10980 8916 11060 8922
rect 10980 8910 11112 8916
rect 11152 8968 11204 8974
rect 11152 8910 11204 8916
rect 10980 8894 11100 8910
rect 10140 8628 10192 8634
rect 10140 8570 10192 8576
rect 10152 8498 10180 8570
rect 10140 8492 10192 8498
rect 10140 8434 10192 8440
rect 10048 8288 10100 8294
rect 10048 8230 10100 8236
rect 10060 7886 10088 8230
rect 8484 7880 8536 7886
rect 8404 7828 8484 7834
rect 8404 7822 8536 7828
rect 8576 7880 8628 7886
rect 8576 7822 8628 7828
rect 8944 7880 8996 7886
rect 8944 7822 8996 7828
rect 9772 7880 9824 7886
rect 9772 7822 9824 7828
rect 9864 7880 9916 7886
rect 9864 7822 9916 7828
rect 10048 7880 10100 7886
rect 10048 7822 10100 7828
rect 8404 7806 8524 7822
rect 9588 7812 9640 7818
rect 8404 7478 8432 7806
rect 9588 7754 9640 7760
rect 8668 7744 8720 7750
rect 8668 7686 8720 7692
rect 9496 7744 9548 7750
rect 9496 7686 9548 7692
rect 8392 7472 8444 7478
rect 8392 7414 8444 7420
rect 8300 7404 8352 7410
rect 8300 7346 8352 7352
rect 8116 7336 8168 7342
rect 8116 7278 8168 7284
rect 8312 6934 8340 7346
rect 8300 6928 8352 6934
rect 8300 6870 8352 6876
rect 7564 6316 7616 6322
rect 7564 6258 7616 6264
rect 7748 6316 7800 6322
rect 7748 6258 7800 6264
rect 7576 5710 7604 6258
rect 7656 5772 7708 5778
rect 7760 5760 7788 6258
rect 7708 5732 7788 5760
rect 7932 5772 7984 5778
rect 7656 5714 7708 5720
rect 7932 5714 7984 5720
rect 7564 5704 7616 5710
rect 7564 5646 7616 5652
rect 7944 5234 7972 5714
rect 8404 5642 8432 7414
rect 8680 7410 8708 7686
rect 9508 7478 9536 7686
rect 9496 7472 9548 7478
rect 9496 7414 9548 7420
rect 8668 7404 8720 7410
rect 8668 7346 8720 7352
rect 8852 7200 8904 7206
rect 8852 7142 8904 7148
rect 8864 6798 8892 7142
rect 8852 6792 8904 6798
rect 8852 6734 8904 6740
rect 9600 5710 9628 7754
rect 9876 7478 9904 7822
rect 9864 7472 9916 7478
rect 9864 7414 9916 7420
rect 10060 7410 10088 7822
rect 10980 7410 11008 8894
rect 11060 8832 11112 8838
rect 11060 8774 11112 8780
rect 11072 7546 11100 8774
rect 11164 8498 11192 8910
rect 11244 8900 11296 8906
rect 11244 8842 11296 8848
rect 11256 8498 11284 8842
rect 11152 8492 11204 8498
rect 11152 8434 11204 8440
rect 11244 8492 11296 8498
rect 11296 8452 11376 8480
rect 11244 8434 11296 8440
rect 11164 8090 11192 8434
rect 11244 8288 11296 8294
rect 11244 8230 11296 8236
rect 11152 8084 11204 8090
rect 11152 8026 11204 8032
rect 11060 7540 11112 7546
rect 11060 7482 11112 7488
rect 10048 7404 10100 7410
rect 10048 7346 10100 7352
rect 10968 7404 11020 7410
rect 10968 7346 11020 7352
rect 9772 6724 9824 6730
rect 9772 6666 9824 6672
rect 9784 5778 9812 6666
rect 10060 6322 10088 7346
rect 10980 7274 11008 7346
rect 10968 7268 11020 7274
rect 10968 7210 11020 7216
rect 10692 7200 10744 7206
rect 10692 7142 10744 7148
rect 10876 7200 10928 7206
rect 10876 7142 10928 7148
rect 10416 6928 10468 6934
rect 10416 6870 10468 6876
rect 10428 6798 10456 6870
rect 10704 6798 10732 7142
rect 10888 6798 10916 7142
rect 11072 6934 11100 7482
rect 11256 7478 11284 8230
rect 11348 7886 11376 8452
rect 11440 7954 11468 9046
rect 11624 8974 11652 11494
rect 11716 11354 11744 11698
rect 11704 11348 11756 11354
rect 11704 11290 11756 11296
rect 11716 9586 11744 11290
rect 11808 11082 11836 11698
rect 12532 11620 12584 11626
rect 12532 11562 12584 11568
rect 12544 11150 12572 11562
rect 12624 11552 12676 11558
rect 12624 11494 12676 11500
rect 12636 11218 12664 11494
rect 12624 11212 12676 11218
rect 12624 11154 12676 11160
rect 12992 11212 13044 11218
rect 12992 11154 13044 11160
rect 12532 11144 12584 11150
rect 12532 11086 12584 11092
rect 11796 11076 11848 11082
rect 11796 11018 11848 11024
rect 11808 10554 11836 11018
rect 12348 10668 12400 10674
rect 12348 10610 12400 10616
rect 12440 10668 12492 10674
rect 12440 10610 12492 10616
rect 11808 10526 11928 10554
rect 11796 10464 11848 10470
rect 11796 10406 11848 10412
rect 11704 9580 11756 9586
rect 11704 9522 11756 9528
rect 11808 9518 11836 10406
rect 11900 10266 11928 10526
rect 11888 10260 11940 10266
rect 11888 10202 11940 10208
rect 11900 9654 11928 10202
rect 11888 9648 11940 9654
rect 11888 9590 11940 9596
rect 11796 9512 11848 9518
rect 11796 9454 11848 9460
rect 12072 9444 12124 9450
rect 12072 9386 12124 9392
rect 11612 8968 11664 8974
rect 11612 8910 11664 8916
rect 11428 7948 11480 7954
rect 11428 7890 11480 7896
rect 11336 7880 11388 7886
rect 11336 7822 11388 7828
rect 11244 7472 11296 7478
rect 11244 7414 11296 7420
rect 12084 7410 12112 9386
rect 12360 8974 12388 10610
rect 12348 8968 12400 8974
rect 12348 8910 12400 8916
rect 12164 7744 12216 7750
rect 12164 7686 12216 7692
rect 12072 7404 12124 7410
rect 12072 7346 12124 7352
rect 11060 6928 11112 6934
rect 11060 6870 11112 6876
rect 10416 6792 10468 6798
rect 10416 6734 10468 6740
rect 10692 6792 10744 6798
rect 10692 6734 10744 6740
rect 10876 6792 10928 6798
rect 10876 6734 10928 6740
rect 11072 6662 11100 6870
rect 10232 6656 10284 6662
rect 10232 6598 10284 6604
rect 10416 6656 10468 6662
rect 10416 6598 10468 6604
rect 11060 6656 11112 6662
rect 11060 6598 11112 6604
rect 10048 6316 10100 6322
rect 10048 6258 10100 6264
rect 9956 6180 10008 6186
rect 9956 6122 10008 6128
rect 9772 5772 9824 5778
rect 9772 5714 9824 5720
rect 8760 5704 8812 5710
rect 8760 5646 8812 5652
rect 9588 5704 9640 5710
rect 9588 5646 9640 5652
rect 8392 5636 8444 5642
rect 8392 5578 8444 5584
rect 8772 5234 8800 5646
rect 9036 5636 9088 5642
rect 9036 5578 9088 5584
rect 7932 5228 7984 5234
rect 7932 5170 7984 5176
rect 8760 5228 8812 5234
rect 8760 5170 8812 5176
rect 8484 5024 8536 5030
rect 8484 4966 8536 4972
rect 7656 4820 7708 4826
rect 7656 4762 7708 4768
rect 7472 4616 7524 4622
rect 7472 4558 7524 4564
rect 7668 4554 7696 4762
rect 8496 4554 8524 4966
rect 7656 4548 7708 4554
rect 7656 4490 7708 4496
rect 8484 4548 8536 4554
rect 8484 4490 8536 4496
rect 8024 4480 8076 4486
rect 8024 4422 8076 4428
rect 6552 4276 6604 4282
rect 6552 4218 6604 4224
rect 8036 4214 8064 4422
rect 8024 4208 8076 4214
rect 8024 4150 8076 4156
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 9048 3534 9076 5578
rect 9784 5234 9812 5714
rect 9772 5228 9824 5234
rect 9772 5170 9824 5176
rect 9588 4684 9640 4690
rect 9588 4626 9640 4632
rect 9600 4554 9628 4626
rect 9588 4548 9640 4554
rect 9588 4490 9640 4496
rect 9496 4480 9548 4486
rect 9496 4422 9548 4428
rect 9508 3534 9536 4422
rect 9968 4282 9996 6122
rect 10244 5846 10272 6598
rect 10428 6254 10456 6598
rect 12084 6390 12112 7346
rect 12176 6934 12204 7686
rect 12164 6928 12216 6934
rect 12164 6870 12216 6876
rect 12072 6384 12124 6390
rect 12072 6326 12124 6332
rect 11980 6316 12032 6322
rect 11980 6258 12032 6264
rect 10416 6248 10468 6254
rect 10416 6190 10468 6196
rect 11888 6248 11940 6254
rect 11888 6190 11940 6196
rect 11796 6112 11848 6118
rect 11796 6054 11848 6060
rect 11808 5846 11836 6054
rect 10232 5840 10284 5846
rect 10232 5782 10284 5788
rect 10968 5840 11020 5846
rect 10968 5782 11020 5788
rect 11796 5840 11848 5846
rect 11796 5782 11848 5788
rect 10508 5364 10560 5370
rect 10508 5306 10560 5312
rect 10520 4622 10548 5306
rect 10692 4820 10744 4826
rect 10692 4762 10744 4768
rect 10704 4622 10732 4762
rect 10980 4758 11008 5782
rect 11900 5710 11928 6190
rect 11992 5914 12020 6258
rect 11980 5908 12032 5914
rect 11980 5850 12032 5856
rect 12176 5846 12204 6870
rect 12360 6798 12388 8910
rect 12452 8022 12480 10610
rect 12544 8956 12572 11086
rect 12636 10674 12664 11154
rect 12716 11008 12768 11014
rect 12716 10950 12768 10956
rect 12728 10674 12756 10950
rect 12624 10668 12676 10674
rect 12624 10610 12676 10616
rect 12716 10668 12768 10674
rect 12716 10610 12768 10616
rect 13004 10538 13032 11154
rect 14844 11150 14872 12406
rect 15304 12238 15332 12582
rect 15488 12306 15516 15438
rect 15580 15434 15608 16526
rect 15660 16448 15712 16454
rect 15660 16390 15712 16396
rect 15568 15428 15620 15434
rect 15568 15370 15620 15376
rect 15580 14890 15608 15370
rect 15672 15366 15700 16390
rect 15844 16108 15896 16114
rect 16408 16096 16436 18935
rect 17052 18714 17080 19207
rect 18340 18766 18368 19722
rect 18708 19378 18736 19858
rect 18696 19372 18748 19378
rect 18696 19314 18748 19320
rect 18696 19236 18748 19242
rect 18696 19178 18748 19184
rect 18708 18766 18736 19178
rect 18328 18760 18380 18766
rect 17052 18686 17172 18714
rect 18328 18702 18380 18708
rect 18420 18760 18472 18766
rect 18420 18702 18472 18708
rect 18696 18760 18748 18766
rect 18696 18702 18748 18708
rect 17040 18624 17092 18630
rect 17040 18566 17092 18572
rect 16764 18284 16816 18290
rect 16764 18226 16816 18232
rect 16776 17882 16804 18226
rect 16764 17876 16816 17882
rect 16764 17818 16816 17824
rect 17052 17678 17080 18566
rect 17144 17678 17172 18686
rect 18052 18216 18104 18222
rect 18052 18158 18104 18164
rect 17684 18148 17736 18154
rect 17684 18090 17736 18096
rect 17696 17678 17724 18090
rect 17960 18080 18012 18086
rect 17960 18022 18012 18028
rect 17040 17672 17092 17678
rect 17040 17614 17092 17620
rect 17132 17672 17184 17678
rect 17132 17614 17184 17620
rect 17592 17672 17644 17678
rect 17592 17614 17644 17620
rect 17684 17672 17736 17678
rect 17684 17614 17736 17620
rect 17868 17672 17920 17678
rect 17868 17614 17920 17620
rect 16670 17368 16726 17377
rect 16670 17303 16726 17312
rect 16684 17270 16712 17303
rect 17144 17270 17172 17614
rect 17408 17604 17460 17610
rect 17408 17546 17460 17552
rect 17420 17338 17448 17546
rect 17604 17338 17632 17614
rect 17408 17332 17460 17338
rect 17408 17274 17460 17280
rect 17592 17332 17644 17338
rect 17592 17274 17644 17280
rect 16672 17264 16724 17270
rect 16672 17206 16724 17212
rect 17132 17264 17184 17270
rect 17132 17206 17184 17212
rect 15844 16050 15896 16056
rect 16224 16068 16436 16096
rect 15752 15632 15804 15638
rect 15752 15574 15804 15580
rect 15660 15360 15712 15366
rect 15660 15302 15712 15308
rect 15672 15026 15700 15302
rect 15764 15026 15792 15574
rect 15856 15162 15884 16050
rect 15844 15156 15896 15162
rect 15844 15098 15896 15104
rect 15660 15020 15712 15026
rect 15660 14962 15712 14968
rect 15752 15020 15804 15026
rect 15752 14962 15804 14968
rect 15568 14884 15620 14890
rect 15568 14826 15620 14832
rect 15844 14816 15896 14822
rect 15844 14758 15896 14764
rect 16028 14816 16080 14822
rect 16028 14758 16080 14764
rect 15856 14414 15884 14758
rect 16040 14618 16068 14758
rect 16028 14612 16080 14618
rect 16028 14554 16080 14560
rect 15844 14408 15896 14414
rect 15844 14350 15896 14356
rect 15856 13734 15884 14350
rect 16028 14272 16080 14278
rect 16028 14214 16080 14220
rect 15844 13728 15896 13734
rect 15844 13670 15896 13676
rect 16040 13394 16068 14214
rect 16028 13388 16080 13394
rect 16028 13330 16080 13336
rect 15752 13252 15804 13258
rect 15752 13194 15804 13200
rect 15764 12986 15792 13194
rect 15752 12980 15804 12986
rect 15752 12922 15804 12928
rect 15660 12912 15712 12918
rect 15658 12880 15660 12889
rect 15712 12880 15714 12889
rect 15658 12815 15714 12824
rect 16120 12776 16172 12782
rect 16120 12718 16172 12724
rect 16132 12442 16160 12718
rect 16120 12436 16172 12442
rect 16120 12378 16172 12384
rect 15476 12300 15528 12306
rect 15476 12242 15528 12248
rect 15292 12232 15344 12238
rect 15292 12174 15344 12180
rect 15476 11280 15528 11286
rect 15476 11222 15528 11228
rect 14924 11212 14976 11218
rect 14924 11154 14976 11160
rect 14188 11144 14240 11150
rect 14188 11086 14240 11092
rect 14832 11144 14884 11150
rect 14832 11086 14884 11092
rect 13912 11008 13964 11014
rect 13912 10950 13964 10956
rect 12992 10532 13044 10538
rect 12992 10474 13044 10480
rect 13924 10062 13952 10950
rect 13912 10056 13964 10062
rect 13912 9998 13964 10004
rect 13924 9586 13952 9998
rect 14096 9920 14148 9926
rect 14096 9862 14148 9868
rect 12808 9580 12860 9586
rect 12808 9522 12860 9528
rect 13912 9580 13964 9586
rect 13912 9522 13964 9528
rect 12820 9178 12848 9522
rect 13636 9444 13688 9450
rect 13636 9386 13688 9392
rect 12808 9172 12860 9178
rect 12808 9114 12860 9120
rect 13648 9042 13676 9386
rect 13636 9036 13688 9042
rect 13636 8978 13688 8984
rect 13820 9036 13872 9042
rect 13820 8978 13872 8984
rect 12624 8968 12676 8974
rect 12544 8928 12624 8956
rect 12624 8910 12676 8916
rect 12636 8498 12664 8910
rect 12624 8492 12676 8498
rect 12624 8434 12676 8440
rect 12900 8084 12952 8090
rect 12900 8026 12952 8032
rect 13176 8084 13228 8090
rect 13176 8026 13228 8032
rect 12440 8016 12492 8022
rect 12440 7958 12492 7964
rect 12912 7886 12940 8026
rect 12900 7880 12952 7886
rect 12530 7848 12586 7857
rect 12900 7822 12952 7828
rect 12530 7783 12532 7792
rect 12584 7783 12586 7792
rect 12532 7754 12584 7760
rect 12912 7342 12940 7822
rect 12992 7472 13044 7478
rect 12992 7414 13044 7420
rect 12900 7336 12952 7342
rect 12900 7278 12952 7284
rect 12716 7268 12768 7274
rect 12716 7210 12768 7216
rect 12348 6792 12400 6798
rect 12348 6734 12400 6740
rect 12624 6316 12676 6322
rect 12624 6258 12676 6264
rect 12636 5914 12664 6258
rect 12728 5914 12756 7210
rect 13004 6458 13032 7414
rect 13188 7410 13216 8026
rect 13452 7948 13504 7954
rect 13452 7890 13504 7896
rect 13268 7812 13320 7818
rect 13268 7754 13320 7760
rect 13280 7410 13308 7754
rect 13176 7404 13228 7410
rect 13176 7346 13228 7352
rect 13268 7404 13320 7410
rect 13268 7346 13320 7352
rect 13464 7342 13492 7890
rect 13648 7886 13676 8978
rect 13636 7880 13688 7886
rect 13636 7822 13688 7828
rect 13648 7410 13676 7822
rect 13728 7812 13780 7818
rect 13728 7754 13780 7760
rect 13544 7404 13596 7410
rect 13544 7346 13596 7352
rect 13636 7404 13688 7410
rect 13636 7346 13688 7352
rect 13452 7336 13504 7342
rect 13452 7278 13504 7284
rect 13268 7268 13320 7274
rect 13268 7210 13320 7216
rect 13176 7200 13228 7206
rect 13176 7142 13228 7148
rect 12992 6452 13044 6458
rect 12992 6394 13044 6400
rect 13004 6322 13032 6394
rect 13188 6322 13216 7142
rect 13280 6934 13308 7210
rect 13268 6928 13320 6934
rect 13268 6870 13320 6876
rect 13280 6322 13308 6870
rect 12992 6316 13044 6322
rect 12992 6258 13044 6264
rect 13176 6316 13228 6322
rect 13176 6258 13228 6264
rect 13268 6316 13320 6322
rect 13268 6258 13320 6264
rect 13084 6180 13136 6186
rect 13084 6122 13136 6128
rect 12808 6112 12860 6118
rect 12808 6054 12860 6060
rect 12900 6112 12952 6118
rect 12900 6054 12952 6060
rect 12624 5908 12676 5914
rect 12624 5850 12676 5856
rect 12716 5908 12768 5914
rect 12716 5850 12768 5856
rect 12164 5840 12216 5846
rect 12164 5782 12216 5788
rect 12532 5772 12584 5778
rect 12532 5714 12584 5720
rect 11888 5704 11940 5710
rect 11888 5646 11940 5652
rect 12348 5704 12400 5710
rect 12348 5646 12400 5652
rect 11888 5568 11940 5574
rect 11888 5510 11940 5516
rect 11900 5370 11928 5510
rect 11796 5364 11848 5370
rect 11796 5306 11848 5312
rect 11888 5364 11940 5370
rect 11888 5306 11940 5312
rect 12072 5364 12124 5370
rect 12072 5306 12124 5312
rect 11704 5228 11756 5234
rect 11704 5170 11756 5176
rect 11060 5092 11112 5098
rect 11060 5034 11112 5040
rect 10968 4752 11020 4758
rect 10968 4694 11020 4700
rect 10508 4616 10560 4622
rect 10508 4558 10560 4564
rect 10692 4616 10744 4622
rect 10692 4558 10744 4564
rect 9956 4276 10008 4282
rect 9956 4218 10008 4224
rect 9968 4146 9996 4218
rect 10232 4208 10284 4214
rect 10232 4150 10284 4156
rect 9956 4140 10008 4146
rect 9956 4082 10008 4088
rect 9036 3528 9088 3534
rect 9036 3470 9088 3476
rect 9496 3528 9548 3534
rect 9496 3470 9548 3476
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 9968 3058 9996 4082
rect 10140 3732 10192 3738
rect 10140 3674 10192 3680
rect 10152 3194 10180 3674
rect 10140 3188 10192 3194
rect 10140 3130 10192 3136
rect 10244 3058 10272 4150
rect 10416 4004 10468 4010
rect 10416 3946 10468 3952
rect 10428 3602 10456 3946
rect 10704 3942 10732 4558
rect 11072 4264 11100 5034
rect 11520 5024 11572 5030
rect 11520 4966 11572 4972
rect 11532 4486 11560 4966
rect 11152 4480 11204 4486
rect 11152 4422 11204 4428
rect 11520 4480 11572 4486
rect 11520 4422 11572 4428
rect 10796 4236 11100 4264
rect 10796 4146 10824 4236
rect 10784 4140 10836 4146
rect 10784 4082 10836 4088
rect 10876 4140 10928 4146
rect 10876 4082 10928 4088
rect 10508 3936 10560 3942
rect 10508 3878 10560 3884
rect 10692 3936 10744 3942
rect 10692 3878 10744 3884
rect 10416 3596 10468 3602
rect 10416 3538 10468 3544
rect 10520 3126 10548 3878
rect 10888 3398 10916 4082
rect 10876 3392 10928 3398
rect 10876 3334 10928 3340
rect 10508 3120 10560 3126
rect 10508 3062 10560 3068
rect 10888 3058 10916 3334
rect 11072 3074 11100 4236
rect 11164 4146 11192 4422
rect 11716 4282 11744 5170
rect 11704 4276 11756 4282
rect 11704 4218 11756 4224
rect 11612 4208 11664 4214
rect 11612 4150 11664 4156
rect 11152 4140 11204 4146
rect 11152 4082 11204 4088
rect 11164 4026 11192 4082
rect 11428 4072 11480 4078
rect 11164 3998 11284 4026
rect 11428 4014 11480 4020
rect 11256 3534 11284 3998
rect 11440 3534 11468 4014
rect 11244 3528 11296 3534
rect 11244 3470 11296 3476
rect 11428 3528 11480 3534
rect 11428 3470 11480 3476
rect 11152 3460 11204 3466
rect 11152 3402 11204 3408
rect 11164 3194 11192 3402
rect 11152 3188 11204 3194
rect 11152 3130 11204 3136
rect 11624 3126 11652 4150
rect 11808 3942 11836 5306
rect 12084 5234 12112 5306
rect 12072 5228 12124 5234
rect 12072 5170 12124 5176
rect 11888 5024 11940 5030
rect 11888 4966 11940 4972
rect 11796 3936 11848 3942
rect 11796 3878 11848 3884
rect 11612 3120 11664 3126
rect 11072 3058 11192 3074
rect 11612 3062 11664 3068
rect 9956 3052 10008 3058
rect 9956 2994 10008 3000
rect 10232 3052 10284 3058
rect 10232 2994 10284 3000
rect 10876 3052 10928 3058
rect 11072 3052 11204 3058
rect 11072 3046 11152 3052
rect 10876 2994 10928 3000
rect 11152 2994 11204 3000
rect 848 2984 900 2990
rect 846 2952 848 2961
rect 900 2952 902 2961
rect 846 2887 902 2896
rect 9968 2854 9996 2994
rect 10416 2984 10468 2990
rect 10416 2926 10468 2932
rect 9956 2848 10008 2854
rect 9956 2790 10008 2796
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 10428 2650 10456 2926
rect 10888 2774 10916 2994
rect 11164 2774 11192 2994
rect 10888 2746 11008 2774
rect 11164 2746 11284 2774
rect 10416 2644 10468 2650
rect 10416 2586 10468 2592
rect 10980 2514 11008 2746
rect 10968 2508 11020 2514
rect 10968 2450 11020 2456
rect 11256 2446 11284 2746
rect 11624 2446 11652 3062
rect 11808 3058 11836 3878
rect 11900 3534 11928 4966
rect 12360 4690 12388 5646
rect 12544 5098 12572 5714
rect 12728 5642 12756 5850
rect 12820 5710 12848 6054
rect 12808 5704 12860 5710
rect 12808 5646 12860 5652
rect 12716 5636 12768 5642
rect 12716 5578 12768 5584
rect 12912 5234 12940 6054
rect 13096 5914 13124 6122
rect 13084 5908 13136 5914
rect 13084 5850 13136 5856
rect 13188 5846 13216 6258
rect 13176 5840 13228 5846
rect 13176 5782 13228 5788
rect 12900 5228 12952 5234
rect 12900 5170 12952 5176
rect 12532 5092 12584 5098
rect 12532 5034 12584 5040
rect 12348 4684 12400 4690
rect 12348 4626 12400 4632
rect 12808 4480 12860 4486
rect 12808 4422 12860 4428
rect 12820 4282 12848 4422
rect 13464 4282 13492 7278
rect 12808 4276 12860 4282
rect 12808 4218 12860 4224
rect 13452 4276 13504 4282
rect 13452 4218 13504 4224
rect 13268 4140 13320 4146
rect 13268 4082 13320 4088
rect 11888 3528 11940 3534
rect 11888 3470 11940 3476
rect 11796 3052 11848 3058
rect 11796 2994 11848 3000
rect 11244 2440 11296 2446
rect 11244 2382 11296 2388
rect 11612 2440 11664 2446
rect 11612 2382 11664 2388
rect 11900 2310 11928 3470
rect 13280 3466 13308 4082
rect 13556 3618 13584 7346
rect 13740 7342 13768 7754
rect 13728 7336 13780 7342
rect 13728 7278 13780 7284
rect 13740 7206 13768 7278
rect 13728 7200 13780 7206
rect 13728 7142 13780 7148
rect 13832 6458 13860 8978
rect 14108 8974 14136 9862
rect 14200 9382 14228 11086
rect 14372 10056 14424 10062
rect 14292 10016 14372 10044
rect 14188 9376 14240 9382
rect 14188 9318 14240 9324
rect 14096 8968 14148 8974
rect 14096 8910 14148 8916
rect 14200 8498 14228 9318
rect 14292 8974 14320 10016
rect 14372 9998 14424 10004
rect 14936 9994 14964 11154
rect 15108 11144 15160 11150
rect 15108 11086 15160 11092
rect 15120 10266 15148 11086
rect 15488 10674 15516 11222
rect 16120 11212 16172 11218
rect 16120 11154 16172 11160
rect 15476 10668 15528 10674
rect 15476 10610 15528 10616
rect 15384 10600 15436 10606
rect 15384 10542 15436 10548
rect 15108 10260 15160 10266
rect 15108 10202 15160 10208
rect 14924 9988 14976 9994
rect 14924 9930 14976 9936
rect 14464 9920 14516 9926
rect 14464 9862 14516 9868
rect 14476 9518 14504 9862
rect 14464 9512 14516 9518
rect 14464 9454 14516 9460
rect 14476 8974 14504 9454
rect 14280 8968 14332 8974
rect 14280 8910 14332 8916
rect 14464 8968 14516 8974
rect 14464 8910 14516 8916
rect 14188 8492 14240 8498
rect 14188 8434 14240 8440
rect 14004 8288 14056 8294
rect 14004 8230 14056 8236
rect 14016 7954 14044 8230
rect 14200 8090 14228 8434
rect 14188 8084 14240 8090
rect 14188 8026 14240 8032
rect 14292 8022 14320 8910
rect 14280 8016 14332 8022
rect 14280 7958 14332 7964
rect 14004 7948 14056 7954
rect 14004 7890 14056 7896
rect 14832 7812 14884 7818
rect 14832 7754 14884 7760
rect 14844 7478 14872 7754
rect 14936 7750 14964 9930
rect 15120 9042 15148 10202
rect 15396 10062 15424 10542
rect 15488 10266 15516 10610
rect 15476 10260 15528 10266
rect 15476 10202 15528 10208
rect 16132 10130 16160 11154
rect 16224 11082 16252 16068
rect 16396 15972 16448 15978
rect 16396 15914 16448 15920
rect 16408 15366 16436 15914
rect 16396 15360 16448 15366
rect 16396 15302 16448 15308
rect 16304 15088 16356 15094
rect 16304 15030 16356 15036
rect 16316 14006 16344 15030
rect 16408 14958 16436 15302
rect 16684 15008 16712 17206
rect 17500 17196 17552 17202
rect 17500 17138 17552 17144
rect 17132 16720 17184 16726
rect 17132 16662 17184 16668
rect 16856 16108 16908 16114
rect 16856 16050 16908 16056
rect 16868 15162 16896 16050
rect 17144 16046 17172 16662
rect 17224 16652 17276 16658
rect 17224 16594 17276 16600
rect 17236 16114 17264 16594
rect 17224 16108 17276 16114
rect 17224 16050 17276 16056
rect 17132 16040 17184 16046
rect 17132 15982 17184 15988
rect 17144 15366 17172 15982
rect 17408 15904 17460 15910
rect 17408 15846 17460 15852
rect 17420 15502 17448 15846
rect 17408 15496 17460 15502
rect 17408 15438 17460 15444
rect 17512 15484 17540 17138
rect 17696 16182 17724 17614
rect 17880 17377 17908 17614
rect 17866 17368 17922 17377
rect 17866 17303 17922 17312
rect 17972 17202 18000 18022
rect 18064 17746 18092 18158
rect 18432 17882 18460 18702
rect 18420 17876 18472 17882
rect 18420 17818 18472 17824
rect 18708 17746 18736 18702
rect 18800 18290 18828 19994
rect 18984 19786 19012 20878
rect 19616 19848 19668 19854
rect 19616 19790 19668 19796
rect 18972 19780 19024 19786
rect 18972 19722 19024 19728
rect 18984 19378 19012 19722
rect 19628 19514 19656 19790
rect 19524 19508 19576 19514
rect 19524 19450 19576 19456
rect 19616 19508 19668 19514
rect 19616 19450 19668 19456
rect 18972 19372 19024 19378
rect 18972 19314 19024 19320
rect 18880 19168 18932 19174
rect 18880 19110 18932 19116
rect 18892 18766 18920 19110
rect 18880 18760 18932 18766
rect 18880 18702 18932 18708
rect 18788 18284 18840 18290
rect 18788 18226 18840 18232
rect 18052 17740 18104 17746
rect 18052 17682 18104 17688
rect 18696 17740 18748 17746
rect 18696 17682 18748 17688
rect 18052 17332 18104 17338
rect 18052 17274 18104 17280
rect 18064 17202 18092 17274
rect 17868 17196 17920 17202
rect 17868 17138 17920 17144
rect 17960 17196 18012 17202
rect 17960 17138 18012 17144
rect 18052 17196 18104 17202
rect 18052 17138 18104 17144
rect 17684 16176 17736 16182
rect 17684 16118 17736 16124
rect 17776 15972 17828 15978
rect 17776 15914 17828 15920
rect 17684 15700 17736 15706
rect 17684 15642 17736 15648
rect 17696 15570 17724 15642
rect 17684 15564 17736 15570
rect 17684 15506 17736 15512
rect 17592 15496 17644 15502
rect 17512 15456 17592 15484
rect 17132 15360 17184 15366
rect 17132 15302 17184 15308
rect 17512 15201 17540 15456
rect 17592 15438 17644 15444
rect 17498 15192 17554 15201
rect 16856 15156 16908 15162
rect 17498 15127 17554 15136
rect 16856 15098 16908 15104
rect 17696 15094 17724 15506
rect 17788 15162 17816 15914
rect 17880 15366 17908 17138
rect 17960 17060 18012 17066
rect 17960 17002 18012 17008
rect 17972 16794 18000 17002
rect 17960 16788 18012 16794
rect 17960 16730 18012 16736
rect 18064 16590 18092 17138
rect 18052 16584 18104 16590
rect 18052 16526 18104 16532
rect 17868 15360 17920 15366
rect 17868 15302 17920 15308
rect 17776 15156 17828 15162
rect 17776 15098 17828 15104
rect 17684 15088 17736 15094
rect 17684 15030 17736 15036
rect 18800 15026 18828 18226
rect 16764 15020 16816 15026
rect 16684 14980 16764 15008
rect 16764 14962 16816 14968
rect 17960 15020 18012 15026
rect 17960 14962 18012 14968
rect 18144 15020 18196 15026
rect 18144 14962 18196 14968
rect 18236 15020 18288 15026
rect 18236 14962 18288 14968
rect 18788 15020 18840 15026
rect 18788 14962 18840 14968
rect 16396 14952 16448 14958
rect 16396 14894 16448 14900
rect 16304 14000 16356 14006
rect 16304 13942 16356 13948
rect 16304 13728 16356 13734
rect 16304 13670 16356 13676
rect 16316 13326 16344 13670
rect 16408 13530 16436 14894
rect 16672 14816 16724 14822
rect 16672 14758 16724 14764
rect 16684 14414 16712 14758
rect 16672 14408 16724 14414
rect 16672 14350 16724 14356
rect 16776 14074 16804 14962
rect 17224 14884 17276 14890
rect 17224 14826 17276 14832
rect 16764 14068 16816 14074
rect 16764 14010 16816 14016
rect 17236 13938 17264 14826
rect 17592 14340 17644 14346
rect 17592 14282 17644 14288
rect 17604 13938 17632 14282
rect 17972 14074 18000 14962
rect 18156 14618 18184 14962
rect 18144 14612 18196 14618
rect 18144 14554 18196 14560
rect 18248 14362 18276 14962
rect 18892 14822 18920 18702
rect 18984 15026 19012 19314
rect 19064 18624 19116 18630
rect 19064 18566 19116 18572
rect 19076 18358 19104 18566
rect 19536 18426 19564 19450
rect 19524 18420 19576 18426
rect 19524 18362 19576 18368
rect 19064 18352 19116 18358
rect 19064 18294 19116 18300
rect 19340 18216 19392 18222
rect 19340 18158 19392 18164
rect 19352 18034 19380 18158
rect 19260 18006 19380 18034
rect 19432 18080 19484 18086
rect 19432 18022 19484 18028
rect 19260 17814 19288 18006
rect 19248 17808 19300 17814
rect 19248 17750 19300 17756
rect 19444 16998 19472 18022
rect 19432 16992 19484 16998
rect 19432 16934 19484 16940
rect 19156 16652 19208 16658
rect 19156 16594 19208 16600
rect 19168 16250 19196 16594
rect 19720 16522 19748 21791
rect 20180 21593 20208 21830
rect 20166 21584 20222 21593
rect 20166 21519 20168 21528
rect 20220 21519 20222 21528
rect 20168 21490 20220 21496
rect 19798 21448 19854 21457
rect 19798 21383 19854 21392
rect 19812 21146 19840 21383
rect 19800 21140 19852 21146
rect 19800 21082 19852 21088
rect 20628 21140 20680 21146
rect 20628 21082 20680 21088
rect 19812 18222 19840 21082
rect 20640 20942 20668 21082
rect 19892 20936 19944 20942
rect 19892 20878 19944 20884
rect 20260 20936 20312 20942
rect 20260 20878 20312 20884
rect 20536 20936 20588 20942
rect 20536 20878 20588 20884
rect 20628 20936 20680 20942
rect 20628 20878 20680 20884
rect 19904 20466 19932 20878
rect 20272 20602 20300 20878
rect 20444 20868 20496 20874
rect 20444 20810 20496 20816
rect 20260 20596 20312 20602
rect 20260 20538 20312 20544
rect 20456 20534 20484 20810
rect 20444 20528 20496 20534
rect 20444 20470 20496 20476
rect 19892 20460 19944 20466
rect 19892 20402 19944 20408
rect 19904 19854 19932 20402
rect 20456 20058 20484 20470
rect 20548 20330 20576 20878
rect 20536 20324 20588 20330
rect 20536 20266 20588 20272
rect 20444 20052 20496 20058
rect 20444 19994 20496 20000
rect 20628 20052 20680 20058
rect 20628 19994 20680 20000
rect 19892 19848 19944 19854
rect 19892 19790 19944 19796
rect 20076 19848 20128 19854
rect 20076 19790 20128 19796
rect 19904 18698 19932 19790
rect 19984 19780 20036 19786
rect 19984 19722 20036 19728
rect 19996 19378 20024 19722
rect 20088 19378 20116 19790
rect 20640 19378 20668 19994
rect 19984 19372 20036 19378
rect 19984 19314 20036 19320
rect 20076 19372 20128 19378
rect 20076 19314 20128 19320
rect 20628 19372 20680 19378
rect 20628 19314 20680 19320
rect 20260 19168 20312 19174
rect 20260 19110 20312 19116
rect 19892 18692 19944 18698
rect 19892 18634 19944 18640
rect 19904 18222 19932 18634
rect 20272 18426 20300 19110
rect 20628 18692 20680 18698
rect 20628 18634 20680 18640
rect 20260 18420 20312 18426
rect 20260 18362 20312 18368
rect 20076 18284 20128 18290
rect 20076 18226 20128 18232
rect 19800 18216 19852 18222
rect 19800 18158 19852 18164
rect 19892 18216 19944 18222
rect 19892 18158 19944 18164
rect 19904 17678 19932 18158
rect 20088 17882 20116 18226
rect 20076 17876 20128 17882
rect 20076 17818 20128 17824
rect 19892 17672 19944 17678
rect 19892 17614 19944 17620
rect 20272 17610 20300 18362
rect 20444 18352 20496 18358
rect 20444 18294 20496 18300
rect 20456 17678 20484 18294
rect 20444 17672 20496 17678
rect 20444 17614 20496 17620
rect 20260 17604 20312 17610
rect 20260 17546 20312 17552
rect 20444 17196 20496 17202
rect 20444 17138 20496 17144
rect 20456 16794 20484 17138
rect 19984 16788 20036 16794
rect 19984 16730 20036 16736
rect 20444 16788 20496 16794
rect 20444 16730 20496 16736
rect 19996 16590 20024 16730
rect 19984 16584 20036 16590
rect 19984 16526 20036 16532
rect 20352 16584 20404 16590
rect 20352 16526 20404 16532
rect 19708 16516 19760 16522
rect 19708 16458 19760 16464
rect 19248 16448 19300 16454
rect 19248 16390 19300 16396
rect 19156 16244 19208 16250
rect 19156 16186 19208 16192
rect 19260 15638 19288 16390
rect 19248 15632 19300 15638
rect 19248 15574 19300 15580
rect 19432 15496 19484 15502
rect 19432 15438 19484 15444
rect 18972 15020 19024 15026
rect 18972 14962 19024 14968
rect 18984 14890 19012 14962
rect 19444 14890 19472 15438
rect 18972 14884 19024 14890
rect 18972 14826 19024 14832
rect 19432 14884 19484 14890
rect 19432 14826 19484 14832
rect 18420 14816 18472 14822
rect 18420 14758 18472 14764
rect 18880 14816 18932 14822
rect 18880 14758 18932 14764
rect 18432 14414 18460 14758
rect 18156 14334 18276 14362
rect 18420 14408 18472 14414
rect 18420 14350 18472 14356
rect 18604 14408 18656 14414
rect 18604 14350 18656 14356
rect 18156 14278 18184 14334
rect 18144 14272 18196 14278
rect 18144 14214 18196 14220
rect 18236 14272 18288 14278
rect 18236 14214 18288 14220
rect 17960 14068 18012 14074
rect 17960 14010 18012 14016
rect 17224 13932 17276 13938
rect 17224 13874 17276 13880
rect 17592 13932 17644 13938
rect 17592 13874 17644 13880
rect 17776 13932 17828 13938
rect 18144 13932 18196 13938
rect 17828 13892 18144 13920
rect 17776 13874 17828 13880
rect 16396 13524 16448 13530
rect 16396 13466 16448 13472
rect 16304 13320 16356 13326
rect 16304 13262 16356 13268
rect 16316 12850 16344 13262
rect 16304 12844 16356 12850
rect 16304 12786 16356 12792
rect 16408 12782 16436 13466
rect 16948 13184 17000 13190
rect 16948 13126 17000 13132
rect 16960 12850 16988 13126
rect 16948 12844 17000 12850
rect 16948 12786 17000 12792
rect 16396 12776 16448 12782
rect 16396 12718 16448 12724
rect 17236 12238 17264 13874
rect 17972 12866 18000 13892
rect 18248 13920 18276 14214
rect 18616 14074 18644 14350
rect 18880 14272 18932 14278
rect 18880 14214 18932 14220
rect 18604 14068 18656 14074
rect 18604 14010 18656 14016
rect 18196 13892 18276 13920
rect 18144 13874 18196 13880
rect 17880 12838 18276 12866
rect 18892 12850 18920 14214
rect 19340 14000 19392 14006
rect 19338 13968 19340 13977
rect 19392 13968 19394 13977
rect 19156 13932 19208 13938
rect 19338 13903 19394 13912
rect 19432 13966 19484 13972
rect 19484 13926 19564 13954
rect 19432 13908 19484 13914
rect 19156 13874 19208 13880
rect 19168 13326 19196 13874
rect 19432 13864 19484 13870
rect 19430 13832 19432 13841
rect 19484 13832 19486 13841
rect 19536 13818 19564 13926
rect 19616 13932 19668 13938
rect 19616 13874 19668 13880
rect 19340 13796 19392 13802
rect 19534 13802 19564 13818
rect 19430 13767 19486 13776
rect 19524 13796 19576 13802
rect 19340 13738 19392 13744
rect 19524 13738 19576 13744
rect 19352 13705 19380 13738
rect 19432 13728 19484 13734
rect 19338 13696 19394 13705
rect 19628 13705 19656 13874
rect 19614 13696 19670 13705
rect 19432 13670 19484 13676
rect 19338 13631 19394 13640
rect 19444 13394 19472 13670
rect 19536 13654 19614 13682
rect 19340 13388 19392 13394
rect 19340 13330 19392 13336
rect 19432 13388 19484 13394
rect 19432 13330 19484 13336
rect 19156 13320 19208 13326
rect 19156 13262 19208 13268
rect 19168 12986 19196 13262
rect 19352 13258 19380 13330
rect 19340 13252 19392 13258
rect 19340 13194 19392 13200
rect 19156 12980 19208 12986
rect 19156 12922 19208 12928
rect 19352 12918 19380 13194
rect 19536 13190 19564 13654
rect 19614 13631 19670 13640
rect 19616 13524 19668 13530
rect 19616 13466 19668 13472
rect 19524 13184 19576 13190
rect 19524 13126 19576 13132
rect 19340 12912 19392 12918
rect 19340 12854 19392 12860
rect 17880 12782 17908 12838
rect 17316 12776 17368 12782
rect 17316 12718 17368 12724
rect 17868 12776 17920 12782
rect 17868 12718 17920 12724
rect 17328 12442 17356 12718
rect 17776 12708 17828 12714
rect 17776 12650 17828 12656
rect 17316 12436 17368 12442
rect 17316 12378 17368 12384
rect 17788 12238 17816 12650
rect 18248 12238 18276 12838
rect 18880 12844 18932 12850
rect 18880 12786 18932 12792
rect 19628 12442 19656 13466
rect 19720 13410 19748 16458
rect 19892 14000 19944 14006
rect 19890 13968 19892 13977
rect 19944 13968 19946 13977
rect 19890 13903 19946 13912
rect 19798 13832 19854 13841
rect 19798 13767 19800 13776
rect 19852 13767 19854 13776
rect 19800 13738 19852 13744
rect 19720 13382 19932 13410
rect 19708 13320 19760 13326
rect 19708 13262 19760 13268
rect 19720 12918 19748 13262
rect 19708 12912 19760 12918
rect 19708 12854 19760 12860
rect 19616 12436 19668 12442
rect 19616 12378 19668 12384
rect 17224 12232 17276 12238
rect 17224 12174 17276 12180
rect 17776 12232 17828 12238
rect 17776 12174 17828 12180
rect 18236 12232 18288 12238
rect 18236 12174 18288 12180
rect 18052 11824 18104 11830
rect 18052 11766 18104 11772
rect 19248 11824 19300 11830
rect 19248 11766 19300 11772
rect 18064 11150 18092 11766
rect 18604 11756 18656 11762
rect 18604 11698 18656 11704
rect 18616 11150 18644 11698
rect 19260 11354 19288 11766
rect 19248 11348 19300 11354
rect 19248 11290 19300 11296
rect 19904 11150 19932 13382
rect 19996 11898 20024 16526
rect 20260 16516 20312 16522
rect 20260 16458 20312 16464
rect 20076 15360 20128 15366
rect 20076 15302 20128 15308
rect 20088 15026 20116 15302
rect 20168 15088 20220 15094
rect 20168 15030 20220 15036
rect 20076 15020 20128 15026
rect 20076 14962 20128 14968
rect 20180 14550 20208 15030
rect 20168 14544 20220 14550
rect 20168 14486 20220 14492
rect 20180 13938 20208 14486
rect 20168 13932 20220 13938
rect 20168 13874 20220 13880
rect 20272 13818 20300 16458
rect 20364 16454 20392 16526
rect 20352 16448 20404 16454
rect 20352 16390 20404 16396
rect 20640 15722 20668 18634
rect 20732 17202 20760 21830
rect 20824 21486 20852 23122
rect 20916 22094 20944 23258
rect 21272 22976 21324 22982
rect 21272 22918 21324 22924
rect 21284 22778 21312 22918
rect 21272 22772 21324 22778
rect 21272 22714 21324 22720
rect 22192 22636 22244 22642
rect 22192 22578 22244 22584
rect 21364 22568 21416 22574
rect 21364 22510 21416 22516
rect 22100 22568 22152 22574
rect 22100 22510 22152 22516
rect 20996 22094 21048 22098
rect 20916 22092 21048 22094
rect 20916 22066 20996 22092
rect 20996 22034 21048 22040
rect 21008 22001 21036 22034
rect 20994 21992 21050 22001
rect 20994 21927 21050 21936
rect 20812 21480 20864 21486
rect 20812 21422 20864 21428
rect 20904 21412 20956 21418
rect 20904 21354 20956 21360
rect 20812 21344 20864 21350
rect 20812 21286 20864 21292
rect 20824 20942 20852 21286
rect 20916 20942 20944 21354
rect 21376 21146 21404 22510
rect 22112 21554 22140 22510
rect 22204 21622 22232 22578
rect 22284 22092 22336 22098
rect 22284 22034 22336 22040
rect 22192 21616 22244 21622
rect 22192 21558 22244 21564
rect 22100 21548 22152 21554
rect 22100 21490 22152 21496
rect 22112 21146 22140 21490
rect 21364 21140 21416 21146
rect 21364 21082 21416 21088
rect 22100 21140 22152 21146
rect 22100 21082 22152 21088
rect 20812 20936 20864 20942
rect 20812 20878 20864 20884
rect 20904 20936 20956 20942
rect 20904 20878 20956 20884
rect 21088 20936 21140 20942
rect 21088 20878 21140 20884
rect 20996 20800 21048 20806
rect 20916 20760 20996 20788
rect 20916 19786 20944 20760
rect 20996 20742 21048 20748
rect 20904 19780 20956 19786
rect 20904 19722 20956 19728
rect 20916 19378 20944 19722
rect 21100 19718 21128 20878
rect 22008 20868 22060 20874
rect 22008 20810 22060 20816
rect 21640 20256 21692 20262
rect 21640 20198 21692 20204
rect 21088 19712 21140 19718
rect 21088 19654 21140 19660
rect 21548 19712 21600 19718
rect 21548 19654 21600 19660
rect 21100 19514 21128 19654
rect 21088 19508 21140 19514
rect 21088 19450 21140 19456
rect 20904 19372 20956 19378
rect 20904 19314 20956 19320
rect 21456 19236 21508 19242
rect 21456 19178 21508 19184
rect 21468 18766 21496 19178
rect 21456 18760 21508 18766
rect 21456 18702 21508 18708
rect 21456 18624 21508 18630
rect 21456 18566 21508 18572
rect 20812 18216 20864 18222
rect 20812 18158 20864 18164
rect 20824 17338 20852 18158
rect 20812 17332 20864 17338
rect 20812 17274 20864 17280
rect 20720 17196 20772 17202
rect 20720 17138 20772 17144
rect 20904 17196 20956 17202
rect 20904 17138 20956 17144
rect 21180 17196 21232 17202
rect 21180 17138 21232 17144
rect 20916 16726 20944 17138
rect 20996 17128 21048 17134
rect 20996 17070 21048 17076
rect 21008 16794 21036 17070
rect 21192 16998 21220 17138
rect 21180 16992 21232 16998
rect 21180 16934 21232 16940
rect 20996 16788 21048 16794
rect 20996 16730 21048 16736
rect 21088 16788 21140 16794
rect 21088 16730 21140 16736
rect 20904 16720 20956 16726
rect 20904 16662 20956 16668
rect 20720 16652 20772 16658
rect 20720 16594 20772 16600
rect 20732 16454 20760 16594
rect 20720 16448 20772 16454
rect 20720 16390 20772 16396
rect 20640 15694 20760 15722
rect 20628 15632 20680 15638
rect 20628 15574 20680 15580
rect 20352 15496 20404 15502
rect 20640 15484 20668 15574
rect 20404 15456 20668 15484
rect 20352 15438 20404 15444
rect 20364 15162 20392 15438
rect 20352 15156 20404 15162
rect 20352 15098 20404 15104
rect 20640 14822 20668 15456
rect 20732 15366 20760 15694
rect 20812 15700 20864 15706
rect 20812 15642 20864 15648
rect 20824 15502 20852 15642
rect 20812 15496 20864 15502
rect 20812 15438 20864 15444
rect 20720 15360 20772 15366
rect 20720 15302 20772 15308
rect 20628 14816 20680 14822
rect 20628 14758 20680 14764
rect 20640 14482 20668 14758
rect 20444 14476 20496 14482
rect 20444 14418 20496 14424
rect 20628 14476 20680 14482
rect 20628 14418 20680 14424
rect 20352 14340 20404 14346
rect 20352 14282 20404 14288
rect 20364 13938 20392 14282
rect 20352 13932 20404 13938
rect 20352 13874 20404 13880
rect 20088 13790 20300 13818
rect 19984 11892 20036 11898
rect 19984 11834 20036 11840
rect 17132 11144 17184 11150
rect 17132 11086 17184 11092
rect 17500 11144 17552 11150
rect 17500 11086 17552 11092
rect 17776 11144 17828 11150
rect 17776 11086 17828 11092
rect 18052 11144 18104 11150
rect 18052 11086 18104 11092
rect 18604 11144 18656 11150
rect 18604 11086 18656 11092
rect 19892 11144 19944 11150
rect 19892 11086 19944 11092
rect 16212 11076 16264 11082
rect 16212 11018 16264 11024
rect 16224 10674 16252 11018
rect 16212 10668 16264 10674
rect 16212 10610 16264 10616
rect 16488 10668 16540 10674
rect 16488 10610 16540 10616
rect 17040 10668 17092 10674
rect 17040 10610 17092 10616
rect 15568 10124 15620 10130
rect 15568 10066 15620 10072
rect 16120 10124 16172 10130
rect 16120 10066 16172 10072
rect 15200 10056 15252 10062
rect 15200 9998 15252 10004
rect 15384 10056 15436 10062
rect 15384 9998 15436 10004
rect 15212 9586 15240 9998
rect 15200 9580 15252 9586
rect 15200 9522 15252 9528
rect 15476 9580 15528 9586
rect 15476 9522 15528 9528
rect 15108 9036 15160 9042
rect 15108 8978 15160 8984
rect 15488 8634 15516 9522
rect 15580 9042 15608 10066
rect 16500 10062 16528 10610
rect 16764 10600 16816 10606
rect 16764 10542 16816 10548
rect 16776 10266 16804 10542
rect 17052 10266 17080 10610
rect 16764 10260 16816 10266
rect 16764 10202 16816 10208
rect 17040 10260 17092 10266
rect 17040 10202 17092 10208
rect 16028 10056 16080 10062
rect 16028 9998 16080 10004
rect 16488 10056 16540 10062
rect 16488 9998 16540 10004
rect 17040 10056 17092 10062
rect 17144 10044 17172 11086
rect 17316 10532 17368 10538
rect 17316 10474 17368 10480
rect 17328 10062 17356 10474
rect 17512 10470 17540 11086
rect 17788 10742 17816 11086
rect 18616 10810 18644 11086
rect 19340 11076 19392 11082
rect 19340 11018 19392 11024
rect 18604 10804 18656 10810
rect 18604 10746 18656 10752
rect 17776 10736 17828 10742
rect 17776 10678 17828 10684
rect 17960 10736 18012 10742
rect 17960 10678 18012 10684
rect 17684 10668 17736 10674
rect 17684 10610 17736 10616
rect 17500 10464 17552 10470
rect 17500 10406 17552 10412
rect 17092 10016 17172 10044
rect 17224 10056 17276 10062
rect 17040 9998 17092 10004
rect 17224 9998 17276 10004
rect 17316 10056 17368 10062
rect 17316 9998 17368 10004
rect 16040 9518 16068 9998
rect 16212 9920 16264 9926
rect 16212 9862 16264 9868
rect 16396 9920 16448 9926
rect 16396 9862 16448 9868
rect 16028 9512 16080 9518
rect 16028 9454 16080 9460
rect 15568 9036 15620 9042
rect 15568 8978 15620 8984
rect 15476 8628 15528 8634
rect 15476 8570 15528 8576
rect 16040 8566 16068 9454
rect 16224 8906 16252 9862
rect 16408 9178 16436 9862
rect 16500 9586 16528 9998
rect 17236 9722 17264 9998
rect 17224 9716 17276 9722
rect 17224 9658 17276 9664
rect 16488 9580 16540 9586
rect 16488 9522 16540 9528
rect 17328 9450 17356 9998
rect 17408 9580 17460 9586
rect 17408 9522 17460 9528
rect 17316 9444 17368 9450
rect 17316 9386 17368 9392
rect 16856 9376 16908 9382
rect 16856 9318 16908 9324
rect 16396 9172 16448 9178
rect 16396 9114 16448 9120
rect 16212 8900 16264 8906
rect 16212 8842 16264 8848
rect 16028 8560 16080 8566
rect 16028 8502 16080 8508
rect 15016 8492 15068 8498
rect 15016 8434 15068 8440
rect 14924 7744 14976 7750
rect 14924 7686 14976 7692
rect 14832 7472 14884 7478
rect 14832 7414 14884 7420
rect 14936 7342 14964 7686
rect 15028 7546 15056 8434
rect 16224 8430 16252 8842
rect 16408 8498 16436 9114
rect 16868 9042 16896 9318
rect 16856 9036 16908 9042
rect 16856 8978 16908 8984
rect 17040 8968 17092 8974
rect 17040 8910 17092 8916
rect 17052 8498 17080 8910
rect 17420 8838 17448 9522
rect 17408 8832 17460 8838
rect 17408 8774 17460 8780
rect 16396 8492 16448 8498
rect 16396 8434 16448 8440
rect 17040 8492 17092 8498
rect 17040 8434 17092 8440
rect 16212 8424 16264 8430
rect 16212 8366 16264 8372
rect 17132 8424 17184 8430
rect 17132 8366 17184 8372
rect 16304 8356 16356 8362
rect 16304 8298 16356 8304
rect 15016 7540 15068 7546
rect 15016 7482 15068 7488
rect 14924 7336 14976 7342
rect 14924 7278 14976 7284
rect 16120 7336 16172 7342
rect 16120 7278 16172 7284
rect 16132 6798 16160 7278
rect 16316 6798 16344 8298
rect 17144 8090 17172 8366
rect 17132 8084 17184 8090
rect 17132 8026 17184 8032
rect 17316 7812 17368 7818
rect 17316 7754 17368 7760
rect 17328 7410 17356 7754
rect 17224 7404 17276 7410
rect 17224 7346 17276 7352
rect 17316 7404 17368 7410
rect 17316 7346 17368 7352
rect 17040 7200 17092 7206
rect 17040 7142 17092 7148
rect 17052 6798 17080 7142
rect 15936 6792 15988 6798
rect 15936 6734 15988 6740
rect 16120 6792 16172 6798
rect 16120 6734 16172 6740
rect 16304 6792 16356 6798
rect 16304 6734 16356 6740
rect 17040 6792 17092 6798
rect 17040 6734 17092 6740
rect 15948 6458 15976 6734
rect 16120 6656 16172 6662
rect 16120 6598 16172 6604
rect 13820 6452 13872 6458
rect 13820 6394 13872 6400
rect 14832 6452 14884 6458
rect 14832 6394 14884 6400
rect 15936 6452 15988 6458
rect 15936 6394 15988 6400
rect 14372 6384 14424 6390
rect 14372 6326 14424 6332
rect 14096 6316 14148 6322
rect 14096 6258 14148 6264
rect 13728 6112 13780 6118
rect 13728 6054 13780 6060
rect 13740 5234 13768 6054
rect 14108 5710 14136 6258
rect 14384 6254 14412 6326
rect 14372 6248 14424 6254
rect 14372 6190 14424 6196
rect 14096 5704 14148 5710
rect 14096 5646 14148 5652
rect 14384 5234 14412 6190
rect 14464 6180 14516 6186
rect 14464 6122 14516 6128
rect 14476 5710 14504 6122
rect 14844 5914 14872 6394
rect 16132 6322 16160 6598
rect 16316 6458 16344 6734
rect 16856 6724 16908 6730
rect 16856 6666 16908 6672
rect 16304 6452 16356 6458
rect 16304 6394 16356 6400
rect 15200 6316 15252 6322
rect 15200 6258 15252 6264
rect 15844 6316 15896 6322
rect 15844 6258 15896 6264
rect 16120 6316 16172 6322
rect 16120 6258 16172 6264
rect 14832 5908 14884 5914
rect 14832 5850 14884 5856
rect 14464 5704 14516 5710
rect 14464 5646 14516 5652
rect 15212 5642 15240 6258
rect 15568 6112 15620 6118
rect 15568 6054 15620 6060
rect 15200 5636 15252 5642
rect 15200 5578 15252 5584
rect 13728 5228 13780 5234
rect 13728 5170 13780 5176
rect 13912 5228 13964 5234
rect 13912 5170 13964 5176
rect 14372 5228 14424 5234
rect 14372 5170 14424 5176
rect 13924 5030 13952 5170
rect 13912 5024 13964 5030
rect 13912 4966 13964 4972
rect 14004 5024 14056 5030
rect 14004 4966 14056 4972
rect 14016 4554 14044 4966
rect 15580 4622 15608 6054
rect 15856 5710 15884 6258
rect 16304 5908 16356 5914
rect 16304 5850 16356 5856
rect 15844 5704 15896 5710
rect 15844 5646 15896 5652
rect 16316 5234 16344 5850
rect 16868 5846 16896 6666
rect 16856 5840 16908 5846
rect 16856 5782 16908 5788
rect 16868 5710 16896 5782
rect 16856 5704 16908 5710
rect 16856 5646 16908 5652
rect 16672 5568 16724 5574
rect 16672 5510 16724 5516
rect 16684 5234 16712 5510
rect 17236 5234 17264 7346
rect 17420 6798 17448 8774
rect 17512 8362 17540 10406
rect 17696 10198 17724 10610
rect 17684 10192 17736 10198
rect 17684 10134 17736 10140
rect 17592 9920 17644 9926
rect 17592 9862 17644 9868
rect 17684 9920 17736 9926
rect 17684 9862 17736 9868
rect 17604 8498 17632 9862
rect 17696 9722 17724 9862
rect 17684 9716 17736 9722
rect 17684 9658 17736 9664
rect 17696 8974 17724 9658
rect 17684 8968 17736 8974
rect 17868 8968 17920 8974
rect 17684 8910 17736 8916
rect 17788 8928 17868 8956
rect 17592 8492 17644 8498
rect 17592 8434 17644 8440
rect 17500 8356 17552 8362
rect 17500 8298 17552 8304
rect 17512 7818 17540 8298
rect 17604 7886 17632 8434
rect 17592 7880 17644 7886
rect 17592 7822 17644 7828
rect 17500 7812 17552 7818
rect 17500 7754 17552 7760
rect 17408 6792 17460 6798
rect 17408 6734 17460 6740
rect 17316 5704 17368 5710
rect 17420 5692 17448 6734
rect 17512 5794 17540 7754
rect 17604 7546 17632 7822
rect 17592 7540 17644 7546
rect 17592 7482 17644 7488
rect 17512 5766 17632 5794
rect 17368 5664 17540 5692
rect 17316 5646 17368 5652
rect 17316 5568 17368 5574
rect 17314 5536 17316 5545
rect 17368 5536 17370 5545
rect 17314 5471 17370 5480
rect 16304 5228 16356 5234
rect 16304 5170 16356 5176
rect 16672 5228 16724 5234
rect 16672 5170 16724 5176
rect 17224 5228 17276 5234
rect 17224 5170 17276 5176
rect 16316 4826 16344 5170
rect 16488 5092 16540 5098
rect 16488 5034 16540 5040
rect 16304 4820 16356 4826
rect 16304 4762 16356 4768
rect 16500 4622 16528 5034
rect 15568 4616 15620 4622
rect 15568 4558 15620 4564
rect 15660 4616 15712 4622
rect 15660 4558 15712 4564
rect 16488 4616 16540 4622
rect 16488 4558 16540 4564
rect 14004 4548 14056 4554
rect 14004 4490 14056 4496
rect 14556 4276 14608 4282
rect 14556 4218 14608 4224
rect 13464 3590 13676 3618
rect 13464 3534 13492 3590
rect 13452 3528 13504 3534
rect 13452 3470 13504 3476
rect 13544 3528 13596 3534
rect 13544 3470 13596 3476
rect 13268 3460 13320 3466
rect 13268 3402 13320 3408
rect 13280 3058 13308 3402
rect 13556 3398 13584 3470
rect 13648 3448 13676 3590
rect 14568 3534 14596 4218
rect 15200 4140 15252 4146
rect 15200 4082 15252 4088
rect 15292 4140 15344 4146
rect 15292 4082 15344 4088
rect 15476 4140 15528 4146
rect 15580 4128 15608 4558
rect 15672 4146 15700 4558
rect 16212 4480 16264 4486
rect 16212 4422 16264 4428
rect 15528 4100 15608 4128
rect 15660 4140 15712 4146
rect 15476 4082 15528 4088
rect 15660 4082 15712 4088
rect 15212 3670 15240 4082
rect 15200 3664 15252 3670
rect 15200 3606 15252 3612
rect 14556 3528 14608 3534
rect 14556 3470 14608 3476
rect 13728 3460 13780 3466
rect 13648 3420 13728 3448
rect 13728 3402 13780 3408
rect 13544 3392 13596 3398
rect 13544 3334 13596 3340
rect 13268 3052 13320 3058
rect 13268 2994 13320 3000
rect 12072 2984 12124 2990
rect 12072 2926 12124 2932
rect 12084 2650 12112 2926
rect 13452 2848 13504 2854
rect 13452 2790 13504 2796
rect 12072 2644 12124 2650
rect 12072 2586 12124 2592
rect 13464 2446 13492 2790
rect 13556 2650 13584 3334
rect 15304 3126 15332 4082
rect 15384 4072 15436 4078
rect 15384 4014 15436 4020
rect 15934 4040 15990 4049
rect 15396 3670 15424 4014
rect 15934 3975 15990 3984
rect 15384 3664 15436 3670
rect 15384 3606 15436 3612
rect 15660 3528 15712 3534
rect 15660 3470 15712 3476
rect 15568 3460 15620 3466
rect 15568 3402 15620 3408
rect 15292 3120 15344 3126
rect 15292 3062 15344 3068
rect 15580 3058 15608 3402
rect 15672 3194 15700 3470
rect 15948 3194 15976 3975
rect 16224 3670 16252 4422
rect 17236 4146 17264 5170
rect 17224 4140 17276 4146
rect 17276 4100 17356 4128
rect 17224 4082 17276 4088
rect 16580 4072 16632 4078
rect 16580 4014 16632 4020
rect 16592 3942 16620 4014
rect 16580 3936 16632 3942
rect 16580 3878 16632 3884
rect 16948 3936 17000 3942
rect 16948 3878 17000 3884
rect 16304 3732 16356 3738
rect 16304 3674 16356 3680
rect 16212 3664 16264 3670
rect 16212 3606 16264 3612
rect 16028 3596 16080 3602
rect 16028 3538 16080 3544
rect 15660 3188 15712 3194
rect 15660 3130 15712 3136
rect 15936 3188 15988 3194
rect 15936 3130 15988 3136
rect 15752 3120 15804 3126
rect 15752 3062 15804 3068
rect 15200 3052 15252 3058
rect 15200 2994 15252 3000
rect 15568 3052 15620 3058
rect 15568 2994 15620 3000
rect 15660 3052 15712 3058
rect 15660 2994 15712 3000
rect 13636 2916 13688 2922
rect 13636 2858 13688 2864
rect 13544 2644 13596 2650
rect 13544 2586 13596 2592
rect 13648 2446 13676 2858
rect 15212 2582 15240 2994
rect 15580 2774 15608 2994
rect 15396 2746 15608 2774
rect 15200 2576 15252 2582
rect 15200 2518 15252 2524
rect 15396 2446 15424 2746
rect 13452 2440 13504 2446
rect 13452 2382 13504 2388
rect 13636 2440 13688 2446
rect 13636 2382 13688 2388
rect 15384 2440 15436 2446
rect 15672 2394 15700 2994
rect 15764 2582 15792 3062
rect 16040 2774 16068 3538
rect 16224 3126 16252 3606
rect 16316 3534 16344 3674
rect 16960 3602 16988 3878
rect 16948 3596 17000 3602
rect 16948 3538 17000 3544
rect 16304 3528 16356 3534
rect 16304 3470 16356 3476
rect 16396 3528 16448 3534
rect 16396 3470 16448 3476
rect 16580 3528 16632 3534
rect 16580 3470 16632 3476
rect 16212 3120 16264 3126
rect 16212 3062 16264 3068
rect 15856 2746 16068 2774
rect 15752 2576 15804 2582
rect 15752 2518 15804 2524
rect 15856 2446 15884 2746
rect 16408 2650 16436 3470
rect 16592 3194 16620 3470
rect 16580 3188 16632 3194
rect 16580 3130 16632 3136
rect 16396 2644 16448 2650
rect 16396 2586 16448 2592
rect 16960 2446 16988 3538
rect 17328 3534 17356 4100
rect 17316 3528 17368 3534
rect 17316 3470 17368 3476
rect 17132 3052 17184 3058
rect 17132 2994 17184 3000
rect 17144 2922 17172 2994
rect 17512 2990 17540 5664
rect 17604 5234 17632 5766
rect 17592 5228 17644 5234
rect 17592 5170 17644 5176
rect 17604 5030 17632 5170
rect 17592 5024 17644 5030
rect 17592 4966 17644 4972
rect 17604 4146 17632 4966
rect 17592 4140 17644 4146
rect 17592 4082 17644 4088
rect 17604 3534 17632 4082
rect 17696 4010 17724 8910
rect 17788 4214 17816 8928
rect 17972 8956 18000 10678
rect 19352 10606 19380 11018
rect 19800 11008 19852 11014
rect 19800 10950 19852 10956
rect 19708 10736 19760 10742
rect 19708 10678 19760 10684
rect 19340 10600 19392 10606
rect 19340 10542 19392 10548
rect 19524 10464 19576 10470
rect 19524 10406 19576 10412
rect 19536 10266 19564 10406
rect 19524 10260 19576 10266
rect 19524 10202 19576 10208
rect 19536 9586 19564 10202
rect 19720 10198 19748 10678
rect 19812 10674 19840 10950
rect 19800 10668 19852 10674
rect 19800 10610 19852 10616
rect 19708 10192 19760 10198
rect 19708 10134 19760 10140
rect 19720 10062 19748 10134
rect 19708 10056 19760 10062
rect 19708 9998 19760 10004
rect 19720 9654 19748 9998
rect 19708 9648 19760 9654
rect 19708 9590 19760 9596
rect 19812 9586 19840 10610
rect 19892 10600 19944 10606
rect 19892 10542 19944 10548
rect 19524 9580 19576 9586
rect 19524 9522 19576 9528
rect 19800 9580 19852 9586
rect 19800 9522 19852 9528
rect 19904 9518 19932 10542
rect 19984 10464 20036 10470
rect 19984 10406 20036 10412
rect 19996 10130 20024 10406
rect 19984 10124 20036 10130
rect 19984 10066 20036 10072
rect 19892 9512 19944 9518
rect 19892 9454 19944 9460
rect 19524 9376 19576 9382
rect 19524 9318 19576 9324
rect 17920 8928 18000 8956
rect 18144 8968 18196 8974
rect 17868 8910 17920 8916
rect 18144 8910 18196 8916
rect 17868 8832 17920 8838
rect 17868 8774 17920 8780
rect 18052 8832 18104 8838
rect 18052 8774 18104 8780
rect 17880 8430 17908 8774
rect 17868 8424 17920 8430
rect 17868 8366 17920 8372
rect 18064 7886 18092 8774
rect 18156 8566 18184 8910
rect 19536 8906 19564 9318
rect 19524 8900 19576 8906
rect 19524 8842 19576 8848
rect 18144 8560 18196 8566
rect 18144 8502 18196 8508
rect 19536 8498 19564 8842
rect 19708 8832 19760 8838
rect 19708 8774 19760 8780
rect 19524 8492 19576 8498
rect 19524 8434 19576 8440
rect 18052 7880 18104 7886
rect 17972 7840 18052 7868
rect 17868 7404 17920 7410
rect 17972 7392 18000 7840
rect 18052 7822 18104 7828
rect 19616 7880 19668 7886
rect 19616 7822 19668 7828
rect 18052 7744 18104 7750
rect 18052 7686 18104 7692
rect 17920 7364 18000 7392
rect 17868 7346 17920 7352
rect 18064 7342 18092 7686
rect 19628 7546 19656 7822
rect 19616 7540 19668 7546
rect 19616 7482 19668 7488
rect 18052 7336 18104 7342
rect 18052 7278 18104 7284
rect 19628 6798 19656 7482
rect 18604 6792 18656 6798
rect 18604 6734 18656 6740
rect 19616 6792 19668 6798
rect 19616 6734 19668 6740
rect 18616 6322 18644 6734
rect 18696 6724 18748 6730
rect 18696 6666 18748 6672
rect 18708 6390 18736 6666
rect 18696 6384 18748 6390
rect 18696 6326 18748 6332
rect 18420 6316 18472 6322
rect 18420 6258 18472 6264
rect 18604 6316 18656 6322
rect 18604 6258 18656 6264
rect 18328 6248 18380 6254
rect 18328 6190 18380 6196
rect 17960 5704 18012 5710
rect 17960 5646 18012 5652
rect 17972 5545 18000 5646
rect 18052 5568 18104 5574
rect 17958 5536 18014 5545
rect 18052 5510 18104 5516
rect 17958 5471 18014 5480
rect 17972 5370 18000 5471
rect 17960 5364 18012 5370
rect 17960 5306 18012 5312
rect 18064 5234 18092 5510
rect 18052 5228 18104 5234
rect 18052 5170 18104 5176
rect 18340 5098 18368 6190
rect 18432 5914 18460 6258
rect 18420 5908 18472 5914
rect 18420 5850 18472 5856
rect 18616 5642 18644 6258
rect 18708 5846 18736 6326
rect 18696 5840 18748 5846
rect 18696 5782 18748 5788
rect 18604 5636 18656 5642
rect 18604 5578 18656 5584
rect 18708 5370 18736 5782
rect 18696 5364 18748 5370
rect 18696 5306 18748 5312
rect 18328 5092 18380 5098
rect 18328 5034 18380 5040
rect 18340 4690 18368 5034
rect 18328 4684 18380 4690
rect 18328 4626 18380 4632
rect 17776 4208 17828 4214
rect 17776 4150 17828 4156
rect 19720 4146 19748 8774
rect 19800 8288 19852 8294
rect 19800 8230 19852 8236
rect 19812 7886 19840 8230
rect 19800 7880 19852 7886
rect 19852 7840 19932 7868
rect 19800 7822 19852 7828
rect 19800 7404 19852 7410
rect 19800 7346 19852 7352
rect 19812 6662 19840 7346
rect 19904 6798 19932 7840
rect 19984 7744 20036 7750
rect 19984 7686 20036 7692
rect 19996 7410 20024 7686
rect 19984 7404 20036 7410
rect 19984 7346 20036 7352
rect 19892 6792 19944 6798
rect 19892 6734 19944 6740
rect 19800 6656 19852 6662
rect 19800 6598 19852 6604
rect 19892 5636 19944 5642
rect 19892 5578 19944 5584
rect 19904 5370 19932 5578
rect 19892 5364 19944 5370
rect 19892 5306 19944 5312
rect 19800 5228 19852 5234
rect 19800 5170 19852 5176
rect 19984 5228 20036 5234
rect 19984 5170 20036 5176
rect 19812 4826 19840 5170
rect 19996 5098 20024 5170
rect 19984 5092 20036 5098
rect 19984 5034 20036 5040
rect 19800 4820 19852 4826
rect 19800 4762 19852 4768
rect 19800 4276 19852 4282
rect 19800 4218 19852 4224
rect 19708 4140 19760 4146
rect 19708 4082 19760 4088
rect 17684 4004 17736 4010
rect 17684 3946 17736 3952
rect 19812 3738 19840 4218
rect 19996 4049 20024 5034
rect 20088 4622 20116 13790
rect 20168 13728 20220 13734
rect 20168 13670 20220 13676
rect 20180 13258 20208 13670
rect 20260 13388 20312 13394
rect 20260 13330 20312 13336
rect 20352 13388 20404 13394
rect 20352 13330 20404 13336
rect 20168 13252 20220 13258
rect 20168 13194 20220 13200
rect 20272 12850 20300 13330
rect 20364 12986 20392 13330
rect 20352 12980 20404 12986
rect 20352 12922 20404 12928
rect 20260 12844 20312 12850
rect 20260 12786 20312 12792
rect 20456 12646 20484 14418
rect 20732 14362 20760 15302
rect 20640 14334 20760 14362
rect 20640 13462 20668 14334
rect 20824 14278 20852 15438
rect 20904 15020 20956 15026
rect 20904 14962 20956 14968
rect 20996 15020 21048 15026
rect 20996 14962 21048 14968
rect 20916 14414 20944 14962
rect 21008 14929 21036 14962
rect 20994 14920 21050 14929
rect 20994 14855 21050 14864
rect 20904 14408 20956 14414
rect 20904 14350 20956 14356
rect 20812 14272 20864 14278
rect 20812 14214 20864 14220
rect 20720 14068 20772 14074
rect 20720 14010 20772 14016
rect 20996 14068 21048 14074
rect 20996 14010 21048 14016
rect 20628 13456 20680 13462
rect 20628 13398 20680 13404
rect 20628 13252 20680 13258
rect 20628 13194 20680 13200
rect 20536 13184 20588 13190
rect 20536 13126 20588 13132
rect 20548 12782 20576 13126
rect 20536 12776 20588 12782
rect 20536 12718 20588 12724
rect 20640 12714 20668 13194
rect 20732 12986 20760 14010
rect 21008 13326 21036 14010
rect 20996 13320 21048 13326
rect 20996 13262 21048 13268
rect 20720 12980 20772 12986
rect 20720 12922 20772 12928
rect 20628 12708 20680 12714
rect 20628 12650 20680 12656
rect 20444 12640 20496 12646
rect 20444 12582 20496 12588
rect 20640 12442 20668 12650
rect 20628 12436 20680 12442
rect 20628 12378 20680 12384
rect 20536 11756 20588 11762
rect 20536 11698 20588 11704
rect 20352 10804 20404 10810
rect 20352 10746 20404 10752
rect 20364 10062 20392 10746
rect 20548 10674 20576 11698
rect 20904 11688 20956 11694
rect 20904 11630 20956 11636
rect 20916 10810 20944 11630
rect 20904 10804 20956 10810
rect 20904 10746 20956 10752
rect 21100 10674 21128 16730
rect 21192 16658 21220 16934
rect 21180 16652 21232 16658
rect 21180 16594 21232 16600
rect 21364 16584 21416 16590
rect 21364 16526 21416 16532
rect 21272 15496 21324 15502
rect 21272 15438 21324 15444
rect 21180 15428 21232 15434
rect 21180 15370 21232 15376
rect 21192 15026 21220 15370
rect 21284 15026 21312 15438
rect 21180 15020 21232 15026
rect 21180 14962 21232 14968
rect 21272 15020 21324 15026
rect 21272 14962 21324 14968
rect 21192 14618 21220 14962
rect 21180 14612 21232 14618
rect 21180 14554 21232 14560
rect 21180 14272 21232 14278
rect 21180 14214 21232 14220
rect 21192 13938 21220 14214
rect 21180 13932 21232 13938
rect 21180 13874 21232 13880
rect 21192 13530 21220 13874
rect 21272 13728 21324 13734
rect 21272 13670 21324 13676
rect 21180 13524 21232 13530
rect 21180 13466 21232 13472
rect 21284 13462 21312 13670
rect 21272 13456 21324 13462
rect 21272 13398 21324 13404
rect 21180 11076 21232 11082
rect 21180 11018 21232 11024
rect 20536 10668 20588 10674
rect 20536 10610 20588 10616
rect 21088 10668 21140 10674
rect 21088 10610 21140 10616
rect 20444 10464 20496 10470
rect 20444 10406 20496 10412
rect 20628 10464 20680 10470
rect 20628 10406 20680 10412
rect 20456 10062 20484 10406
rect 20640 10130 20668 10406
rect 21100 10198 21128 10610
rect 21192 10606 21220 11018
rect 21180 10600 21232 10606
rect 21180 10542 21232 10548
rect 21088 10192 21140 10198
rect 21088 10134 21140 10140
rect 20628 10124 20680 10130
rect 20628 10066 20680 10072
rect 20168 10056 20220 10062
rect 20168 9998 20220 10004
rect 20352 10056 20404 10062
rect 20352 9998 20404 10004
rect 20444 10056 20496 10062
rect 20444 9998 20496 10004
rect 21088 10056 21140 10062
rect 21088 9998 21140 10004
rect 20180 9178 20208 9998
rect 20168 9172 20220 9178
rect 20168 9114 20220 9120
rect 20076 4616 20128 4622
rect 20076 4558 20128 4564
rect 20088 4282 20116 4558
rect 20076 4276 20128 4282
rect 20076 4218 20128 4224
rect 20076 4140 20128 4146
rect 20076 4082 20128 4088
rect 19982 4040 20038 4049
rect 19982 3975 20038 3984
rect 18880 3732 18932 3738
rect 18880 3674 18932 3680
rect 19800 3732 19852 3738
rect 19800 3674 19852 3680
rect 18420 3596 18472 3602
rect 18420 3538 18472 3544
rect 17592 3528 17644 3534
rect 17592 3470 17644 3476
rect 18236 3528 18288 3534
rect 18236 3470 18288 3476
rect 18248 3058 18276 3470
rect 18432 3058 18460 3538
rect 18892 3058 18920 3674
rect 20088 3534 20116 4082
rect 20076 3528 20128 3534
rect 20076 3470 20128 3476
rect 20088 3194 20116 3470
rect 20180 3194 20208 9114
rect 20260 8968 20312 8974
rect 20260 8910 20312 8916
rect 20272 8634 20300 8910
rect 20364 8838 20392 9998
rect 21100 9874 21128 9998
rect 21192 9994 21220 10542
rect 21272 10260 21324 10266
rect 21272 10202 21324 10208
rect 21284 10062 21312 10202
rect 21272 10056 21324 10062
rect 21272 9998 21324 10004
rect 21376 9994 21404 16526
rect 21468 15502 21496 18566
rect 21560 15502 21588 19654
rect 21652 19310 21680 20198
rect 21732 19848 21784 19854
rect 21732 19790 21784 19796
rect 21916 19848 21968 19854
rect 21916 19790 21968 19796
rect 21640 19304 21692 19310
rect 21640 19246 21692 19252
rect 21652 18970 21680 19246
rect 21640 18964 21692 18970
rect 21640 18906 21692 18912
rect 21744 18766 21772 19790
rect 21928 19174 21956 19790
rect 21916 19168 21968 19174
rect 21916 19110 21968 19116
rect 21732 18760 21784 18766
rect 21732 18702 21784 18708
rect 21928 18358 21956 19110
rect 21916 18352 21968 18358
rect 21916 18294 21968 18300
rect 21824 18284 21876 18290
rect 21824 18226 21876 18232
rect 21836 17338 21864 18226
rect 21824 17332 21876 17338
rect 21824 17274 21876 17280
rect 21640 17196 21692 17202
rect 21640 17138 21692 17144
rect 21652 16726 21680 17138
rect 21640 16720 21692 16726
rect 21640 16662 21692 16668
rect 21916 16584 21968 16590
rect 21916 16526 21968 16532
rect 21824 16244 21876 16250
rect 21824 16186 21876 16192
rect 21640 15700 21692 15706
rect 21640 15642 21692 15648
rect 21456 15496 21508 15502
rect 21456 15438 21508 15444
rect 21548 15496 21600 15502
rect 21548 15438 21600 15444
rect 21468 13938 21496 15438
rect 21560 14074 21588 15438
rect 21652 15026 21680 15642
rect 21836 15026 21864 16186
rect 21640 15020 21692 15026
rect 21640 14962 21692 14968
rect 21824 15020 21876 15026
rect 21824 14962 21876 14968
rect 21732 14408 21784 14414
rect 21732 14350 21784 14356
rect 21548 14068 21600 14074
rect 21548 14010 21600 14016
rect 21456 13932 21508 13938
rect 21456 13874 21508 13880
rect 21468 13326 21496 13874
rect 21456 13320 21508 13326
rect 21456 13262 21508 13268
rect 21744 12442 21772 14350
rect 21836 12850 21864 14962
rect 21824 12844 21876 12850
rect 21824 12786 21876 12792
rect 21732 12436 21784 12442
rect 21928 12434 21956 16526
rect 22020 15706 22048 20810
rect 22192 17536 22244 17542
rect 22192 17478 22244 17484
rect 22204 17338 22232 17478
rect 22296 17338 22324 22034
rect 22572 21690 22784 21706
rect 22560 21684 22796 21690
rect 22612 21678 22744 21684
rect 22560 21626 22612 21632
rect 22744 21626 22796 21632
rect 23020 21616 23072 21622
rect 23020 21558 23072 21564
rect 22652 21548 22704 21554
rect 22652 21490 22704 21496
rect 22744 21548 22796 21554
rect 22744 21490 22796 21496
rect 22376 21480 22428 21486
rect 22376 21422 22428 21428
rect 22468 21480 22520 21486
rect 22468 21422 22520 21428
rect 22388 20806 22416 21422
rect 22480 21078 22508 21422
rect 22664 21146 22692 21490
rect 22652 21140 22704 21146
rect 22652 21082 22704 21088
rect 22468 21072 22520 21078
rect 22468 21014 22520 21020
rect 22376 20800 22428 20806
rect 22376 20742 22428 20748
rect 22388 19786 22416 20742
rect 22480 20058 22508 21014
rect 22756 20806 22784 21490
rect 22836 21140 22888 21146
rect 22836 21082 22888 21088
rect 22848 20942 22876 21082
rect 22836 20936 22888 20942
rect 22836 20878 22888 20884
rect 22744 20800 22796 20806
rect 22744 20742 22796 20748
rect 22468 20052 22520 20058
rect 22468 19994 22520 20000
rect 22480 19922 22508 19994
rect 22468 19916 22520 19922
rect 22468 19858 22520 19864
rect 22376 19780 22428 19786
rect 22376 19722 22428 19728
rect 22848 18970 22876 20878
rect 22836 18964 22888 18970
rect 22836 18906 22888 18912
rect 22652 18692 22704 18698
rect 22652 18634 22704 18640
rect 22836 18692 22888 18698
rect 22836 18634 22888 18640
rect 22376 18284 22428 18290
rect 22376 18226 22428 18232
rect 22192 17332 22244 17338
rect 22192 17274 22244 17280
rect 22284 17332 22336 17338
rect 22284 17274 22336 17280
rect 22388 17202 22416 18226
rect 22664 17678 22692 18634
rect 22848 18290 22876 18634
rect 22836 18284 22888 18290
rect 22836 18226 22888 18232
rect 22848 17882 22876 18226
rect 22836 17876 22888 17882
rect 22836 17818 22888 17824
rect 22652 17672 22704 17678
rect 22652 17614 22704 17620
rect 22848 17338 22876 17818
rect 23032 17678 23060 21558
rect 23388 21548 23440 21554
rect 23388 21490 23440 21496
rect 23204 21480 23256 21486
rect 23204 21422 23256 21428
rect 23216 19854 23244 21422
rect 23296 21140 23348 21146
rect 23296 21082 23348 21088
rect 23308 20874 23336 21082
rect 23400 20942 23428 21490
rect 23388 20936 23440 20942
rect 23388 20878 23440 20884
rect 25320 20936 25372 20942
rect 25320 20878 25372 20884
rect 23296 20868 23348 20874
rect 23296 20810 23348 20816
rect 24216 20392 24268 20398
rect 24216 20334 24268 20340
rect 24228 20058 24256 20334
rect 24400 20324 24452 20330
rect 24400 20266 24452 20272
rect 24032 20052 24084 20058
rect 24032 19994 24084 20000
rect 24216 20052 24268 20058
rect 24216 19994 24268 20000
rect 23204 19848 23256 19854
rect 23480 19848 23532 19854
rect 23256 19808 23336 19836
rect 23204 19790 23256 19796
rect 23112 19168 23164 19174
rect 23112 19110 23164 19116
rect 23124 18970 23152 19110
rect 23112 18964 23164 18970
rect 23112 18906 23164 18912
rect 23020 17672 23072 17678
rect 23020 17614 23072 17620
rect 23308 17610 23336 19808
rect 23400 19808 23480 19836
rect 23400 19446 23428 19808
rect 23480 19790 23532 19796
rect 23848 19780 23900 19786
rect 23848 19722 23900 19728
rect 23664 19712 23716 19718
rect 23664 19654 23716 19660
rect 23756 19712 23808 19718
rect 23756 19654 23808 19660
rect 23388 19440 23440 19446
rect 23388 19382 23440 19388
rect 23572 19440 23624 19446
rect 23572 19382 23624 19388
rect 23400 18698 23428 19382
rect 23584 19174 23612 19382
rect 23676 19378 23704 19654
rect 23768 19378 23796 19654
rect 23860 19514 23888 19722
rect 23848 19508 23900 19514
rect 23848 19450 23900 19456
rect 24044 19378 24072 19994
rect 24412 19854 24440 20266
rect 24400 19848 24452 19854
rect 24400 19790 24452 19796
rect 25228 19848 25280 19854
rect 25228 19790 25280 19796
rect 23664 19372 23716 19378
rect 23664 19314 23716 19320
rect 23756 19372 23808 19378
rect 23756 19314 23808 19320
rect 24032 19372 24084 19378
rect 24032 19314 24084 19320
rect 23572 19168 23624 19174
rect 23572 19110 23624 19116
rect 23388 18692 23440 18698
rect 23388 18634 23440 18640
rect 23400 18358 23428 18634
rect 23572 18624 23624 18630
rect 23572 18566 23624 18572
rect 23388 18352 23440 18358
rect 23388 18294 23440 18300
rect 23584 18290 23612 18566
rect 23572 18284 23624 18290
rect 23572 18226 23624 18232
rect 23204 17604 23256 17610
rect 23204 17546 23256 17552
rect 23296 17604 23348 17610
rect 23296 17546 23348 17552
rect 23216 17338 23244 17546
rect 22836 17332 22888 17338
rect 22836 17274 22888 17280
rect 23204 17332 23256 17338
rect 23204 17274 23256 17280
rect 22376 17196 22428 17202
rect 22376 17138 22428 17144
rect 22836 16992 22888 16998
rect 22836 16934 22888 16940
rect 23388 16992 23440 16998
rect 23388 16934 23440 16940
rect 22848 16522 22876 16934
rect 23112 16584 23164 16590
rect 23112 16526 23164 16532
rect 22836 16516 22888 16522
rect 22836 16458 22888 16464
rect 22008 15700 22060 15706
rect 22008 15642 22060 15648
rect 22192 15496 22244 15502
rect 22192 15438 22244 15444
rect 22008 15020 22060 15026
rect 22008 14962 22060 14968
rect 22020 14346 22048 14962
rect 22008 14340 22060 14346
rect 22008 14282 22060 14288
rect 21732 12378 21784 12384
rect 21836 12406 21956 12434
rect 21836 10690 21864 12406
rect 21456 10668 21508 10674
rect 21456 10610 21508 10616
rect 21744 10662 21864 10690
rect 22204 10674 22232 15438
rect 22284 15156 22336 15162
rect 22284 15098 22336 15104
rect 22296 15026 22324 15098
rect 22284 15020 22336 15026
rect 22284 14962 22336 14968
rect 22282 14920 22338 14929
rect 22282 14855 22284 14864
rect 22336 14855 22338 14864
rect 22284 14826 22336 14832
rect 22296 14414 22324 14826
rect 22744 14544 22796 14550
rect 22744 14486 22796 14492
rect 22284 14408 22336 14414
rect 22284 14350 22336 14356
rect 22560 14408 22612 14414
rect 22560 14350 22612 14356
rect 22296 13802 22324 14350
rect 22572 14074 22600 14350
rect 22560 14068 22612 14074
rect 22560 14010 22612 14016
rect 22284 13796 22336 13802
rect 22284 13738 22336 13744
rect 22756 11694 22784 14486
rect 22848 14346 22876 16458
rect 23124 14550 23152 16526
rect 23400 16454 23428 16934
rect 23584 16794 23612 18226
rect 23676 18222 23704 19314
rect 23756 18964 23808 18970
rect 23756 18906 23808 18912
rect 23768 18290 23796 18906
rect 23848 18692 23900 18698
rect 23848 18634 23900 18640
rect 23860 18290 23888 18634
rect 24044 18630 24072 19314
rect 24412 19310 24440 19790
rect 25240 19378 25268 19790
rect 25228 19372 25280 19378
rect 25228 19314 25280 19320
rect 24400 19304 24452 19310
rect 24400 19246 24452 19252
rect 24952 19304 25004 19310
rect 24952 19246 25004 19252
rect 24676 18760 24728 18766
rect 24676 18702 24728 18708
rect 24032 18624 24084 18630
rect 24032 18566 24084 18572
rect 24688 18426 24716 18702
rect 24676 18420 24728 18426
rect 24676 18362 24728 18368
rect 24964 18290 24992 19246
rect 23756 18284 23808 18290
rect 23756 18226 23808 18232
rect 23848 18284 23900 18290
rect 23848 18226 23900 18232
rect 24400 18284 24452 18290
rect 24400 18226 24452 18232
rect 24952 18284 25004 18290
rect 24952 18226 25004 18232
rect 23664 18216 23716 18222
rect 23664 18158 23716 18164
rect 23676 17882 23704 18158
rect 24412 17882 24440 18226
rect 24584 18080 24636 18086
rect 24584 18022 24636 18028
rect 24596 17882 24624 18022
rect 23664 17876 23716 17882
rect 23664 17818 23716 17824
rect 24400 17876 24452 17882
rect 24400 17818 24452 17824
rect 24584 17876 24636 17882
rect 24584 17818 24636 17824
rect 24596 17678 24624 17818
rect 24584 17672 24636 17678
rect 24584 17614 24636 17620
rect 24860 17672 24912 17678
rect 24860 17614 24912 17620
rect 23664 17536 23716 17542
rect 23664 17478 23716 17484
rect 23676 17202 23704 17478
rect 24596 17202 24624 17614
rect 24872 17202 24900 17614
rect 24964 17338 24992 18226
rect 25044 18216 25096 18222
rect 25044 18158 25096 18164
rect 25056 17882 25084 18158
rect 25044 17876 25096 17882
rect 25044 17818 25096 17824
rect 24952 17332 25004 17338
rect 24952 17274 25004 17280
rect 23664 17196 23716 17202
rect 23664 17138 23716 17144
rect 24584 17196 24636 17202
rect 24584 17138 24636 17144
rect 24860 17196 24912 17202
rect 24860 17138 24912 17144
rect 23572 16788 23624 16794
rect 23572 16730 23624 16736
rect 23388 16448 23440 16454
rect 23388 16390 23440 16396
rect 23572 15496 23624 15502
rect 23572 15438 23624 15444
rect 23204 15020 23256 15026
rect 23204 14962 23256 14968
rect 23112 14544 23164 14550
rect 23112 14486 23164 14492
rect 23216 14346 23244 14962
rect 22836 14340 22888 14346
rect 22836 14282 22888 14288
rect 23204 14340 23256 14346
rect 23204 14282 23256 14288
rect 22744 11688 22796 11694
rect 22744 11630 22796 11636
rect 22376 11144 22428 11150
rect 22376 11086 22428 11092
rect 22284 11008 22336 11014
rect 22284 10950 22336 10956
rect 22008 10668 22060 10674
rect 21468 10130 21496 10610
rect 21640 10464 21692 10470
rect 21640 10406 21692 10412
rect 21456 10124 21508 10130
rect 21456 10066 21508 10072
rect 21180 9988 21232 9994
rect 21180 9930 21232 9936
rect 21364 9988 21416 9994
rect 21364 9930 21416 9936
rect 21376 9874 21404 9930
rect 21100 9846 21404 9874
rect 21376 8974 21404 9846
rect 21468 9178 21496 10066
rect 21652 10062 21680 10406
rect 21640 10056 21692 10062
rect 21640 9998 21692 10004
rect 21456 9172 21508 9178
rect 21456 9114 21508 9120
rect 21640 9172 21692 9178
rect 21640 9114 21692 9120
rect 21652 8974 21680 9114
rect 21364 8968 21416 8974
rect 21364 8910 21416 8916
rect 21640 8968 21692 8974
rect 21640 8910 21692 8916
rect 20352 8832 20404 8838
rect 20352 8774 20404 8780
rect 20444 8832 20496 8838
rect 20444 8774 20496 8780
rect 20260 8628 20312 8634
rect 20260 8570 20312 8576
rect 20352 8492 20404 8498
rect 20352 8434 20404 8440
rect 20364 8090 20392 8434
rect 20352 8084 20404 8090
rect 20352 8026 20404 8032
rect 20456 7954 20484 8774
rect 20536 8492 20588 8498
rect 20536 8434 20588 8440
rect 20444 7948 20496 7954
rect 20444 7890 20496 7896
rect 20260 6792 20312 6798
rect 20260 6734 20312 6740
rect 20272 6662 20300 6734
rect 20260 6656 20312 6662
rect 20260 6598 20312 6604
rect 20352 6656 20404 6662
rect 20352 6598 20404 6604
rect 20260 5772 20312 5778
rect 20260 5714 20312 5720
rect 20272 4622 20300 5714
rect 20364 5710 20392 6598
rect 20352 5704 20404 5710
rect 20352 5646 20404 5652
rect 20444 5568 20496 5574
rect 20444 5510 20496 5516
rect 20456 4826 20484 5510
rect 20444 4820 20496 4826
rect 20444 4762 20496 4768
rect 20260 4616 20312 4622
rect 20260 4558 20312 4564
rect 20272 4146 20300 4558
rect 20352 4276 20404 4282
rect 20352 4218 20404 4224
rect 20260 4140 20312 4146
rect 20260 4082 20312 4088
rect 20272 3534 20300 4082
rect 20364 3534 20392 4218
rect 20456 4214 20484 4762
rect 20548 4690 20576 8434
rect 20720 8356 20772 8362
rect 20720 8298 20772 8304
rect 20732 6730 20760 8298
rect 21272 8084 21324 8090
rect 21272 8026 21324 8032
rect 21284 7886 21312 8026
rect 21272 7880 21324 7886
rect 21272 7822 21324 7828
rect 21088 7812 21140 7818
rect 21088 7754 21140 7760
rect 21100 7410 21128 7754
rect 21180 7540 21232 7546
rect 21180 7482 21232 7488
rect 21088 7404 21140 7410
rect 21088 7346 21140 7352
rect 20720 6724 20772 6730
rect 20720 6666 20772 6672
rect 20904 6724 20956 6730
rect 20904 6666 20956 6672
rect 20996 6724 21048 6730
rect 20996 6666 21048 6672
rect 20732 6322 20760 6666
rect 20916 6390 20944 6666
rect 21008 6458 21036 6666
rect 20996 6452 21048 6458
rect 20996 6394 21048 6400
rect 20904 6384 20956 6390
rect 20904 6326 20956 6332
rect 20720 6316 20772 6322
rect 20720 6258 20772 6264
rect 20732 5778 20760 6258
rect 20720 5772 20772 5778
rect 20720 5714 20772 5720
rect 20916 5574 20944 6326
rect 21100 6118 21128 7346
rect 21192 7002 21220 7482
rect 21180 6996 21232 7002
rect 21180 6938 21232 6944
rect 21088 6112 21140 6118
rect 21088 6054 21140 6060
rect 21284 5846 21312 7822
rect 21376 6866 21404 8910
rect 21652 8634 21680 8910
rect 21640 8628 21692 8634
rect 21560 8588 21640 8616
rect 21560 7002 21588 8588
rect 21640 8570 21692 8576
rect 21640 7336 21692 7342
rect 21640 7278 21692 7284
rect 21548 6996 21600 7002
rect 21548 6938 21600 6944
rect 21364 6860 21416 6866
rect 21364 6802 21416 6808
rect 21376 6186 21404 6802
rect 21560 6322 21588 6938
rect 21652 6934 21680 7278
rect 21640 6928 21692 6934
rect 21640 6870 21692 6876
rect 21548 6316 21600 6322
rect 21548 6258 21600 6264
rect 21364 6180 21416 6186
rect 21364 6122 21416 6128
rect 21272 5840 21324 5846
rect 21272 5782 21324 5788
rect 21652 5710 21680 6870
rect 21640 5704 21692 5710
rect 21192 5652 21640 5658
rect 21192 5646 21692 5652
rect 21192 5642 21680 5646
rect 21180 5636 21680 5642
rect 21232 5630 21680 5636
rect 21180 5578 21232 5584
rect 20904 5568 20956 5574
rect 20904 5510 20956 5516
rect 20536 4684 20588 4690
rect 20536 4626 20588 4632
rect 20548 4282 20576 4626
rect 21744 4622 21772 10662
rect 22008 10610 22060 10616
rect 22192 10668 22244 10674
rect 22192 10610 22244 10616
rect 21824 10600 21876 10606
rect 21824 10542 21876 10548
rect 21836 10266 21864 10542
rect 21824 10260 21876 10266
rect 21824 10202 21876 10208
rect 22020 10198 22048 10610
rect 22008 10192 22060 10198
rect 22008 10134 22060 10140
rect 22100 9920 22152 9926
rect 22100 9862 22152 9868
rect 22112 9110 22140 9862
rect 22100 9104 22152 9110
rect 22100 9046 22152 9052
rect 21916 8968 21968 8974
rect 21916 8910 21968 8916
rect 22008 8968 22060 8974
rect 22008 8910 22060 8916
rect 21928 8362 21956 8910
rect 22020 8498 22048 8910
rect 22008 8492 22060 8498
rect 22008 8434 22060 8440
rect 21916 8356 21968 8362
rect 21916 8298 21968 8304
rect 22112 7274 22140 9046
rect 22204 8974 22232 10610
rect 22296 10470 22324 10950
rect 22284 10464 22336 10470
rect 22284 10406 22336 10412
rect 22296 10062 22324 10406
rect 22388 10062 22416 11086
rect 22560 10668 22612 10674
rect 22560 10610 22612 10616
rect 22572 10266 22600 10610
rect 22848 10606 22876 14282
rect 22928 14000 22980 14006
rect 22928 13942 22980 13948
rect 23018 13968 23074 13977
rect 22940 13530 22968 13942
rect 23018 13903 23020 13912
rect 23072 13903 23074 13912
rect 23020 13874 23072 13880
rect 22928 13524 22980 13530
rect 22928 13466 22980 13472
rect 22928 13184 22980 13190
rect 23032 13172 23060 13874
rect 22980 13144 23060 13172
rect 22928 13126 22980 13132
rect 23216 12434 23244 14282
rect 23386 13968 23442 13977
rect 23386 13903 23388 13912
rect 23440 13903 23442 13912
rect 23388 13874 23440 13880
rect 23296 13864 23348 13870
rect 23296 13806 23348 13812
rect 23308 13258 23336 13806
rect 23296 13252 23348 13258
rect 23296 13194 23348 13200
rect 23124 12406 23244 12434
rect 23020 12232 23072 12238
rect 23020 12174 23072 12180
rect 22928 12096 22980 12102
rect 22928 12038 22980 12044
rect 22836 10600 22888 10606
rect 22836 10542 22888 10548
rect 22560 10260 22612 10266
rect 22560 10202 22612 10208
rect 22284 10056 22336 10062
rect 22284 9998 22336 10004
rect 22376 10056 22428 10062
rect 22376 9998 22428 10004
rect 22940 9994 22968 12038
rect 23032 11830 23060 12174
rect 23020 11824 23072 11830
rect 23020 11766 23072 11772
rect 23124 11354 23152 12406
rect 23204 12232 23256 12238
rect 23204 12174 23256 12180
rect 23216 11898 23244 12174
rect 23204 11892 23256 11898
rect 23204 11834 23256 11840
rect 23308 11540 23336 13194
rect 23388 13184 23440 13190
rect 23388 13126 23440 13132
rect 23400 12238 23428 13126
rect 23584 12434 23612 15438
rect 23492 12406 23612 12434
rect 23388 12232 23440 12238
rect 23388 12174 23440 12180
rect 23492 11762 23520 12406
rect 23676 12050 23704 17138
rect 24032 16584 24084 16590
rect 24032 16526 24084 16532
rect 24044 15366 24072 16526
rect 24596 16114 24624 17138
rect 24872 16114 24900 17138
rect 25136 16448 25188 16454
rect 25136 16390 25188 16396
rect 24952 16176 25004 16182
rect 24952 16118 25004 16124
rect 24584 16108 24636 16114
rect 24584 16050 24636 16056
rect 24860 16108 24912 16114
rect 24860 16050 24912 16056
rect 24676 15564 24728 15570
rect 24676 15506 24728 15512
rect 24124 15496 24176 15502
rect 24124 15438 24176 15444
rect 24216 15496 24268 15502
rect 24216 15438 24268 15444
rect 24032 15360 24084 15366
rect 24032 15302 24084 15308
rect 24136 15162 24164 15438
rect 24124 15156 24176 15162
rect 24124 15098 24176 15104
rect 23940 15020 23992 15026
rect 23940 14962 23992 14968
rect 23952 14482 23980 14962
rect 24124 14612 24176 14618
rect 24124 14554 24176 14560
rect 23940 14476 23992 14482
rect 23940 14418 23992 14424
rect 24136 14278 24164 14554
rect 24124 14272 24176 14278
rect 24124 14214 24176 14220
rect 24136 13530 24164 14214
rect 24124 13524 24176 13530
rect 24124 13466 24176 13472
rect 23848 13252 23900 13258
rect 23848 13194 23900 13200
rect 23860 12918 23888 13194
rect 23848 12912 23900 12918
rect 23848 12854 23900 12860
rect 24032 12164 24084 12170
rect 24032 12106 24084 12112
rect 23584 12022 23704 12050
rect 23940 12096 23992 12102
rect 23940 12038 23992 12044
rect 23480 11756 23532 11762
rect 23480 11698 23532 11704
rect 23388 11552 23440 11558
rect 23308 11512 23388 11540
rect 23388 11494 23440 11500
rect 23112 11348 23164 11354
rect 23112 11290 23164 11296
rect 22928 9988 22980 9994
rect 22928 9930 22980 9936
rect 22284 9036 22336 9042
rect 22284 8978 22336 8984
rect 22192 8968 22244 8974
rect 22192 8910 22244 8916
rect 22192 8832 22244 8838
rect 22192 8774 22244 8780
rect 22204 8498 22232 8774
rect 22192 8492 22244 8498
rect 22192 8434 22244 8440
rect 22296 7886 22324 8978
rect 22376 8968 22428 8974
rect 22376 8910 22428 8916
rect 22388 8634 22416 8910
rect 22652 8832 22704 8838
rect 22652 8774 22704 8780
rect 22744 8832 22796 8838
rect 22744 8774 22796 8780
rect 22376 8628 22428 8634
rect 22376 8570 22428 8576
rect 22388 7886 22416 8570
rect 22284 7880 22336 7886
rect 22284 7822 22336 7828
rect 22376 7880 22428 7886
rect 22376 7822 22428 7828
rect 22376 7540 22428 7546
rect 22376 7482 22428 7488
rect 22100 7268 22152 7274
rect 22100 7210 22152 7216
rect 22284 7268 22336 7274
rect 22284 7210 22336 7216
rect 21916 6316 21968 6322
rect 21916 6258 21968 6264
rect 21824 6180 21876 6186
rect 21824 6122 21876 6128
rect 21836 5030 21864 6122
rect 21928 5302 21956 6258
rect 22192 5840 22244 5846
rect 22192 5782 22244 5788
rect 22204 5710 22232 5782
rect 22296 5778 22324 7210
rect 22388 6934 22416 7482
rect 22664 7478 22692 8774
rect 22756 8498 22784 8774
rect 22744 8492 22796 8498
rect 22744 8434 22796 8440
rect 22940 7750 22968 9930
rect 23296 8968 23348 8974
rect 23296 8910 23348 8916
rect 23308 8498 23336 8910
rect 23296 8492 23348 8498
rect 23296 8434 23348 8440
rect 23400 8362 23428 11494
rect 23492 11218 23520 11698
rect 23584 11694 23612 12022
rect 23952 11830 23980 12038
rect 23940 11824 23992 11830
rect 23940 11766 23992 11772
rect 23572 11688 23624 11694
rect 23570 11656 23572 11665
rect 23848 11688 23900 11694
rect 23624 11656 23626 11665
rect 23848 11630 23900 11636
rect 23570 11591 23626 11600
rect 23480 11212 23532 11218
rect 23480 11154 23532 11160
rect 23756 11212 23808 11218
rect 23756 11154 23808 11160
rect 23572 10124 23624 10130
rect 23572 10066 23624 10072
rect 23480 10056 23532 10062
rect 23480 9998 23532 10004
rect 23388 8356 23440 8362
rect 23388 8298 23440 8304
rect 23492 7886 23520 9998
rect 23584 9722 23612 10066
rect 23572 9716 23624 9722
rect 23572 9658 23624 9664
rect 23768 9586 23796 11154
rect 23860 9586 23888 11630
rect 23940 10056 23992 10062
rect 24044 10044 24072 12106
rect 24228 10674 24256 15438
rect 24584 15360 24636 15366
rect 24584 15302 24636 15308
rect 24492 15156 24544 15162
rect 24492 15098 24544 15104
rect 24308 14816 24360 14822
rect 24308 14758 24360 14764
rect 24320 11354 24348 14758
rect 24504 14618 24532 15098
rect 24596 14822 24624 15302
rect 24688 15026 24716 15506
rect 24872 15162 24900 16050
rect 24964 15434 24992 16118
rect 25044 15564 25096 15570
rect 25044 15506 25096 15512
rect 24952 15428 25004 15434
rect 24952 15370 25004 15376
rect 24860 15156 24912 15162
rect 24860 15098 24912 15104
rect 24676 15020 24728 15026
rect 24676 14962 24728 14968
rect 24584 14816 24636 14822
rect 24584 14758 24636 14764
rect 24492 14612 24544 14618
rect 24492 14554 24544 14560
rect 24400 12640 24452 12646
rect 24400 12582 24452 12588
rect 24412 11762 24440 12582
rect 24492 12300 24544 12306
rect 24492 12242 24544 12248
rect 24504 11898 24532 12242
rect 24492 11892 24544 11898
rect 24492 11834 24544 11840
rect 24400 11756 24452 11762
rect 24400 11698 24452 11704
rect 24308 11348 24360 11354
rect 24308 11290 24360 11296
rect 24320 10674 24348 11290
rect 24216 10668 24268 10674
rect 24216 10610 24268 10616
rect 24308 10668 24360 10674
rect 24308 10610 24360 10616
rect 24412 10198 24440 11698
rect 24596 11150 24624 14758
rect 25056 13938 25084 15506
rect 25148 15366 25176 16390
rect 25240 16182 25268 19314
rect 25332 17338 25360 20878
rect 25596 18284 25648 18290
rect 25596 18226 25648 18232
rect 25608 18086 25636 18226
rect 25596 18080 25648 18086
rect 25596 18022 25648 18028
rect 25320 17332 25372 17338
rect 25320 17274 25372 17280
rect 25504 17196 25556 17202
rect 25504 17138 25556 17144
rect 25228 16176 25280 16182
rect 25228 16118 25280 16124
rect 25516 16114 25544 17138
rect 25608 16998 25636 18022
rect 25780 17536 25832 17542
rect 25780 17478 25832 17484
rect 25792 17202 25820 17478
rect 26424 17332 26476 17338
rect 26424 17274 26476 17280
rect 25780 17196 25832 17202
rect 25780 17138 25832 17144
rect 25872 17196 25924 17202
rect 25872 17138 25924 17144
rect 25596 16992 25648 16998
rect 25596 16934 25648 16940
rect 25504 16108 25556 16114
rect 25504 16050 25556 16056
rect 25320 15904 25372 15910
rect 25320 15846 25372 15852
rect 25228 15496 25280 15502
rect 25228 15438 25280 15444
rect 25136 15360 25188 15366
rect 25240 15337 25268 15438
rect 25332 15434 25360 15846
rect 25516 15706 25544 16050
rect 25504 15700 25556 15706
rect 25504 15642 25556 15648
rect 25320 15428 25372 15434
rect 25320 15370 25372 15376
rect 25136 15302 25188 15308
rect 25226 15328 25282 15337
rect 25148 15162 25176 15302
rect 25226 15263 25282 15272
rect 25332 15178 25360 15370
rect 25136 15156 25188 15162
rect 25136 15098 25188 15104
rect 25240 15150 25360 15178
rect 25240 13938 25268 15150
rect 25044 13932 25096 13938
rect 25044 13874 25096 13880
rect 25228 13932 25280 13938
rect 25228 13874 25280 13880
rect 24768 13252 24820 13258
rect 24768 13194 24820 13200
rect 24952 13252 25004 13258
rect 24952 13194 25004 13200
rect 24676 12912 24728 12918
rect 24676 12854 24728 12860
rect 24688 12646 24716 12854
rect 24780 12646 24808 13194
rect 24860 12980 24912 12986
rect 24860 12922 24912 12928
rect 24872 12782 24900 12922
rect 24860 12776 24912 12782
rect 24860 12718 24912 12724
rect 24676 12640 24728 12646
rect 24676 12582 24728 12588
rect 24768 12640 24820 12646
rect 24768 12582 24820 12588
rect 24872 11898 24900 12718
rect 24964 12646 24992 13194
rect 24952 12640 25004 12646
rect 24952 12582 25004 12588
rect 24860 11892 24912 11898
rect 24860 11834 24912 11840
rect 24964 11762 24992 12582
rect 25240 12170 25268 13874
rect 25412 13864 25464 13870
rect 25412 13806 25464 13812
rect 25596 13864 25648 13870
rect 25596 13806 25648 13812
rect 25320 13456 25372 13462
rect 25320 13398 25372 13404
rect 25228 12164 25280 12170
rect 25228 12106 25280 12112
rect 24952 11756 25004 11762
rect 24952 11698 25004 11704
rect 24584 11144 24636 11150
rect 24584 11086 24636 11092
rect 24492 10668 24544 10674
rect 24492 10610 24544 10616
rect 24400 10192 24452 10198
rect 24400 10134 24452 10140
rect 23992 10016 24072 10044
rect 23940 9998 23992 10004
rect 23756 9580 23808 9586
rect 23756 9522 23808 9528
rect 23848 9580 23900 9586
rect 23848 9522 23900 9528
rect 23860 9042 23888 9522
rect 23848 9036 23900 9042
rect 23848 8978 23900 8984
rect 23952 8922 23980 9998
rect 24032 9920 24084 9926
rect 24032 9862 24084 9868
rect 24044 9586 24072 9862
rect 24032 9580 24084 9586
rect 24032 9522 24084 9528
rect 23860 8894 23980 8922
rect 24216 8968 24268 8974
rect 24216 8910 24268 8916
rect 24400 8968 24452 8974
rect 24400 8910 24452 8916
rect 23480 7880 23532 7886
rect 23480 7822 23532 7828
rect 22928 7744 22980 7750
rect 22928 7686 22980 7692
rect 22940 7478 22968 7686
rect 23492 7546 23520 7822
rect 23860 7750 23888 8894
rect 24124 8832 24176 8838
rect 24124 8774 24176 8780
rect 23848 7744 23900 7750
rect 23848 7686 23900 7692
rect 23480 7540 23532 7546
rect 23480 7482 23532 7488
rect 22652 7472 22704 7478
rect 22652 7414 22704 7420
rect 22928 7472 22980 7478
rect 22928 7414 22980 7420
rect 23860 7410 23888 7686
rect 24136 7410 24164 8774
rect 24228 8566 24256 8910
rect 24216 8560 24268 8566
rect 24216 8502 24268 8508
rect 24228 7954 24256 8502
rect 24412 8498 24440 8910
rect 24504 8838 24532 10610
rect 24596 9654 24624 11086
rect 24676 10668 24728 10674
rect 24676 10610 24728 10616
rect 24584 9648 24636 9654
rect 24584 9590 24636 9596
rect 24596 9110 24624 9590
rect 24584 9104 24636 9110
rect 24584 9046 24636 9052
rect 24688 8974 24716 10610
rect 24676 8968 24728 8974
rect 24676 8910 24728 8916
rect 24492 8832 24544 8838
rect 24492 8774 24544 8780
rect 24400 8492 24452 8498
rect 24400 8434 24452 8440
rect 24412 8090 24440 8434
rect 24400 8084 24452 8090
rect 24400 8026 24452 8032
rect 24216 7948 24268 7954
rect 24216 7890 24268 7896
rect 24308 7812 24360 7818
rect 24308 7754 24360 7760
rect 24320 7410 24348 7754
rect 23848 7404 23900 7410
rect 23848 7346 23900 7352
rect 24124 7404 24176 7410
rect 24124 7346 24176 7352
rect 24308 7404 24360 7410
rect 24308 7346 24360 7352
rect 23756 7336 23808 7342
rect 23756 7278 23808 7284
rect 23388 7200 23440 7206
rect 23388 7142 23440 7148
rect 22376 6928 22428 6934
rect 22376 6870 22428 6876
rect 23400 6798 23428 7142
rect 23768 7002 23796 7278
rect 23756 6996 23808 7002
rect 23756 6938 23808 6944
rect 23388 6792 23440 6798
rect 23388 6734 23440 6740
rect 23572 6792 23624 6798
rect 23572 6734 23624 6740
rect 23756 6792 23808 6798
rect 23756 6734 23808 6740
rect 23584 6458 23612 6734
rect 23664 6656 23716 6662
rect 23664 6598 23716 6604
rect 23572 6452 23624 6458
rect 23572 6394 23624 6400
rect 23204 6316 23256 6322
rect 23204 6258 23256 6264
rect 23480 6316 23532 6322
rect 23480 6258 23532 6264
rect 23216 5914 23244 6258
rect 23492 6186 23520 6258
rect 23480 6180 23532 6186
rect 23480 6122 23532 6128
rect 23204 5908 23256 5914
rect 23204 5850 23256 5856
rect 22376 5840 22428 5846
rect 22376 5782 22428 5788
rect 22284 5772 22336 5778
rect 22284 5714 22336 5720
rect 22192 5704 22244 5710
rect 22192 5646 22244 5652
rect 22100 5364 22152 5370
rect 22100 5306 22152 5312
rect 21916 5296 21968 5302
rect 21916 5238 21968 5244
rect 21824 5024 21876 5030
rect 21824 4966 21876 4972
rect 21732 4616 21784 4622
rect 21732 4558 21784 4564
rect 20628 4480 20680 4486
rect 20628 4422 20680 4428
rect 21640 4480 21692 4486
rect 21640 4422 21692 4428
rect 20536 4276 20588 4282
rect 20536 4218 20588 4224
rect 20444 4208 20496 4214
rect 20444 4150 20496 4156
rect 20456 3738 20484 4150
rect 20536 4140 20588 4146
rect 20536 4082 20588 4088
rect 20444 3732 20496 3738
rect 20444 3674 20496 3680
rect 20260 3528 20312 3534
rect 20260 3470 20312 3476
rect 20352 3528 20404 3534
rect 20352 3470 20404 3476
rect 20548 3398 20576 4082
rect 20640 4010 20668 4422
rect 20628 4004 20680 4010
rect 20628 3946 20680 3952
rect 21456 4004 21508 4010
rect 21456 3946 21508 3952
rect 20640 3602 20668 3946
rect 21272 3664 21324 3670
rect 21272 3606 21324 3612
rect 20628 3596 20680 3602
rect 20628 3538 20680 3544
rect 21284 3534 21312 3606
rect 21272 3528 21324 3534
rect 21272 3470 21324 3476
rect 21468 3466 21496 3946
rect 21652 3534 21680 4422
rect 21640 3528 21692 3534
rect 21640 3470 21692 3476
rect 21456 3460 21508 3466
rect 21456 3402 21508 3408
rect 20536 3392 20588 3398
rect 20536 3334 20588 3340
rect 21744 3194 21772 4558
rect 21836 4486 21864 4966
rect 21928 4758 21956 5238
rect 22112 5098 22140 5306
rect 22100 5092 22152 5098
rect 22100 5034 22152 5040
rect 21916 4752 21968 4758
rect 21916 4694 21968 4700
rect 21824 4480 21876 4486
rect 21824 4422 21876 4428
rect 21824 4072 21876 4078
rect 21824 4014 21876 4020
rect 21836 3602 21864 4014
rect 21928 3738 21956 4694
rect 22296 4146 22324 5714
rect 22388 5234 22416 5782
rect 22928 5704 22980 5710
rect 22928 5646 22980 5652
rect 23492 5658 23520 6122
rect 23584 5846 23612 6394
rect 23572 5840 23624 5846
rect 23572 5782 23624 5788
rect 22560 5636 22612 5642
rect 22560 5578 22612 5584
rect 22572 5234 22600 5578
rect 22940 5370 22968 5646
rect 23492 5630 23612 5658
rect 23204 5568 23256 5574
rect 23204 5510 23256 5516
rect 23480 5568 23532 5574
rect 23480 5510 23532 5516
rect 22928 5364 22980 5370
rect 22928 5306 22980 5312
rect 22376 5228 22428 5234
rect 22376 5170 22428 5176
rect 22560 5228 22612 5234
rect 22560 5170 22612 5176
rect 22940 5166 22968 5306
rect 23216 5166 23244 5510
rect 22928 5160 22980 5166
rect 22928 5102 22980 5108
rect 23204 5160 23256 5166
rect 23204 5102 23256 5108
rect 22376 5024 22428 5030
rect 22376 4966 22428 4972
rect 22388 4826 22416 4966
rect 22376 4820 22428 4826
rect 22376 4762 22428 4768
rect 23492 4146 23520 5510
rect 23584 4826 23612 5630
rect 23572 4820 23624 4826
rect 23572 4762 23624 4768
rect 22284 4140 22336 4146
rect 22284 4082 22336 4088
rect 22376 4140 22428 4146
rect 22376 4082 22428 4088
rect 23204 4140 23256 4146
rect 23204 4082 23256 4088
rect 23480 4140 23532 4146
rect 23480 4082 23532 4088
rect 21916 3732 21968 3738
rect 21916 3674 21968 3680
rect 22388 3670 22416 4082
rect 23216 3738 23244 4082
rect 23676 4078 23704 6598
rect 23768 5710 23796 6734
rect 24320 5846 24348 7346
rect 24504 7342 24532 8774
rect 24688 8566 24716 8910
rect 24676 8560 24728 8566
rect 24676 8502 24728 8508
rect 24964 7546 24992 11698
rect 25136 8832 25188 8838
rect 25136 8774 25188 8780
rect 25148 8430 25176 8774
rect 25136 8424 25188 8430
rect 25136 8366 25188 8372
rect 24952 7540 25004 7546
rect 24952 7482 25004 7488
rect 25228 7472 25280 7478
rect 25228 7414 25280 7420
rect 25136 7404 25188 7410
rect 25136 7346 25188 7352
rect 24492 7336 24544 7342
rect 24492 7278 24544 7284
rect 25044 6996 25096 7002
rect 25044 6938 25096 6944
rect 24952 6860 25004 6866
rect 24952 6802 25004 6808
rect 24308 5840 24360 5846
rect 24308 5782 24360 5788
rect 24964 5710 24992 6802
rect 25056 6798 25084 6938
rect 25044 6792 25096 6798
rect 25044 6734 25096 6740
rect 23756 5704 23808 5710
rect 23756 5646 23808 5652
rect 24032 5704 24084 5710
rect 24032 5646 24084 5652
rect 24952 5704 25004 5710
rect 24952 5646 25004 5652
rect 23768 5234 23796 5646
rect 24044 5370 24072 5646
rect 24860 5568 24912 5574
rect 24398 5536 24454 5545
rect 24860 5510 24912 5516
rect 24398 5471 24454 5480
rect 24032 5364 24084 5370
rect 24032 5306 24084 5312
rect 23756 5228 23808 5234
rect 23756 5170 23808 5176
rect 24308 4820 24360 4826
rect 24308 4762 24360 4768
rect 24320 4146 24348 4762
rect 24412 4622 24440 5471
rect 24872 5234 24900 5510
rect 24860 5228 24912 5234
rect 24860 5170 24912 5176
rect 24400 4616 24452 4622
rect 24400 4558 24452 4564
rect 24676 4616 24728 4622
rect 24676 4558 24728 4564
rect 24308 4140 24360 4146
rect 24308 4082 24360 4088
rect 23664 4072 23716 4078
rect 23664 4014 23716 4020
rect 23480 4004 23532 4010
rect 23480 3946 23532 3952
rect 23204 3732 23256 3738
rect 23204 3674 23256 3680
rect 22376 3664 22428 3670
rect 22376 3606 22428 3612
rect 21824 3596 21876 3602
rect 21824 3538 21876 3544
rect 22388 3534 22416 3606
rect 22376 3528 22428 3534
rect 22376 3470 22428 3476
rect 23492 3466 23520 3946
rect 24412 3942 24440 4558
rect 24688 4146 24716 4558
rect 24964 4146 24992 5646
rect 25056 5574 25084 6734
rect 25148 6662 25176 7346
rect 25240 7206 25268 7414
rect 25228 7200 25280 7206
rect 25228 7142 25280 7148
rect 25240 6798 25268 7142
rect 25228 6792 25280 6798
rect 25228 6734 25280 6740
rect 25136 6656 25188 6662
rect 25136 6598 25188 6604
rect 25148 6254 25176 6598
rect 25136 6248 25188 6254
rect 25136 6190 25188 6196
rect 25240 5778 25268 6734
rect 25228 5772 25280 5778
rect 25228 5714 25280 5720
rect 25044 5568 25096 5574
rect 25044 5510 25096 5516
rect 25056 4826 25084 5510
rect 25332 5370 25360 13398
rect 25424 12102 25452 13806
rect 25608 13530 25636 13806
rect 25780 13796 25832 13802
rect 25780 13738 25832 13744
rect 25596 13524 25648 13530
rect 25596 13466 25648 13472
rect 25792 13394 25820 13738
rect 25780 13388 25832 13394
rect 25780 13330 25832 13336
rect 25688 12844 25740 12850
rect 25688 12786 25740 12792
rect 25700 12306 25728 12786
rect 25792 12714 25820 13330
rect 25780 12708 25832 12714
rect 25780 12650 25832 12656
rect 25792 12442 25820 12650
rect 25780 12436 25832 12442
rect 25884 12434 25912 17138
rect 26436 15502 26464 17274
rect 26424 15496 26476 15502
rect 26424 15438 26476 15444
rect 26436 13938 26464 15438
rect 26608 14408 26660 14414
rect 26608 14350 26660 14356
rect 26700 14408 26752 14414
rect 26700 14350 26752 14356
rect 26620 14074 26648 14350
rect 26608 14068 26660 14074
rect 26608 14010 26660 14016
rect 26424 13932 26476 13938
rect 26424 13874 26476 13880
rect 26240 13864 26292 13870
rect 26240 13806 26292 13812
rect 26332 13864 26384 13870
rect 26332 13806 26384 13812
rect 26148 13456 26200 13462
rect 26148 13398 26200 13404
rect 26160 13326 26188 13398
rect 26148 13320 26200 13326
rect 26148 13262 26200 13268
rect 26160 13002 26188 13262
rect 26068 12974 26188 13002
rect 26068 12782 26096 12974
rect 26252 12918 26280 13806
rect 26344 13394 26372 13806
rect 26424 13728 26476 13734
rect 26424 13670 26476 13676
rect 26332 13388 26384 13394
rect 26332 13330 26384 13336
rect 26344 12986 26372 13330
rect 26332 12980 26384 12986
rect 26332 12922 26384 12928
rect 26240 12912 26292 12918
rect 26240 12854 26292 12860
rect 26148 12844 26200 12850
rect 26148 12786 26200 12792
rect 26056 12776 26108 12782
rect 26056 12718 26108 12724
rect 25884 12406 26004 12434
rect 25780 12378 25832 12384
rect 25688 12300 25740 12306
rect 25688 12242 25740 12248
rect 25976 12238 26004 12406
rect 25504 12232 25556 12238
rect 25504 12174 25556 12180
rect 25964 12232 26016 12238
rect 25964 12174 26016 12180
rect 25412 12096 25464 12102
rect 25412 12038 25464 12044
rect 25412 11824 25464 11830
rect 25412 11766 25464 11772
rect 25424 11150 25452 11766
rect 25516 11762 25544 12174
rect 25688 12096 25740 12102
rect 25688 12038 25740 12044
rect 25504 11756 25556 11762
rect 25504 11698 25556 11704
rect 25700 11626 25728 12038
rect 25688 11620 25740 11626
rect 25688 11562 25740 11568
rect 25412 11144 25464 11150
rect 25412 11086 25464 11092
rect 25700 10742 25728 11562
rect 25688 10736 25740 10742
rect 25688 10678 25740 10684
rect 25976 10266 26004 12174
rect 26056 11688 26108 11694
rect 26056 11630 26108 11636
rect 26068 11354 26096 11630
rect 26056 11348 26108 11354
rect 26056 11290 26108 11296
rect 25964 10260 26016 10266
rect 25964 10202 26016 10208
rect 25688 10192 25740 10198
rect 25688 10134 25740 10140
rect 25700 10062 25728 10134
rect 25504 10056 25556 10062
rect 25504 9998 25556 10004
rect 25688 10056 25740 10062
rect 25688 9998 25740 10004
rect 25320 5364 25372 5370
rect 25320 5306 25372 5312
rect 25136 5228 25188 5234
rect 25136 5170 25188 5176
rect 25044 4820 25096 4826
rect 25044 4762 25096 4768
rect 25148 4690 25176 5170
rect 25516 4758 25544 9998
rect 25596 9104 25648 9110
rect 25596 9046 25648 9052
rect 25608 7410 25636 9046
rect 25596 7404 25648 7410
rect 25596 7346 25648 7352
rect 25608 7002 25636 7346
rect 25596 6996 25648 7002
rect 25596 6938 25648 6944
rect 25596 6792 25648 6798
rect 25596 6734 25648 6740
rect 25608 6186 25636 6734
rect 25596 6180 25648 6186
rect 25596 6122 25648 6128
rect 25504 4752 25556 4758
rect 25504 4694 25556 4700
rect 25136 4684 25188 4690
rect 25136 4626 25188 4632
rect 25148 4282 25176 4626
rect 25136 4276 25188 4282
rect 25136 4218 25188 4224
rect 24676 4140 24728 4146
rect 24676 4082 24728 4088
rect 24952 4140 25004 4146
rect 24952 4082 25004 4088
rect 25504 4140 25556 4146
rect 25504 4082 25556 4088
rect 24400 3936 24452 3942
rect 24400 3878 24452 3884
rect 23664 3528 23716 3534
rect 23664 3470 23716 3476
rect 22468 3460 22520 3466
rect 22468 3402 22520 3408
rect 23480 3460 23532 3466
rect 23480 3402 23532 3408
rect 21916 3392 21968 3398
rect 21916 3334 21968 3340
rect 20076 3188 20128 3194
rect 20076 3130 20128 3136
rect 20168 3188 20220 3194
rect 20168 3130 20220 3136
rect 21732 3188 21784 3194
rect 21732 3130 21784 3136
rect 17776 3052 17828 3058
rect 17776 2994 17828 3000
rect 18236 3052 18288 3058
rect 18236 2994 18288 3000
rect 18420 3052 18472 3058
rect 18420 2994 18472 3000
rect 18696 3052 18748 3058
rect 18696 2994 18748 3000
rect 18880 3052 18932 3058
rect 18880 2994 18932 3000
rect 17500 2984 17552 2990
rect 17500 2926 17552 2932
rect 17132 2916 17184 2922
rect 17132 2858 17184 2864
rect 17788 2446 17816 2994
rect 18708 2922 18736 2994
rect 21928 2990 21956 3334
rect 22480 3194 22508 3402
rect 23676 3194 23704 3470
rect 24688 3466 24716 4082
rect 25516 4049 25544 4082
rect 25502 4040 25558 4049
rect 25502 3975 25558 3984
rect 24860 3936 24912 3942
rect 24860 3878 24912 3884
rect 24872 3670 24900 3878
rect 25516 3738 25544 3975
rect 25504 3732 25556 3738
rect 25504 3674 25556 3680
rect 25700 3670 25728 9998
rect 25780 9512 25832 9518
rect 25780 9454 25832 9460
rect 25792 8974 25820 9454
rect 25780 8968 25832 8974
rect 25780 8910 25832 8916
rect 25792 7546 25820 8910
rect 25780 7540 25832 7546
rect 25780 7482 25832 7488
rect 25792 6934 25820 7482
rect 25872 7268 25924 7274
rect 25872 7210 25924 7216
rect 25780 6928 25832 6934
rect 25780 6870 25832 6876
rect 25884 6798 25912 7210
rect 25872 6792 25924 6798
rect 25872 6734 25924 6740
rect 25780 6724 25832 6730
rect 25780 6666 25832 6672
rect 25792 6458 25820 6666
rect 26160 6662 26188 12786
rect 26436 12434 26464 13670
rect 26712 13258 26740 14350
rect 26700 13252 26752 13258
rect 26700 13194 26752 13200
rect 26608 12912 26660 12918
rect 26608 12854 26660 12860
rect 26344 12406 26464 12434
rect 26344 10266 26372 12406
rect 26516 11552 26568 11558
rect 26516 11494 26568 11500
rect 26332 10260 26384 10266
rect 26332 10202 26384 10208
rect 26424 10260 26476 10266
rect 26424 10202 26476 10208
rect 26436 10130 26464 10202
rect 26424 10124 26476 10130
rect 26424 10066 26476 10072
rect 26528 10062 26556 11494
rect 26620 11218 26648 12854
rect 26712 12850 26740 13194
rect 26700 12844 26752 12850
rect 26700 12786 26752 12792
rect 27160 12368 27212 12374
rect 27160 12310 27212 12316
rect 27172 11762 27200 12310
rect 27160 11756 27212 11762
rect 27160 11698 27212 11704
rect 27252 11756 27304 11762
rect 27252 11698 27304 11704
rect 27172 11286 27200 11698
rect 27160 11280 27212 11286
rect 27160 11222 27212 11228
rect 27264 11218 27292 11698
rect 26608 11212 26660 11218
rect 26608 11154 26660 11160
rect 27252 11212 27304 11218
rect 27252 11154 27304 11160
rect 26516 10056 26568 10062
rect 26516 9998 26568 10004
rect 26148 6656 26200 6662
rect 26148 6598 26200 6604
rect 25780 6452 25832 6458
rect 25780 6394 25832 6400
rect 24860 3664 24912 3670
rect 24860 3606 24912 3612
rect 25688 3664 25740 3670
rect 25688 3606 25740 3612
rect 24676 3460 24728 3466
rect 24676 3402 24728 3408
rect 22468 3188 22520 3194
rect 22468 3130 22520 3136
rect 23664 3188 23716 3194
rect 23664 3130 23716 3136
rect 21916 2984 21968 2990
rect 21916 2926 21968 2932
rect 27528 2984 27580 2990
rect 27528 2926 27580 2932
rect 18696 2916 18748 2922
rect 18696 2858 18748 2864
rect 18708 2650 18736 2858
rect 27540 2825 27568 2926
rect 27526 2816 27582 2825
rect 27526 2751 27582 2760
rect 18696 2644 18748 2650
rect 18696 2586 18748 2592
rect 15384 2382 15436 2388
rect 15580 2378 15700 2394
rect 15844 2440 15896 2446
rect 15844 2382 15896 2388
rect 16948 2440 17000 2446
rect 16948 2382 17000 2388
rect 17776 2440 17828 2446
rect 17776 2382 17828 2388
rect 15568 2372 15700 2378
rect 15620 2366 15700 2372
rect 15568 2314 15620 2320
rect 11888 2304 11940 2310
rect 11888 2246 11940 2252
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
<< via2 >>
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 1306 27920 1362 27976
rect 1214 26580 1270 26616
rect 1214 26560 1216 26580
rect 1216 26560 1268 26580
rect 1268 26560 1270 26580
rect 846 25372 848 25392
rect 848 25372 900 25392
rect 900 25372 902 25392
rect 846 25336 902 25372
rect 846 24676 902 24712
rect 846 24656 848 24676
rect 848 24656 900 24676
rect 900 24656 902 24676
rect 1214 23860 1270 23896
rect 1214 23840 1216 23860
rect 1216 23840 1268 23860
rect 1268 23840 1270 23860
rect 846 21256 902 21312
rect 1490 25880 1546 25936
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4880 28314 4936 28316
rect 4960 28314 5016 28316
rect 5040 28314 5096 28316
rect 5120 28314 5176 28316
rect 4880 28262 4926 28314
rect 4926 28262 4936 28314
rect 4960 28262 4990 28314
rect 4990 28262 5002 28314
rect 5002 28262 5016 28314
rect 5040 28262 5054 28314
rect 5054 28262 5066 28314
rect 5066 28262 5096 28314
rect 5120 28262 5130 28314
rect 5130 28262 5176 28314
rect 4880 28260 4936 28262
rect 4960 28260 5016 28262
rect 5040 28260 5096 28262
rect 5120 28260 5176 28262
rect 4880 27226 4936 27228
rect 4960 27226 5016 27228
rect 5040 27226 5096 27228
rect 5120 27226 5176 27228
rect 4880 27174 4926 27226
rect 4926 27174 4936 27226
rect 4960 27174 4990 27226
rect 4990 27174 5002 27226
rect 5002 27174 5016 27226
rect 5040 27174 5054 27226
rect 5054 27174 5066 27226
rect 5066 27174 5096 27226
rect 5120 27174 5130 27226
rect 5130 27174 5176 27226
rect 4880 27172 4936 27174
rect 4960 27172 5016 27174
rect 5040 27172 5096 27174
rect 5120 27172 5176 27174
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4986 26424 5042 26480
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4880 26138 4936 26140
rect 4960 26138 5016 26140
rect 5040 26138 5096 26140
rect 5120 26138 5176 26140
rect 4880 26086 4926 26138
rect 4926 26086 4936 26138
rect 4960 26086 4990 26138
rect 4990 26086 5002 26138
rect 5002 26086 5016 26138
rect 5040 26086 5054 26138
rect 5054 26086 5066 26138
rect 5066 26086 5096 26138
rect 5120 26086 5130 26138
rect 5130 26086 5176 26138
rect 4880 26084 4936 26086
rect 4960 26084 5016 26086
rect 5040 26084 5096 26086
rect 5120 26084 5176 26086
rect 4880 25050 4936 25052
rect 4960 25050 5016 25052
rect 5040 25050 5096 25052
rect 5120 25050 5176 25052
rect 4880 24998 4926 25050
rect 4926 24998 4936 25050
rect 4960 24998 4990 25050
rect 4990 24998 5002 25050
rect 5002 24998 5016 25050
rect 5040 24998 5054 25050
rect 5054 24998 5066 25050
rect 5066 24998 5096 25050
rect 5120 24998 5130 25050
rect 5130 24998 5176 25050
rect 4880 24996 4936 24998
rect 4960 24996 5016 24998
rect 5040 24996 5096 24998
rect 5120 24996 5176 24998
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 1950 23160 2006 23216
rect 4880 23962 4936 23964
rect 4960 23962 5016 23964
rect 5040 23962 5096 23964
rect 5120 23962 5176 23964
rect 4880 23910 4926 23962
rect 4926 23910 4936 23962
rect 4960 23910 4990 23962
rect 4990 23910 5002 23962
rect 5002 23910 5016 23962
rect 5040 23910 5054 23962
rect 5054 23910 5066 23962
rect 5066 23910 5096 23962
rect 5120 23910 5130 23962
rect 5130 23910 5176 23962
rect 4880 23908 4936 23910
rect 4960 23908 5016 23910
rect 5040 23908 5096 23910
rect 5120 23908 5176 23910
rect 7102 26460 7104 26480
rect 7104 26460 7156 26480
rect 7156 26460 7158 26480
rect 7102 26424 7158 26460
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4880 22874 4936 22876
rect 4960 22874 5016 22876
rect 5040 22874 5096 22876
rect 5120 22874 5176 22876
rect 4880 22822 4926 22874
rect 4926 22822 4936 22874
rect 4960 22822 4990 22874
rect 4990 22822 5002 22874
rect 5002 22822 5016 22874
rect 5040 22822 5054 22874
rect 5054 22822 5066 22874
rect 5066 22822 5096 22874
rect 5120 22822 5130 22874
rect 5130 22822 5176 22874
rect 4880 22820 4936 22822
rect 4960 22820 5016 22822
rect 5040 22820 5096 22822
rect 5120 22820 5176 22822
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4880 21786 4936 21788
rect 4960 21786 5016 21788
rect 5040 21786 5096 21788
rect 5120 21786 5176 21788
rect 4880 21734 4926 21786
rect 4926 21734 4936 21786
rect 4960 21734 4990 21786
rect 4990 21734 5002 21786
rect 5002 21734 5016 21786
rect 5040 21734 5054 21786
rect 5054 21734 5066 21786
rect 5066 21734 5096 21786
rect 5120 21734 5130 21786
rect 5130 21734 5176 21786
rect 4880 21732 4936 21734
rect 4960 21732 5016 21734
rect 5040 21732 5096 21734
rect 5120 21732 5176 21734
rect 6826 21528 6882 21584
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 846 19896 902 19952
rect 4880 20698 4936 20700
rect 4960 20698 5016 20700
rect 5040 20698 5096 20700
rect 5120 20698 5176 20700
rect 4880 20646 4926 20698
rect 4926 20646 4936 20698
rect 4960 20646 4990 20698
rect 4990 20646 5002 20698
rect 5002 20646 5016 20698
rect 5040 20646 5054 20698
rect 5054 20646 5066 20698
rect 5066 20646 5096 20698
rect 5120 20646 5130 20698
rect 5130 20646 5176 20698
rect 4880 20644 4936 20646
rect 4960 20644 5016 20646
rect 5040 20644 5096 20646
rect 5120 20644 5176 20646
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4880 19610 4936 19612
rect 4960 19610 5016 19612
rect 5040 19610 5096 19612
rect 5120 19610 5176 19612
rect 4880 19558 4926 19610
rect 4926 19558 4936 19610
rect 4960 19558 4990 19610
rect 4990 19558 5002 19610
rect 5002 19558 5016 19610
rect 5040 19558 5054 19610
rect 5054 19558 5066 19610
rect 5066 19558 5096 19610
rect 5120 19558 5130 19610
rect 5130 19558 5176 19610
rect 4880 19556 4936 19558
rect 4960 19556 5016 19558
rect 5040 19556 5096 19558
rect 5120 19556 5176 19558
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4880 18522 4936 18524
rect 4960 18522 5016 18524
rect 5040 18522 5096 18524
rect 5120 18522 5176 18524
rect 4880 18470 4926 18522
rect 4926 18470 4936 18522
rect 4960 18470 4990 18522
rect 4990 18470 5002 18522
rect 5002 18470 5016 18522
rect 5040 18470 5054 18522
rect 5054 18470 5066 18522
rect 5066 18470 5096 18522
rect 5120 18470 5130 18522
rect 5130 18470 5176 18522
rect 4880 18468 4936 18470
rect 4960 18468 5016 18470
rect 5040 18468 5096 18470
rect 5120 18468 5176 18470
rect 7102 21548 7158 21584
rect 7102 21528 7104 21548
rect 7104 21528 7156 21548
rect 7156 21528 7158 21548
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4880 17434 4936 17436
rect 4960 17434 5016 17436
rect 5040 17434 5096 17436
rect 5120 17434 5176 17436
rect 4880 17382 4926 17434
rect 4926 17382 4936 17434
rect 4960 17382 4990 17434
rect 4990 17382 5002 17434
rect 5002 17382 5016 17434
rect 5040 17382 5054 17434
rect 5054 17382 5066 17434
rect 5066 17382 5096 17434
rect 5120 17382 5130 17434
rect 5130 17382 5176 17434
rect 4880 17380 4936 17382
rect 4960 17380 5016 17382
rect 5040 17380 5096 17382
rect 5120 17380 5176 17382
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4880 16346 4936 16348
rect 4960 16346 5016 16348
rect 5040 16346 5096 16348
rect 5120 16346 5176 16348
rect 4880 16294 4926 16346
rect 4926 16294 4936 16346
rect 4960 16294 4990 16346
rect 4990 16294 5002 16346
rect 5002 16294 5016 16346
rect 5040 16294 5054 16346
rect 5054 16294 5066 16346
rect 5066 16294 5096 16346
rect 5120 16294 5130 16346
rect 5130 16294 5176 16346
rect 4880 16292 4936 16294
rect 4960 16292 5016 16294
rect 5040 16292 5096 16294
rect 5120 16292 5176 16294
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4880 15258 4936 15260
rect 4960 15258 5016 15260
rect 5040 15258 5096 15260
rect 5120 15258 5176 15260
rect 4880 15206 4926 15258
rect 4926 15206 4936 15258
rect 4960 15206 4990 15258
rect 4990 15206 5002 15258
rect 5002 15206 5016 15258
rect 5040 15206 5054 15258
rect 5054 15206 5066 15258
rect 5066 15206 5096 15258
rect 5120 15206 5130 15258
rect 5130 15206 5176 15258
rect 4880 15204 4936 15206
rect 4960 15204 5016 15206
rect 5040 15204 5096 15206
rect 5120 15204 5176 15206
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4880 14170 4936 14172
rect 4960 14170 5016 14172
rect 5040 14170 5096 14172
rect 5120 14170 5176 14172
rect 4880 14118 4926 14170
rect 4926 14118 4936 14170
rect 4960 14118 4990 14170
rect 4990 14118 5002 14170
rect 5002 14118 5016 14170
rect 5040 14118 5054 14170
rect 5054 14118 5066 14170
rect 5066 14118 5096 14170
rect 5120 14118 5130 14170
rect 5130 14118 5176 14170
rect 4880 14116 4936 14118
rect 4960 14116 5016 14118
rect 5040 14116 5096 14118
rect 5120 14116 5176 14118
rect 4880 13082 4936 13084
rect 4960 13082 5016 13084
rect 5040 13082 5096 13084
rect 5120 13082 5176 13084
rect 4880 13030 4926 13082
rect 4926 13030 4936 13082
rect 4960 13030 4990 13082
rect 4990 13030 5002 13082
rect 5002 13030 5016 13082
rect 5040 13030 5054 13082
rect 5054 13030 5066 13082
rect 5066 13030 5096 13082
rect 5120 13030 5130 13082
rect 5130 13030 5176 13082
rect 4880 13028 4936 13030
rect 4960 13028 5016 13030
rect 5040 13028 5096 13030
rect 5120 13028 5176 13030
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 12162 21664 12218 21720
rect 12254 21548 12310 21584
rect 12254 21528 12256 21548
rect 12256 21528 12308 21548
rect 12308 21528 12310 21548
rect 10782 20476 10784 20496
rect 10784 20476 10836 20496
rect 10836 20476 10838 20496
rect 10782 20440 10838 20476
rect 5538 9424 5594 9480
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 5446 7792 5502 7848
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 6550 9424 6606 9480
rect 13082 21664 13138 21720
rect 12990 21528 13046 21584
rect 11334 15972 11390 16008
rect 11334 15952 11336 15972
rect 11336 15952 11388 15972
rect 11388 15952 11390 15972
rect 11150 15020 11206 15056
rect 11150 15000 11152 15020
rect 11152 15000 11204 15020
rect 11204 15000 11206 15020
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 13174 18964 13230 19000
rect 13174 18944 13176 18964
rect 13176 18944 13228 18964
rect 13228 18944 13230 18964
rect 14370 21120 14426 21176
rect 14186 20460 14242 20496
rect 14186 20440 14188 20460
rect 14188 20440 14240 20460
rect 14240 20440 14242 20460
rect 14186 19216 14242 19272
rect 13542 15136 13598 15192
rect 13450 15000 13506 15056
rect 13542 12844 13598 12880
rect 13542 12824 13544 12844
rect 13544 12824 13596 12844
rect 13596 12824 13598 12844
rect 15290 21564 15292 21584
rect 15292 21564 15344 21584
rect 15344 21564 15346 21584
rect 15290 21528 15346 21564
rect 15934 21800 15990 21856
rect 16026 20984 16082 21040
rect 17774 21936 17830 21992
rect 16302 20848 16358 20904
rect 17590 21800 17646 21856
rect 17038 21392 17094 21448
rect 18050 21836 18052 21856
rect 18052 21836 18104 21856
rect 18104 21836 18106 21856
rect 18050 21800 18106 21836
rect 19706 21800 19762 21856
rect 17774 20984 17830 21040
rect 18970 21120 19026 21176
rect 17866 20848 17922 20904
rect 17038 19216 17094 19272
rect 16394 18944 16450 19000
rect 15106 15952 15162 16008
rect 15106 15136 15162 15192
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 16670 17312 16726 17368
rect 15658 12860 15660 12880
rect 15660 12860 15712 12880
rect 15712 12860 15714 12880
rect 15658 12824 15714 12860
rect 12530 7812 12586 7848
rect 12530 7792 12532 7812
rect 12532 7792 12584 7812
rect 12584 7792 12586 7812
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 846 2932 848 2952
rect 848 2932 900 2952
rect 900 2932 902 2952
rect 846 2896 902 2932
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 17866 17312 17922 17368
rect 17498 15136 17554 15192
rect 20166 21548 20222 21584
rect 20166 21528 20168 21548
rect 20168 21528 20220 21548
rect 20220 21528 20222 21548
rect 19798 21392 19854 21448
rect 19338 13948 19340 13968
rect 19340 13948 19392 13968
rect 19392 13948 19394 13968
rect 19338 13912 19394 13948
rect 19430 13812 19432 13832
rect 19432 13812 19484 13832
rect 19484 13812 19486 13832
rect 19430 13776 19486 13812
rect 19338 13640 19394 13696
rect 19614 13640 19670 13696
rect 19890 13948 19892 13968
rect 19892 13948 19944 13968
rect 19944 13948 19946 13968
rect 19890 13912 19946 13948
rect 19798 13796 19854 13832
rect 19798 13776 19800 13796
rect 19800 13776 19852 13796
rect 19852 13776 19854 13796
rect 20994 21936 21050 21992
rect 17314 5516 17316 5536
rect 17316 5516 17368 5536
rect 17368 5516 17370 5536
rect 17314 5480 17370 5516
rect 15934 3984 15990 4040
rect 17958 5480 18014 5536
rect 20994 14864 21050 14920
rect 19982 3984 20038 4040
rect 22282 14884 22338 14920
rect 22282 14864 22284 14884
rect 22284 14864 22336 14884
rect 22336 14864 22338 14884
rect 23018 13932 23074 13968
rect 23018 13912 23020 13932
rect 23020 13912 23072 13932
rect 23072 13912 23074 13932
rect 23386 13932 23442 13968
rect 23386 13912 23388 13932
rect 23388 13912 23440 13932
rect 23440 13912 23442 13932
rect 23570 11636 23572 11656
rect 23572 11636 23624 11656
rect 23624 11636 23626 11656
rect 23570 11600 23626 11636
rect 25226 15272 25282 15328
rect 24398 5480 24454 5536
rect 25502 3984 25558 4040
rect 27526 2760 27582 2816
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
<< metal3 >>
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 4870 28320 5186 28321
rect 4870 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5186 28320
rect 4870 28255 5186 28256
rect 0 27978 800 28008
rect 1301 27978 1367 27981
rect 0 27976 1367 27978
rect 0 27920 1306 27976
rect 1362 27920 1367 27976
rect 0 27918 1367 27920
rect 0 27888 800 27918
rect 1301 27915 1367 27918
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 4870 27232 5186 27233
rect 4870 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5186 27232
rect 4870 27167 5186 27168
rect 4210 26688 4526 26689
rect 0 26618 800 26648
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 1209 26618 1275 26621
rect 0 26616 1275 26618
rect 0 26560 1214 26616
rect 1270 26560 1275 26616
rect 0 26558 1275 26560
rect 0 26528 800 26558
rect 1209 26555 1275 26558
rect 4981 26482 5047 26485
rect 7097 26482 7163 26485
rect 4981 26480 7163 26482
rect 4981 26424 4986 26480
rect 5042 26424 7102 26480
rect 7158 26424 7163 26480
rect 4981 26422 7163 26424
rect 4981 26419 5047 26422
rect 7097 26419 7163 26422
rect 4870 26144 5186 26145
rect 4870 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5186 26144
rect 4870 26079 5186 26080
rect 0 25938 800 25968
rect 1485 25938 1551 25941
rect 0 25936 1551 25938
rect 0 25880 1490 25936
rect 1546 25880 1551 25936
rect 0 25878 1551 25880
rect 0 25848 800 25878
rect 1485 25875 1551 25878
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 841 25394 907 25397
rect 798 25392 907 25394
rect 798 25336 846 25392
rect 902 25336 907 25392
rect 798 25331 907 25336
rect 798 25288 858 25331
rect 0 25198 858 25288
rect 0 25168 800 25198
rect 4870 25056 5186 25057
rect 4870 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5186 25056
rect 4870 24991 5186 24992
rect 841 24714 907 24717
rect 798 24712 907 24714
rect 798 24656 846 24712
rect 902 24656 907 24712
rect 798 24651 907 24656
rect 798 24608 858 24651
rect 0 24518 858 24608
rect 0 24488 800 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 4870 23968 5186 23969
rect 0 23898 800 23928
rect 4870 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5186 23968
rect 4870 23903 5186 23904
rect 1209 23898 1275 23901
rect 0 23896 1275 23898
rect 0 23840 1214 23896
rect 1270 23840 1275 23896
rect 0 23838 1275 23840
rect 0 23808 800 23838
rect 1209 23835 1275 23838
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 0 23218 800 23248
rect 1945 23218 2011 23221
rect 0 23216 2011 23218
rect 0 23160 1950 23216
rect 2006 23160 2011 23216
rect 0 23158 2011 23160
rect 0 23128 800 23158
rect 1945 23155 2011 23158
rect 4870 22880 5186 22881
rect 4870 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5186 22880
rect 4870 22815 5186 22816
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 17769 21994 17835 21997
rect 20989 21994 21055 21997
rect 17769 21992 21055 21994
rect 17769 21936 17774 21992
rect 17830 21936 20994 21992
rect 21050 21936 21055 21992
rect 17769 21934 21055 21936
rect 17769 21931 17835 21934
rect 20989 21931 21055 21934
rect 15929 21858 15995 21861
rect 17585 21858 17651 21861
rect 18045 21858 18111 21861
rect 19701 21858 19767 21861
rect 15929 21856 19767 21858
rect 15929 21800 15934 21856
rect 15990 21800 17590 21856
rect 17646 21800 18050 21856
rect 18106 21800 19706 21856
rect 19762 21800 19767 21856
rect 15929 21798 19767 21800
rect 15929 21795 15995 21798
rect 17585 21795 17651 21798
rect 18045 21795 18111 21798
rect 19701 21795 19767 21798
rect 4870 21792 5186 21793
rect 4870 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5186 21792
rect 4870 21727 5186 21728
rect 12157 21722 12223 21725
rect 13077 21722 13143 21725
rect 12157 21720 13143 21722
rect 12157 21664 12162 21720
rect 12218 21664 13082 21720
rect 13138 21664 13143 21720
rect 12157 21662 13143 21664
rect 12157 21659 12223 21662
rect 13077 21659 13143 21662
rect 6821 21586 6887 21589
rect 7097 21586 7163 21589
rect 6821 21584 7163 21586
rect 6821 21528 6826 21584
rect 6882 21528 7102 21584
rect 7158 21528 7163 21584
rect 6821 21526 7163 21528
rect 6821 21523 6887 21526
rect 7097 21523 7163 21526
rect 12249 21586 12315 21589
rect 12985 21586 13051 21589
rect 12249 21584 13051 21586
rect 12249 21528 12254 21584
rect 12310 21528 12990 21584
rect 13046 21528 13051 21584
rect 12249 21526 13051 21528
rect 12249 21523 12315 21526
rect 12985 21523 13051 21526
rect 15285 21586 15351 21589
rect 20161 21586 20227 21589
rect 15285 21584 20227 21586
rect 15285 21528 15290 21584
rect 15346 21528 20166 21584
rect 20222 21528 20227 21584
rect 15285 21526 20227 21528
rect 15285 21523 15351 21526
rect 20161 21523 20227 21526
rect 17033 21450 17099 21453
rect 19793 21450 19859 21453
rect 17033 21448 19859 21450
rect 17033 21392 17038 21448
rect 17094 21392 19798 21448
rect 19854 21392 19859 21448
rect 17033 21390 19859 21392
rect 17033 21387 17099 21390
rect 19793 21387 19859 21390
rect 841 21314 907 21317
rect 798 21312 907 21314
rect 798 21256 846 21312
rect 902 21256 907 21312
rect 798 21251 907 21256
rect 798 21208 858 21251
rect 0 21118 858 21208
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 14365 21178 14431 21181
rect 18965 21178 19031 21181
rect 14365 21176 19031 21178
rect 14365 21120 14370 21176
rect 14426 21120 18970 21176
rect 19026 21120 19031 21176
rect 14365 21118 19031 21120
rect 0 21088 800 21118
rect 14365 21115 14431 21118
rect 18965 21115 19031 21118
rect 16021 21042 16087 21045
rect 17769 21042 17835 21045
rect 16021 21040 17835 21042
rect 16021 20984 16026 21040
rect 16082 20984 17774 21040
rect 17830 20984 17835 21040
rect 16021 20982 17835 20984
rect 16021 20979 16087 20982
rect 17769 20979 17835 20982
rect 16297 20906 16363 20909
rect 17861 20906 17927 20909
rect 16297 20904 17927 20906
rect 16297 20848 16302 20904
rect 16358 20848 17866 20904
rect 17922 20848 17927 20904
rect 16297 20846 17927 20848
rect 16297 20843 16363 20846
rect 17861 20843 17927 20846
rect 4870 20704 5186 20705
rect 4870 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5186 20704
rect 4870 20639 5186 20640
rect 10777 20498 10843 20501
rect 14181 20498 14247 20501
rect 10777 20496 14247 20498
rect 10777 20440 10782 20496
rect 10838 20440 14186 20496
rect 14242 20440 14247 20496
rect 10777 20438 14247 20440
rect 10777 20435 10843 20438
rect 14181 20435 14247 20438
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 841 19954 907 19957
rect 798 19952 907 19954
rect 798 19896 846 19952
rect 902 19896 907 19952
rect 798 19891 907 19896
rect 798 19848 858 19891
rect 0 19758 858 19848
rect 0 19728 800 19758
rect 4870 19616 5186 19617
rect 4870 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5186 19616
rect 4870 19551 5186 19552
rect 14181 19274 14247 19277
rect 17033 19274 17099 19277
rect 14181 19272 17099 19274
rect 14181 19216 14186 19272
rect 14242 19216 17038 19272
rect 17094 19216 17099 19272
rect 14181 19214 17099 19216
rect 14181 19211 14247 19214
rect 17033 19211 17099 19214
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 13169 19002 13235 19005
rect 16389 19002 16455 19005
rect 13169 19000 16455 19002
rect 13169 18944 13174 19000
rect 13230 18944 16394 19000
rect 16450 18944 16455 19000
rect 13169 18942 16455 18944
rect 13169 18939 13235 18942
rect 16389 18939 16455 18942
rect 4870 18528 5186 18529
rect 4870 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5186 18528
rect 4870 18463 5186 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 4870 17440 5186 17441
rect 4870 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5186 17440
rect 4870 17375 5186 17376
rect 16665 17370 16731 17373
rect 17861 17370 17927 17373
rect 16665 17368 17927 17370
rect 16665 17312 16670 17368
rect 16726 17312 17866 17368
rect 17922 17312 17927 17368
rect 16665 17310 17927 17312
rect 16665 17307 16731 17310
rect 17861 17307 17927 17310
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 4870 16352 5186 16353
rect 4870 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5186 16352
rect 4870 16287 5186 16288
rect 11329 16010 11395 16013
rect 15101 16010 15167 16013
rect 11329 16008 15167 16010
rect 11329 15952 11334 16008
rect 11390 15952 15106 16008
rect 15162 15952 15167 16008
rect 11329 15950 15167 15952
rect 11329 15947 11395 15950
rect 15101 15947 15167 15950
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 25221 15330 25287 15333
rect 25630 15330 25636 15332
rect 25221 15328 25636 15330
rect 25221 15272 25226 15328
rect 25282 15272 25636 15328
rect 25221 15270 25636 15272
rect 25221 15267 25287 15270
rect 25630 15268 25636 15270
rect 25700 15268 25706 15332
rect 4870 15264 5186 15265
rect 4870 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5186 15264
rect 4870 15199 5186 15200
rect 13537 15194 13603 15197
rect 15101 15194 15167 15197
rect 17493 15194 17559 15197
rect 13537 15192 17559 15194
rect 13537 15136 13542 15192
rect 13598 15136 15106 15192
rect 15162 15136 17498 15192
rect 17554 15136 17559 15192
rect 13537 15134 17559 15136
rect 13537 15131 13603 15134
rect 15101 15131 15167 15134
rect 17493 15131 17559 15134
rect 11145 15058 11211 15061
rect 13445 15058 13511 15061
rect 11145 15056 13511 15058
rect 11145 15000 11150 15056
rect 11206 15000 13450 15056
rect 13506 15000 13511 15056
rect 11145 14998 13511 15000
rect 11145 14995 11211 14998
rect 13445 14995 13511 14998
rect 20989 14922 21055 14925
rect 22277 14922 22343 14925
rect 20989 14920 22343 14922
rect 20989 14864 20994 14920
rect 21050 14864 22282 14920
rect 22338 14864 22343 14920
rect 20989 14862 22343 14864
rect 20989 14859 21055 14862
rect 22277 14859 22343 14862
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 4870 14176 5186 14177
rect 4870 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5186 14176
rect 4870 14111 5186 14112
rect 19333 13970 19399 13973
rect 19885 13970 19951 13973
rect 19333 13968 19951 13970
rect 19333 13912 19338 13968
rect 19394 13912 19890 13968
rect 19946 13912 19951 13968
rect 19333 13910 19951 13912
rect 19333 13907 19399 13910
rect 19885 13907 19951 13910
rect 23013 13970 23079 13973
rect 23381 13970 23447 13973
rect 23013 13968 23447 13970
rect 23013 13912 23018 13968
rect 23074 13912 23386 13968
rect 23442 13912 23447 13968
rect 23013 13910 23447 13912
rect 23013 13907 23079 13910
rect 23381 13907 23447 13910
rect 19425 13834 19491 13837
rect 19793 13834 19859 13837
rect 19425 13832 19859 13834
rect 19425 13776 19430 13832
rect 19486 13776 19798 13832
rect 19854 13776 19859 13832
rect 19425 13774 19859 13776
rect 19425 13771 19491 13774
rect 19793 13771 19859 13774
rect 19333 13698 19399 13701
rect 19609 13698 19675 13701
rect 19333 13696 19675 13698
rect 19333 13640 19338 13696
rect 19394 13640 19614 13696
rect 19670 13640 19675 13696
rect 19333 13638 19675 13640
rect 19333 13635 19399 13638
rect 19609 13635 19675 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 4870 13088 5186 13089
rect 4870 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5186 13088
rect 4870 13023 5186 13024
rect 13537 12882 13603 12885
rect 15653 12882 15719 12885
rect 13537 12880 15719 12882
rect 13537 12824 13542 12880
rect 13598 12824 15658 12880
rect 15714 12824 15719 12880
rect 13537 12822 15719 12824
rect 13537 12819 13603 12822
rect 15653 12819 15719 12822
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 23565 11658 23631 11661
rect 23790 11658 23796 11660
rect 23565 11656 23796 11658
rect 23565 11600 23570 11656
rect 23626 11600 23796 11656
rect 23565 11598 23796 11600
rect 23565 11595 23631 11598
rect 23790 11596 23796 11598
rect 23860 11596 23866 11660
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 4870 10847 5186 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 5533 9482 5599 9485
rect 6545 9482 6611 9485
rect 5533 9480 6611 9482
rect 5533 9424 5538 9480
rect 5594 9424 6550 9480
rect 6606 9424 6611 9480
rect 5533 9422 6611 9424
rect 5533 9419 5599 9422
rect 6545 9419 6611 9422
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 5441 7850 5507 7853
rect 12525 7850 12591 7853
rect 5441 7848 12591 7850
rect 5441 7792 5446 7848
rect 5502 7792 12530 7848
rect 12586 7792 12591 7848
rect 5441 7790 12591 7792
rect 5441 7787 5507 7790
rect 12525 7787 12591 7790
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 17309 5538 17375 5541
rect 17953 5538 18019 5541
rect 17309 5536 18019 5538
rect 17309 5480 17314 5536
rect 17370 5480 17958 5536
rect 18014 5480 18019 5536
rect 17309 5478 18019 5480
rect 17309 5475 17375 5478
rect 17953 5475 18019 5478
rect 23790 5476 23796 5540
rect 23860 5538 23866 5540
rect 24393 5538 24459 5541
rect 23860 5536 24459 5538
rect 23860 5480 24398 5536
rect 24454 5480 24459 5536
rect 23860 5478 24459 5480
rect 23860 5476 23866 5478
rect 24393 5475 24459 5478
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 4870 5407 5186 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 15929 4042 15995 4045
rect 19977 4042 20043 4045
rect 15929 4040 20043 4042
rect 15929 3984 15934 4040
rect 15990 3984 19982 4040
rect 20038 3984 20043 4040
rect 15929 3982 20043 3984
rect 15929 3979 15995 3982
rect 19977 3979 20043 3982
rect 25497 4042 25563 4045
rect 25630 4042 25636 4044
rect 25497 4040 25636 4042
rect 25497 3984 25502 4040
rect 25558 3984 25636 4040
rect 25497 3982 25636 3984
rect 25497 3979 25563 3982
rect 25630 3980 25636 3982
rect 25700 3980 25706 4044
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 841 2954 907 2957
rect 798 2952 907 2954
rect 798 2896 846 2952
rect 902 2896 907 2952
rect 798 2891 907 2896
rect 798 2848 858 2891
rect 0 2758 858 2848
rect 27521 2818 27587 2821
rect 28220 2818 29020 2848
rect 27521 2816 29020 2818
rect 27521 2760 27526 2816
rect 27582 2760 29020 2816
rect 27521 2758 29020 2760
rect 0 2728 800 2758
rect 27521 2755 27587 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 28220 2728 29020 2758
rect 4210 2687 4526 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
<< via3 >>
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 4876 28316 4940 28320
rect 4876 28260 4880 28316
rect 4880 28260 4936 28316
rect 4936 28260 4940 28316
rect 4876 28256 4940 28260
rect 4956 28316 5020 28320
rect 4956 28260 4960 28316
rect 4960 28260 5016 28316
rect 5016 28260 5020 28316
rect 4956 28256 5020 28260
rect 5036 28316 5100 28320
rect 5036 28260 5040 28316
rect 5040 28260 5096 28316
rect 5096 28260 5100 28316
rect 5036 28256 5100 28260
rect 5116 28316 5180 28320
rect 5116 28260 5120 28316
rect 5120 28260 5176 28316
rect 5176 28260 5180 28316
rect 5116 28256 5180 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 4876 27228 4940 27232
rect 4876 27172 4880 27228
rect 4880 27172 4936 27228
rect 4936 27172 4940 27228
rect 4876 27168 4940 27172
rect 4956 27228 5020 27232
rect 4956 27172 4960 27228
rect 4960 27172 5016 27228
rect 5016 27172 5020 27228
rect 4956 27168 5020 27172
rect 5036 27228 5100 27232
rect 5036 27172 5040 27228
rect 5040 27172 5096 27228
rect 5096 27172 5100 27228
rect 5036 27168 5100 27172
rect 5116 27228 5180 27232
rect 5116 27172 5120 27228
rect 5120 27172 5176 27228
rect 5176 27172 5180 27228
rect 5116 27168 5180 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 4876 26140 4940 26144
rect 4876 26084 4880 26140
rect 4880 26084 4936 26140
rect 4936 26084 4940 26140
rect 4876 26080 4940 26084
rect 4956 26140 5020 26144
rect 4956 26084 4960 26140
rect 4960 26084 5016 26140
rect 5016 26084 5020 26140
rect 4956 26080 5020 26084
rect 5036 26140 5100 26144
rect 5036 26084 5040 26140
rect 5040 26084 5096 26140
rect 5096 26084 5100 26140
rect 5036 26080 5100 26084
rect 5116 26140 5180 26144
rect 5116 26084 5120 26140
rect 5120 26084 5176 26140
rect 5176 26084 5180 26140
rect 5116 26080 5180 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 4876 25052 4940 25056
rect 4876 24996 4880 25052
rect 4880 24996 4936 25052
rect 4936 24996 4940 25052
rect 4876 24992 4940 24996
rect 4956 25052 5020 25056
rect 4956 24996 4960 25052
rect 4960 24996 5016 25052
rect 5016 24996 5020 25052
rect 4956 24992 5020 24996
rect 5036 25052 5100 25056
rect 5036 24996 5040 25052
rect 5040 24996 5096 25052
rect 5096 24996 5100 25052
rect 5036 24992 5100 24996
rect 5116 25052 5180 25056
rect 5116 24996 5120 25052
rect 5120 24996 5176 25052
rect 5176 24996 5180 25052
rect 5116 24992 5180 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 4876 23964 4940 23968
rect 4876 23908 4880 23964
rect 4880 23908 4936 23964
rect 4936 23908 4940 23964
rect 4876 23904 4940 23908
rect 4956 23964 5020 23968
rect 4956 23908 4960 23964
rect 4960 23908 5016 23964
rect 5016 23908 5020 23964
rect 4956 23904 5020 23908
rect 5036 23964 5100 23968
rect 5036 23908 5040 23964
rect 5040 23908 5096 23964
rect 5096 23908 5100 23964
rect 5036 23904 5100 23908
rect 5116 23964 5180 23968
rect 5116 23908 5120 23964
rect 5120 23908 5176 23964
rect 5176 23908 5180 23964
rect 5116 23904 5180 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 4876 22876 4940 22880
rect 4876 22820 4880 22876
rect 4880 22820 4936 22876
rect 4936 22820 4940 22876
rect 4876 22816 4940 22820
rect 4956 22876 5020 22880
rect 4956 22820 4960 22876
rect 4960 22820 5016 22876
rect 5016 22820 5020 22876
rect 4956 22816 5020 22820
rect 5036 22876 5100 22880
rect 5036 22820 5040 22876
rect 5040 22820 5096 22876
rect 5096 22820 5100 22876
rect 5036 22816 5100 22820
rect 5116 22876 5180 22880
rect 5116 22820 5120 22876
rect 5120 22820 5176 22876
rect 5176 22820 5180 22876
rect 5116 22816 5180 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 4876 21788 4940 21792
rect 4876 21732 4880 21788
rect 4880 21732 4936 21788
rect 4936 21732 4940 21788
rect 4876 21728 4940 21732
rect 4956 21788 5020 21792
rect 4956 21732 4960 21788
rect 4960 21732 5016 21788
rect 5016 21732 5020 21788
rect 4956 21728 5020 21732
rect 5036 21788 5100 21792
rect 5036 21732 5040 21788
rect 5040 21732 5096 21788
rect 5096 21732 5100 21788
rect 5036 21728 5100 21732
rect 5116 21788 5180 21792
rect 5116 21732 5120 21788
rect 5120 21732 5176 21788
rect 5176 21732 5180 21788
rect 5116 21728 5180 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 4876 20700 4940 20704
rect 4876 20644 4880 20700
rect 4880 20644 4936 20700
rect 4936 20644 4940 20700
rect 4876 20640 4940 20644
rect 4956 20700 5020 20704
rect 4956 20644 4960 20700
rect 4960 20644 5016 20700
rect 5016 20644 5020 20700
rect 4956 20640 5020 20644
rect 5036 20700 5100 20704
rect 5036 20644 5040 20700
rect 5040 20644 5096 20700
rect 5096 20644 5100 20700
rect 5036 20640 5100 20644
rect 5116 20700 5180 20704
rect 5116 20644 5120 20700
rect 5120 20644 5176 20700
rect 5176 20644 5180 20700
rect 5116 20640 5180 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 4876 19612 4940 19616
rect 4876 19556 4880 19612
rect 4880 19556 4936 19612
rect 4936 19556 4940 19612
rect 4876 19552 4940 19556
rect 4956 19612 5020 19616
rect 4956 19556 4960 19612
rect 4960 19556 5016 19612
rect 5016 19556 5020 19612
rect 4956 19552 5020 19556
rect 5036 19612 5100 19616
rect 5036 19556 5040 19612
rect 5040 19556 5096 19612
rect 5096 19556 5100 19612
rect 5036 19552 5100 19556
rect 5116 19612 5180 19616
rect 5116 19556 5120 19612
rect 5120 19556 5176 19612
rect 5176 19556 5180 19612
rect 5116 19552 5180 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 4876 18524 4940 18528
rect 4876 18468 4880 18524
rect 4880 18468 4936 18524
rect 4936 18468 4940 18524
rect 4876 18464 4940 18468
rect 4956 18524 5020 18528
rect 4956 18468 4960 18524
rect 4960 18468 5016 18524
rect 5016 18468 5020 18524
rect 4956 18464 5020 18468
rect 5036 18524 5100 18528
rect 5036 18468 5040 18524
rect 5040 18468 5096 18524
rect 5096 18468 5100 18524
rect 5036 18464 5100 18468
rect 5116 18524 5180 18528
rect 5116 18468 5120 18524
rect 5120 18468 5176 18524
rect 5176 18468 5180 18524
rect 5116 18464 5180 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 4876 17436 4940 17440
rect 4876 17380 4880 17436
rect 4880 17380 4936 17436
rect 4936 17380 4940 17436
rect 4876 17376 4940 17380
rect 4956 17436 5020 17440
rect 4956 17380 4960 17436
rect 4960 17380 5016 17436
rect 5016 17380 5020 17436
rect 4956 17376 5020 17380
rect 5036 17436 5100 17440
rect 5036 17380 5040 17436
rect 5040 17380 5096 17436
rect 5096 17380 5100 17436
rect 5036 17376 5100 17380
rect 5116 17436 5180 17440
rect 5116 17380 5120 17436
rect 5120 17380 5176 17436
rect 5176 17380 5180 17436
rect 5116 17376 5180 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 4876 16348 4940 16352
rect 4876 16292 4880 16348
rect 4880 16292 4936 16348
rect 4936 16292 4940 16348
rect 4876 16288 4940 16292
rect 4956 16348 5020 16352
rect 4956 16292 4960 16348
rect 4960 16292 5016 16348
rect 5016 16292 5020 16348
rect 4956 16288 5020 16292
rect 5036 16348 5100 16352
rect 5036 16292 5040 16348
rect 5040 16292 5096 16348
rect 5096 16292 5100 16348
rect 5036 16288 5100 16292
rect 5116 16348 5180 16352
rect 5116 16292 5120 16348
rect 5120 16292 5176 16348
rect 5176 16292 5180 16348
rect 5116 16288 5180 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 25636 15268 25700 15332
rect 4876 15260 4940 15264
rect 4876 15204 4880 15260
rect 4880 15204 4936 15260
rect 4936 15204 4940 15260
rect 4876 15200 4940 15204
rect 4956 15260 5020 15264
rect 4956 15204 4960 15260
rect 4960 15204 5016 15260
rect 5016 15204 5020 15260
rect 4956 15200 5020 15204
rect 5036 15260 5100 15264
rect 5036 15204 5040 15260
rect 5040 15204 5096 15260
rect 5096 15204 5100 15260
rect 5036 15200 5100 15204
rect 5116 15260 5180 15264
rect 5116 15204 5120 15260
rect 5120 15204 5176 15260
rect 5176 15204 5180 15260
rect 5116 15200 5180 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 4876 14172 4940 14176
rect 4876 14116 4880 14172
rect 4880 14116 4936 14172
rect 4936 14116 4940 14172
rect 4876 14112 4940 14116
rect 4956 14172 5020 14176
rect 4956 14116 4960 14172
rect 4960 14116 5016 14172
rect 5016 14116 5020 14172
rect 4956 14112 5020 14116
rect 5036 14172 5100 14176
rect 5036 14116 5040 14172
rect 5040 14116 5096 14172
rect 5096 14116 5100 14172
rect 5036 14112 5100 14116
rect 5116 14172 5180 14176
rect 5116 14116 5120 14172
rect 5120 14116 5176 14172
rect 5176 14116 5180 14172
rect 5116 14112 5180 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 4876 13084 4940 13088
rect 4876 13028 4880 13084
rect 4880 13028 4936 13084
rect 4936 13028 4940 13084
rect 4876 13024 4940 13028
rect 4956 13084 5020 13088
rect 4956 13028 4960 13084
rect 4960 13028 5016 13084
rect 5016 13028 5020 13084
rect 4956 13024 5020 13028
rect 5036 13084 5100 13088
rect 5036 13028 5040 13084
rect 5040 13028 5096 13084
rect 5096 13028 5100 13084
rect 5036 13024 5100 13028
rect 5116 13084 5180 13088
rect 5116 13028 5120 13084
rect 5120 13028 5176 13084
rect 5176 13028 5180 13084
rect 5116 13024 5180 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 23796 11596 23860 11660
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 23796 5476 23860 5540
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 25636 3980 25700 4044
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
<< metal4 >>
rect 4208 28864 4528 28880
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 28320 5188 28880
rect 4868 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5188 28320
rect 4868 27232 5188 28256
rect 4868 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5188 27232
rect 4868 26144 5188 27168
rect 4868 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5188 26144
rect 4868 25056 5188 26080
rect 4868 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5188 25056
rect 4868 23968 5188 24992
rect 4868 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5188 23968
rect 4868 22880 5188 23904
rect 4868 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5188 22880
rect 4868 21792 5188 22816
rect 4868 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5188 21792
rect 4868 20704 5188 21728
rect 4868 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5188 20704
rect 4868 19616 5188 20640
rect 4868 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5188 19616
rect 4868 18528 5188 19552
rect 4868 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5188 18528
rect 4868 17440 5188 18464
rect 4868 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5188 17440
rect 4868 16352 5188 17376
rect 4868 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5188 16352
rect 4868 15264 5188 16288
rect 25635 15332 25701 15333
rect 25635 15268 25636 15332
rect 25700 15268 25701 15332
rect 25635 15267 25701 15268
rect 4868 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5188 15264
rect 4868 14176 5188 15200
rect 4868 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5188 14176
rect 4868 13088 5188 14112
rect 4868 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5188 13088
rect 4868 12000 5188 13024
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4868 10912 5188 11936
rect 23795 11660 23861 11661
rect 23795 11596 23796 11660
rect 23860 11596 23861 11660
rect 23795 11595 23861 11596
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 5472 5188 6496
rect 23798 5541 23858 11595
rect 23795 5540 23861 5541
rect 23795 5476 23796 5540
rect 23860 5476 23861 5540
rect 23795 5475 23861 5476
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 25638 4045 25698 15267
rect 25635 4044 25701 4045
rect 25635 3980 25636 4044
rect 25700 3980 25701 4044
rect 25635 3979 25701 3980
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
use sky130_fd_sc_hd__inv_2  _0787_
timestamp 1
transform -1 0 8556 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0788_
timestamp 1
transform 1 0 6808 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0789_
timestamp 1
transform 1 0 8096 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0790_
timestamp 1
transform -1 0 7268 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0791_
timestamp 1
transform -1 0 18860 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0792_
timestamp 1
transform 1 0 8924 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0793_
timestamp 1
transform 1 0 5152 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0794_
timestamp 1
transform 1 0 18216 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0795_
timestamp 1
transform 1 0 20792 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0796_
timestamp 1
transform 1 0 23644 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0797_
timestamp 1
transform -1 0 10120 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0798_
timestamp 1
transform -1 0 12052 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0799_
timestamp 1
transform -1 0 9476 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0800_
timestamp 1
transform -1 0 5336 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _0801_
timestamp 1
transform -1 0 2944 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _0802_
timestamp 1
transform 1 0 2944 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0803_
timestamp 1
transform -1 0 3128 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0804_
timestamp 1
transform 1 0 1656 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0805_
timestamp 1
transform 1 0 6348 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0806_
timestamp 1
transform -1 0 7452 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a2111o_1  _0807_
timestamp 1
transform 1 0 5336 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0808_
timestamp 1
transform -1 0 6808 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0809_
timestamp 1
transform -1 0 2024 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _0810_
timestamp 1
transform 1 0 7728 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a41o_1  _0811_
timestamp 1
transform 1 0 6164 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or4bb_1  _0812_
timestamp 1
transform 1 0 3220 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__or4bb_1  _0813_
timestamp 1
transform 1 0 3772 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0814_
timestamp 1
transform -1 0 4692 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0815_
timestamp 1
transform 1 0 3864 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0816_
timestamp 1
transform 1 0 3956 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0817_
timestamp 1
transform 1 0 4508 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0818_
timestamp 1
transform -1 0 6532 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0819_
timestamp 1
transform 1 0 5244 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0820_
timestamp 1
transform -1 0 6072 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0821_
timestamp 1
transform 1 0 5336 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o311a_1  _0822_
timestamp 1
transform 1 0 4600 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0823_
timestamp 1
transform 1 0 4048 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0824_
timestamp 1
transform -1 0 7636 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0825_
timestamp 1
transform -1 0 5980 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0826_
timestamp 1
transform -1 0 5336 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a211oi_1  _0827_
timestamp 1
transform -1 0 6624 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _0828_
timestamp 1
transform 1 0 3956 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_1  _0829_
timestamp 1
transform 1 0 4508 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0830_
timestamp 1
transform 1 0 4692 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _0831_
timestamp 1
transform -1 0 6256 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0832_
timestamp 1
transform 1 0 6532 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0833_
timestamp 1
transform 1 0 4692 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0834_
timestamp 1
transform 1 0 6348 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0835_
timestamp 1
transform 1 0 19228 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0836_
timestamp 1
transform 1 0 20700 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0837_
timestamp 1
transform -1 0 19688 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0838_
timestamp 1
transform 1 0 21160 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0839_
timestamp 1
transform -1 0 21252 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0840_
timestamp 1
transform -1 0 16468 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0841_
timestamp 1
transform 1 0 19596 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0842_
timestamp 1
transform -1 0 18584 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _0843_
timestamp 1
transform 1 0 12420 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _0844_
timestamp 1
transform 1 0 15456 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or4bb_1  _0845_
timestamp 1
transform 1 0 15732 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__or4_2  _0846_
timestamp 1
transform -1 0 16284 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0847_
timestamp 1
transform -1 0 17296 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0848_
timestamp 1
transform -1 0 16560 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0849_
timestamp 1
transform 1 0 16008 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0850_
timestamp 1
transform 1 0 17112 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0851_
timestamp 1
transform -1 0 17296 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0852_
timestamp 1
transform -1 0 17572 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0853_
timestamp 1
transform 1 0 17112 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0854_
timestamp 1
transform 1 0 16284 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0855_
timestamp 1
transform 1 0 15732 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0856_
timestamp 1
transform -1 0 16560 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0857_
timestamp 1
transform -1 0 15640 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0858_
timestamp 1
transform -1 0 15732 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_1  _0859_
timestamp 1
transform 1 0 13064 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0860_
timestamp 1
transform 1 0 14628 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0861_
timestamp 1
transform 1 0 14076 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0862_
timestamp 1
transform -1 0 14076 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0863_
timestamp 1
transform 1 0 13616 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0864_
timestamp 1
transform 1 0 13524 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0865_
timestamp 1
transform 1 0 14076 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0866_
timestamp 1
transform -1 0 13616 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0867_
timestamp 1
transform -1 0 13984 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0868_
timestamp 1
transform -1 0 12604 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0869_
timestamp 1
transform -1 0 13616 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0870_
timestamp 1
transform 1 0 12420 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0871_
timestamp 1
transform -1 0 13248 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0872_
timestamp 1
transform 1 0 13156 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0873_
timestamp 1
transform -1 0 11408 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0874_
timestamp 1
transform 1 0 10764 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0875_
timestamp 1
transform 1 0 6440 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0876_
timestamp 1
transform 1 0 7452 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0877_
timestamp 1
transform 1 0 11776 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0878_
timestamp 1
transform -1 0 10856 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _0879_
timestamp 1
transform 1 0 11684 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0880_
timestamp 1
transform -1 0 10488 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0881_
timestamp 1
transform 1 0 10120 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0882_
timestamp 1
transform 1 0 8096 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _0883_
timestamp 1
transform 1 0 11500 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0884_
timestamp 1
transform 1 0 14076 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0885_
timestamp 1
transform 1 0 3772 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0886_
timestamp 1
transform 1 0 4416 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0887_
timestamp 1
transform -1 0 4968 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0888_
timestamp 1
transform -1 0 13340 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0889_
timestamp 1
transform -1 0 9200 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0890_
timestamp 1
transform -1 0 11224 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0891_
timestamp 1
transform -1 0 12144 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _0892_
timestamp 1
transform -1 0 12236 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _0893_
timestamp 1
transform 1 0 11684 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0894_
timestamp 1
transform 1 0 12420 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0895_
timestamp 1
transform -1 0 11684 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _0896_
timestamp 1
transform -1 0 12604 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _0897_
timestamp 1
transform 1 0 11132 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _0898_
timestamp 1
transform 1 0 10396 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_1  _0899_
timestamp 1
transform 1 0 10120 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _0900_
timestamp 1
transform -1 0 10212 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0901_
timestamp 1
transform 1 0 7728 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0902_
timestamp 1
transform -1 0 5980 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _0903_
timestamp 1
transform 1 0 4968 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0904_
timestamp 1
transform 1 0 7360 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0905_
timestamp 1
transform 1 0 7084 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _0906_
timestamp 1
transform 1 0 6348 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a31oi_1  _0907_
timestamp 1
transform 1 0 5244 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0908_
timestamp 1
transform 1 0 6072 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0909_
timestamp 1
transform -1 0 6992 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0910_
timestamp 1
transform -1 0 5888 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0911_
timestamp 1
transform 1 0 6348 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0912_
timestamp 1
transform -1 0 7636 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0913_
timestamp 1
transform 1 0 5612 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0914_
timestamp 1
transform 1 0 6440 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0915_
timestamp 1
transform 1 0 5428 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _0916_
timestamp 1
transform 1 0 9568 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0917_
timestamp 1
transform 1 0 10856 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_1  _0918_
timestamp 1
transform 1 0 13064 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _0919_
timestamp 1
transform -1 0 13616 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _0920_
timestamp 1
transform -1 0 13616 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0921_
timestamp 1
transform 1 0 11684 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0922_
timestamp 1
transform -1 0 8740 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a2111o_1  _0923_
timestamp 1
transform 1 0 9936 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _0924_
timestamp 1
transform -1 0 9936 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0925_
timestamp 1
transform 1 0 6348 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0926_
timestamp 1
transform -1 0 4692 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0927_
timestamp 1
transform 1 0 9752 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0928_
timestamp 1
transform -1 0 19044 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0929_
timestamp 1
transform -1 0 9200 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0930_
timestamp 1
transform 1 0 8740 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0931_
timestamp 1
transform -1 0 10488 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0932_
timestamp 1
transform 1 0 9384 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0933_
timestamp 1
transform 1 0 8832 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0934_
timestamp 1
transform 1 0 10212 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0935_
timestamp 1
transform 1 0 9844 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0936_
timestamp 1
transform -1 0 11408 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0937_
timestamp 1
transform 1 0 10304 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0938_
timestamp 1
transform 1 0 11684 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0939_
timestamp 1
transform 1 0 12236 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0940_
timestamp 1
transform -1 0 11684 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0941_
timestamp 1
transform 1 0 11868 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0942_
timestamp 1
transform -1 0 12880 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0943_
timestamp 1
transform -1 0 13340 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0944_
timestamp 1
transform -1 0 13064 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0945_
timestamp 1
transform 1 0 13340 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0946_
timestamp 1
transform -1 0 3496 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0947_
timestamp 1
transform -1 0 5520 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0948_
timestamp 1
transform 1 0 3864 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0949_
timestamp 1
transform 1 0 5520 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _0950_
timestamp 1
transform -1 0 11316 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0951_
timestamp 1
transform 1 0 15456 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0952_
timestamp 1
transform -1 0 10672 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0953_
timestamp 1
transform 1 0 7636 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a41oi_4  _0954_
timestamp 1
transform 1 0 3956 0 -1 16320
box -38 -48 2062 592
use sky130_fd_sc_hd__a41o_1  _0955_
timestamp 1
transform 1 0 4140 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0956_
timestamp 1
transform 1 0 11224 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0957_
timestamp 1
transform 1 0 10304 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0958_
timestamp 1
transform -1 0 10672 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0959_
timestamp 1
transform 1 0 10028 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0960_
timestamp 1
transform 1 0 9476 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _0961_
timestamp 1
transform -1 0 10120 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0962_
timestamp 1
transform -1 0 9200 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0963_
timestamp 1
transform -1 0 10396 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0964_
timestamp 1
transform -1 0 9752 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0965_
timestamp 1
transform -1 0 10028 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0966_
timestamp 1
transform -1 0 9660 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0967_
timestamp 1
transform -1 0 9200 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0968_
timestamp 1
transform -1 0 9200 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0969_
timestamp 1
transform 1 0 8004 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0970_
timestamp 1
transform -1 0 8464 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0971_
timestamp 1
transform 1 0 8188 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0972_
timestamp 1
transform -1 0 8740 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0973_
timestamp 1
transform 1 0 6900 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0974_
timestamp 1
transform -1 0 6900 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0975_
timestamp 1
transform 1 0 8188 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _0976_
timestamp 1
transform 1 0 7176 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0977_
timestamp 1
transform 1 0 6440 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_4  _0978_
timestamp 1
transform -1 0 8372 0 -1 15232
box -38 -48 2062 592
use sky130_fd_sc_hd__nor2_1  _0979_
timestamp 1
transform 1 0 8004 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0980_
timestamp 1
transform 1 0 8280 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _0981_
timestamp 1
transform 1 0 8372 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _0982_
timestamp 1
transform -1 0 8004 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _0983_
timestamp 1
transform -1 0 7820 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0984_
timestamp 1
transform -1 0 7360 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a2111o_1  _0985_
timestamp 1
transform 1 0 7820 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _0986_
timestamp 1
transform 1 0 7360 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0987_
timestamp 1
transform -1 0 11868 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0988_
timestamp 1
transform -1 0 10856 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _0989_
timestamp 1
transform 1 0 10948 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0990_
timestamp 1
transform -1 0 11224 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0991_
timestamp 1
transform 1 0 10488 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _0992_
timestamp 1
transform 1 0 9844 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0993_
timestamp 1
transform -1 0 8464 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0994_
timestamp 1
transform -1 0 5796 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0995_
timestamp 1
transform 1 0 6992 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0996_
timestamp 1
transform 1 0 3680 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0997_
timestamp 1
transform -1 0 4048 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0998_
timestamp 1
transform 1 0 2944 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0999_
timestamp 1
transform -1 0 4600 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _1000_
timestamp 1
transform 1 0 3772 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1001_
timestamp 1
transform -1 0 3956 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1002_
timestamp 1
transform -1 0 6256 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1003_
timestamp 1
transform 1 0 5704 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _1004_
timestamp 1
transform -1 0 6624 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2b_1  _1005_
timestamp 1
transform -1 0 5612 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_2  _1006_
timestamp 1
transform 1 0 3404 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1007_
timestamp 1
transform 1 0 4600 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _1008_
timestamp 1
transform -1 0 4416 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1009_
timestamp 1
transform 1 0 5704 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1010_
timestamp 1
transform -1 0 6900 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _1011_
timestamp 1
transform 1 0 5612 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _1012_
timestamp 1
transform 1 0 4416 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1013_
timestamp 1
transform -1 0 4968 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a2111o_4  _1014_
timestamp 1
transform 1 0 4692 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__and3_1  _1015_
timestamp 1
transform 1 0 4048 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a221oi_4  _1016_
timestamp 1
transform 1 0 4508 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__and2_2  _1017_
timestamp 1
transform -1 0 5704 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1018_
timestamp 1
transform -1 0 5704 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1019_
timestamp 1
transform -1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1020_
timestamp 1
transform -1 0 12696 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1021_
timestamp 1
transform 1 0 11960 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1022_
timestamp 1
transform 1 0 12420 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_4  _1023_
timestamp 1
transform 1 0 10304 0 1 9792
box -38 -48 2062 592
use sky130_fd_sc_hd__nor2_1  _1024_
timestamp 1
transform -1 0 12788 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1025_
timestamp 1
transform -1 0 8464 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1026_
timestamp 1
transform -1 0 8280 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1027_
timestamp 1
transform 1 0 7360 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1028_
timestamp 1
transform -1 0 6900 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a221oi_4  _1029_
timestamp 1
transform 1 0 6348 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__xnor2_2  _1030_
timestamp 1
transform -1 0 7544 0 -1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1031_
timestamp 1
transform 1 0 6624 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _1032_
timestamp 1
transform 1 0 6348 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__a21boi_1  _1033_
timestamp 1
transform 1 0 6348 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _1034_
timestamp 1
transform 1 0 6348 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _1035_
timestamp 1
transform 1 0 7728 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1036_
timestamp 1
transform -1 0 7544 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__or3_2  _1037_
timestamp 1
transform -1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _1038_
timestamp 1
transform 1 0 7176 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_1  _1039_
timestamp 1
transform 1 0 7176 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_2  _1040_
timestamp 1
transform 1 0 8740 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_2  _1041_
timestamp 1
transform 1 0 8924 0 1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1042_
timestamp 1
transform 1 0 9936 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1043_
timestamp 1
transform -1 0 11408 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1044_
timestamp 1
transform 1 0 9752 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_2  _1045_
timestamp 1
transform 1 0 9752 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _1046_
timestamp 1
transform 1 0 9292 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1047_
timestamp 1
transform 1 0 8924 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1048_
timestamp 1
transform 1 0 9108 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1049_
timestamp 1
transform 1 0 7544 0 -1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1050_
timestamp 1
transform -1 0 8832 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor3b_1  _1051_
timestamp 1
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1052_
timestamp 1
transform 1 0 9476 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1053_
timestamp 1
transform 1 0 7176 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1054_
timestamp 1
transform 1 0 10396 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1055_
timestamp 1
transform 1 0 11592 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _1056_
timestamp 1
transform -1 0 10580 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1057_
timestamp 1
transform -1 0 9200 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand4b_1  _1058_
timestamp 1
transform 1 0 7544 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1059_
timestamp 1
transform -1 0 6624 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1060_
timestamp 1
transform -1 0 6532 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1061_
timestamp 1
transform 1 0 5060 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1062_
timestamp 1
transform -1 0 5980 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1063_
timestamp 1
transform 1 0 5060 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1064_
timestamp 1
transform 1 0 6348 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_2  _1065_
timestamp 1
transform 1 0 5060 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _1066_
timestamp 1
transform -1 0 6164 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a311o_1  _1067_
timestamp 1
transform -1 0 6256 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1068_
timestamp 1
transform 1 0 4784 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1069_
timestamp 1
transform -1 0 5152 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1070_
timestamp 1
transform 1 0 4232 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1071_
timestamp 1
transform -1 0 3864 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1072_
timestamp 1
transform 1 0 3864 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1073_
timestamp 1
transform 1 0 3772 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1074_
timestamp 1
transform -1 0 4692 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1075_
timestamp 1
transform 1 0 3312 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1076_
timestamp 1
transform 1 0 4324 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1077_
timestamp 1
transform 1 0 4232 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_2  _1078_
timestamp 1
transform 1 0 3036 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_2  _1079_
timestamp 1
transform 1 0 6348 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1080_
timestamp 1
transform -1 0 13156 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1081_
timestamp 1
transform 1 0 12144 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1082_
timestamp 1
transform 1 0 12788 0 1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__a21o_1  _1083_
timestamp 1
transform -1 0 12880 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_4  _1084_
timestamp 1
transform 1 0 12512 0 -1 9792
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_4  _1085_
timestamp 1
transform 1 0 11960 0 -1 8704
box -38 -48 2062 592
use sky130_fd_sc_hd__nor2_1  _1086_
timestamp 1
transform 1 0 13984 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1087_
timestamp 1
transform -1 0 4968 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_2  _1088_
timestamp 1
transform 1 0 5060 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _1089_
timestamp 1
transform 1 0 4784 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _1090_
timestamp 1
transform 1 0 4968 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1091_
timestamp 1
transform 1 0 4600 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1092_
timestamp 1
transform -1 0 5888 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1093_
timestamp 1
transform -1 0 6256 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1094_
timestamp 1
transform -1 0 6992 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1095_
timestamp 1
transform 1 0 4416 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _1096_
timestamp 1
transform 1 0 5244 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1097_
timestamp 1
transform -1 0 10764 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1098_
timestamp 1
transform 1 0 11040 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1099_
timestamp 1
transform -1 0 10948 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1100_
timestamp 1
transform 1 0 10764 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1101_
timestamp 1
transform 1 0 10120 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1102_
timestamp 1
transform 1 0 9384 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1103_
timestamp 1
transform 1 0 8832 0 -1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_1  _1104_
timestamp 1
transform -1 0 11408 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_2  _1105_
timestamp 1
transform 1 0 10948 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _1106_
timestamp 1
transform 1 0 11500 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1107_
timestamp 1
transform 1 0 12696 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_4  _1108_
timestamp 1
transform -1 0 16100 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__xnor2_1  _1109_
timestamp 1
transform 1 0 10120 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1110_
timestamp 1
transform -1 0 11316 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_2  _1111_
timestamp 1
transform 1 0 11500 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_1  _1112_
timestamp 1
transform -1 0 13524 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _1113_
timestamp 1
transform -1 0 8556 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1114_
timestamp 1
transform -1 0 8832 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _1115_
timestamp 1
transform 1 0 7360 0 1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__a22o_1  _1116_
timestamp 1
transform 1 0 8280 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1117_
timestamp 1
transform 1 0 8924 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__and2b_1  _1118_
timestamp 1
transform 1 0 10764 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1119_
timestamp 1
transform -1 0 12880 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _1120_
timestamp 1
transform 1 0 11868 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1121_
timestamp 1
transform 1 0 11776 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _1122_
timestamp 1
transform -1 0 12972 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1123_
timestamp 1
transform -1 0 12328 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1124_
timestamp 1
transform -1 0 11960 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1125_
timestamp 1
transform 1 0 5980 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1126_
timestamp 1
transform 1 0 5980 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1127_
timestamp 1
transform 1 0 6348 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1128_
timestamp 1
transform -1 0 10028 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1129_
timestamp 1
transform 1 0 10672 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _1130_
timestamp 1
transform 1 0 11224 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _1131_
timestamp 1
transform -1 0 12236 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1132_
timestamp 1
transform 1 0 11500 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1133_
timestamp 1
transform 1 0 12512 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a31oi_2  _1134_
timestamp 1
transform 1 0 12972 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _1135_
timestamp 1
transform 1 0 14076 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _1136_
timestamp 1
transform 1 0 13340 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _1137_
timestamp 1
transform -1 0 10672 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1138_
timestamp 1
transform -1 0 12144 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1139_
timestamp 1
transform -1 0 12696 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1140_
timestamp 1
transform 1 0 11776 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1141_
timestamp 1
transform -1 0 10488 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1142_
timestamp 1
transform -1 0 11316 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1143_
timestamp 1
transform 1 0 10212 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1144_
timestamp 1
transform 1 0 13432 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_4  _1145_
timestamp 1
transform 1 0 12788 0 -1 3264
box -38 -48 2062 592
use sky130_fd_sc_hd__a32oi_4  _1146_
timestamp 1
transform -1 0 16100 0 1 3264
box -38 -48 2062 592
use sky130_fd_sc_hd__a21oi_1  _1147_
timestamp 1
transform -1 0 13340 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1148_
timestamp 1
transform 1 0 13800 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1149_
timestamp 1
transform 1 0 14444 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1150_
timestamp 1
transform 1 0 13340 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _1151_
timestamp 1
transform -1 0 14996 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1152_
timestamp 1
transform -1 0 13708 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_2  _1153_
timestamp 1
transform 1 0 14904 0 1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _1154_
timestamp 1
transform 1 0 14260 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1155_
timestamp 1
transform 1 0 14168 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _1156_
timestamp 1
transform 1 0 14812 0 -1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _1157_
timestamp 1
transform -1 0 16836 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1158_
timestamp 1
transform 1 0 16008 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1159_
timestamp 1
transform 1 0 15180 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1160_
timestamp 1
transform 1 0 15456 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1161_
timestamp 1
transform 1 0 16008 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _1162_
timestamp 1
transform 1 0 14260 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1163_
timestamp 1
transform 1 0 14168 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _1164_
timestamp 1
transform 1 0 14628 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1165_
timestamp 1
transform -1 0 18216 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1166_
timestamp 1
transform 1 0 16652 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1167_
timestamp 1
transform 1 0 14996 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1168_
timestamp 1
transform 1 0 15088 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _1169_
timestamp 1
transform -1 0 16192 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1170_
timestamp 1
transform 1 0 16192 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1171_
timestamp 1
transform -1 0 16928 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1172_
timestamp 1
transform 1 0 15640 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1173_
timestamp 1
transform -1 0 14076 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1174_
timestamp 1
transform -1 0 13432 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1175_
timestamp 1
transform 1 0 12328 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1176_
timestamp 1
transform 1 0 14260 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _1177_
timestamp 1
transform 1 0 14812 0 -1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_1  _1178_
timestamp 1
transform 1 0 14076 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1179_
timestamp 1
transform 1 0 16284 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1180_
timestamp 1
transform -1 0 16560 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1181_
timestamp 1
transform 1 0 15456 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1182_
timestamp 1
transform 1 0 9568 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1183_
timestamp 1
transform -1 0 9568 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_2  _1184_
timestamp 1
transform 1 0 8924 0 1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _1185_
timestamp 1
transform 1 0 15640 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1186_
timestamp 1
transform 1 0 16008 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _1187_
timestamp 1
transform 1 0 13524 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1188_
timestamp 1
transform -1 0 15824 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1189_
timestamp 1
transform -1 0 17388 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1190_
timestamp 1
transform -1 0 17940 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1191_
timestamp 1
transform 1 0 16100 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1192_
timestamp 1
transform 1 0 16836 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1193_
timestamp 1
transform 1 0 16468 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__and3_1  _1194_
timestamp 1
transform 1 0 16744 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1195_
timestamp 1
transform -1 0 17940 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _1196_
timestamp 1
transform 1 0 18584 0 -1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_1  _1197_
timestamp 1
transform 1 0 19780 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1198_
timestamp 1
transform 1 0 17388 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1199_
timestamp 1
transform 1 0 17940 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _1200_
timestamp 1
transform -1 0 17940 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _1201_
timestamp 1
transform -1 0 17940 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1202_
timestamp 1
transform -1 0 17296 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1203_
timestamp 1
transform 1 0 17940 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1204_
timestamp 1
transform 1 0 21436 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1205_
timestamp 1
transform 1 0 16836 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1206_
timestamp 1
transform 1 0 15088 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _1207_
timestamp 1
transform 1 0 14812 0 -1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _1208_
timestamp 1
transform -1 0 20056 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1209_
timestamp 1
transform -1 0 17940 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _1210_
timestamp 1
transform -1 0 17664 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1211_
timestamp 1
transform 1 0 19228 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _1212_
timestamp 1
transform 1 0 17940 0 -1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__nand3_1  _1213_
timestamp 1
transform -1 0 19044 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1214_
timestamp 1
transform -1 0 18124 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1215_
timestamp 1
transform 1 0 17020 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1216_
timestamp 1
transform 1 0 17664 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_2  _1217_
timestamp 1
transform 1 0 17480 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_4  _1218_
timestamp 1
transform 1 0 18124 0 -1 8704
box -38 -48 2062 592
use sky130_fd_sc_hd__or2_1  _1219_
timestamp 1
transform -1 0 19872 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a22oi_2  _1220_
timestamp 1
transform 1 0 16744 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _1221_
timestamp 1
transform 1 0 21620 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _1222_
timestamp 1
transform -1 0 20424 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_2  _1223_
timestamp 1
transform 1 0 19780 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _1224_
timestamp 1
transform 1 0 17480 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1225_
timestamp 1
transform 1 0 16836 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1226_
timestamp 1
transform 1 0 17940 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _1227_
timestamp 1
transform 1 0 17204 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1228_
timestamp 1
transform 1 0 17940 0 1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__and3_1  _1229_
timestamp 1
transform 1 0 17756 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1230_
timestamp 1
transform 1 0 18584 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1231_
timestamp 1
transform 1 0 19228 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1232_
timestamp 1
transform 1 0 19412 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1233_
timestamp 1
transform 1 0 19964 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a22oi_2  _1234_
timestamp 1
transform 1 0 16836 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _1235_
timestamp 1
transform -1 0 20056 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1236_
timestamp 1
transform 1 0 21160 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1237_
timestamp 1
transform -1 0 21160 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _1238_
timestamp 1
transform -1 0 21252 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1239_
timestamp 1
transform 1 0 20056 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1240_
timestamp 1
transform 1 0 17940 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1241_
timestamp 1
transform 1 0 16192 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1242_
timestamp 1
transform 1 0 21068 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1243_
timestamp 1
transform 1 0 20608 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1244_
timestamp 1
transform -1 0 21528 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1245_
timestamp 1
transform -1 0 20884 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__o2111a_1  _1246_
timestamp 1
transform 1 0 19780 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__o2111ai_4  _1247_
timestamp 1
transform 1 0 19780 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__nor2_1  _1248_
timestamp 1
transform 1 0 21528 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _1249_
timestamp 1
transform 1 0 21804 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1250_
timestamp 1
transform 1 0 19504 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _1251_
timestamp 1
transform 1 0 19964 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__or4_1  _1252_
timestamp 1
transform 1 0 21344 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_1  _1253_
timestamp 1
transform 1 0 20792 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1254_
timestamp 1
transform 1 0 21804 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1255_
timestamp 1
transform 1 0 20424 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a31oi_2  _1256_
timestamp 1
transform -1 0 20516 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__a21oi_1  _1257_
timestamp 1
transform 1 0 22080 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1258_
timestamp 1
transform -1 0 21436 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1259_
timestamp 1
transform -1 0 21804 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1260_
timestamp 1
transform -1 0 21712 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o31ai_1  _1261_
timestamp 1
transform 1 0 19504 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1262_
timestamp 1
transform 1 0 20056 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1263_
timestamp 1
transform -1 0 21436 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1264_
timestamp 1
transform -1 0 21160 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1265_
timestamp 1
transform 1 0 20608 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1266_
timestamp 1
transform 1 0 20884 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1267_
timestamp 1
transform 1 0 23000 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1268_
timestamp 1
transform -1 0 24012 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1269_
timestamp 1
transform 1 0 21896 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o311a_2  _1270_
timestamp 1
transform -1 0 23092 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1271_
timestamp 1
transform -1 0 20700 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1272_
timestamp 1
transform 1 0 20608 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _1273_
timestamp 1
transform 1 0 21068 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1274_
timestamp 1
transform 1 0 21252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1275_
timestamp 1
transform -1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1276_
timestamp 1
transform -1 0 19044 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1277_
timestamp 1
transform -1 0 21620 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1278_
timestamp 1
transform 1 0 21896 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1279_
timestamp 1
transform 1 0 23736 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1280_
timestamp 1
transform 1 0 26128 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1281_
timestamp 1
transform 1 0 22540 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1282_
timestamp 1
transform -1 0 22448 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1283_
timestamp 1
transform 1 0 21896 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1284_
timestamp 1
transform -1 0 23736 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1285_
timestamp 1
transform 1 0 25300 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_4  _1286_
timestamp 1
transform 1 0 22632 0 -1 8704
box -38 -48 2062 592
use sky130_fd_sc_hd__o41a_1  _1287_
timestamp 1
transform -1 0 22632 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a21boi_1  _1288_
timestamp 1
transform 1 0 22356 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1289_
timestamp 1
transform -1 0 24288 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1290_
timestamp 1
transform 1 0 21804 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_4  _1291_
timestamp 1
transform 1 0 18860 0 -1 7616
box -38 -48 2062 592
use sky130_fd_sc_hd__or2_1  _1292_
timestamp 1
transform 1 0 20700 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_2  _1293_
timestamp 1
transform 1 0 20884 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1294_
timestamp 1
transform 1 0 23920 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1295_
timestamp 1
transform 1 0 22816 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _1296_
timestamp 1
transform 1 0 23276 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _1297_
timestamp 1
transform -1 0 22816 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o2111a_1  _1298_
timestamp 1
transform 1 0 23368 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _1299_
timestamp 1
transform 1 0 23092 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _1300_
timestamp 1
transform 1 0 23552 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1301_
timestamp 1
transform 1 0 23644 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1302_
timestamp 1
transform -1 0 22632 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_1  _1303_
timestamp 1
transform 1 0 21804 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _1304_
timestamp 1
transform 1 0 21436 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1305_
timestamp 1
transform 1 0 22540 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1306_
timestamp 1
transform 1 0 22172 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1307_
timestamp 1
transform 1 0 22816 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1308_
timestamp 1
transform -1 0 23920 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1309_
timestamp 1
transform -1 0 23644 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1310_
timestamp 1
transform 1 0 23000 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1311_
timestamp 1
transform 1 0 24472 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1312_
timestamp 1
transform -1 0 25484 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o22ai_2  _1313_
timestamp 1
transform 1 0 24380 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__o21a_1  _1314_
timestamp 1
transform -1 0 24564 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _1315_
timestamp 1
transform 1 0 24840 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _1316_
timestamp 1
transform -1 0 25392 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1317_
timestamp 1
transform -1 0 25944 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1318_
timestamp 1
transform 1 0 24840 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1319_
timestamp 1
transform 1 0 25484 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1320_
timestamp 1
transform 1 0 26220 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1321_
timestamp 1
transform -1 0 25576 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _1322_
timestamp 1
transform 1 0 23276 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1323_
timestamp 1
transform 1 0 23460 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1324_
timestamp 1
transform 1 0 23276 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1325_
timestamp 1
transform 1 0 24380 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1326_
timestamp 1
transform -1 0 25944 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1327_
timestamp 1
transform -1 0 25300 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1328_
timestamp 1
transform 1 0 22172 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1329_
timestamp 1
transform -1 0 22172 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1330_
timestamp 1
transform 1 0 23920 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _1331_
timestamp 1
transform 1 0 23552 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1332_
timestamp 1
transform 1 0 24288 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _1333_
timestamp 1
transform 1 0 24564 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_1  _1334_
timestamp 1
transform 1 0 24932 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _1335_
timestamp 1
transform 1 0 24380 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_2  _1336_
timestamp 1
transform 1 0 22356 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _1337_
timestamp 1
transform 1 0 25300 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1338_
timestamp 1
transform 1 0 24380 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _1339_
timestamp 1
transform -1 0 24932 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _1340_
timestamp 1
transform -1 0 23184 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1341_
timestamp 1
transform -1 0 23644 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1342_
timestamp 1
transform 1 0 22632 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1343_
timestamp 1
transform 1 0 22632 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _1344_
timestamp 1
transform 1 0 21804 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1345_
timestamp 1
transform 1 0 23552 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_2  _1346_
timestamp 1
transform 1 0 20516 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _1347_
timestamp 1
transform 1 0 22264 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__and3_1  _1348_
timestamp 1
transform 1 0 22908 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1349_
timestamp 1
transform 1 0 24288 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1350_
timestamp 1
transform 1 0 22908 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1351_
timestamp 1
transform -1 0 24104 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1352_
timestamp 1
transform 1 0 24748 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1353_
timestamp 1
transform -1 0 25300 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1354_
timestamp 1
transform -1 0 25300 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _1355_
timestamp 1
transform 1 0 25024 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1356_
timestamp 1
transform 1 0 25760 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1357_
timestamp 1
transform -1 0 27416 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1358_
timestamp 1
transform 1 0 25944 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1359_
timestamp 1
transform 1 0 25392 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1360_
timestamp 1
transform -1 0 26588 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1361_
timestamp 1
transform 1 0 24748 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1362_
timestamp 1
transform 1 0 24288 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1363_
timestamp 1
transform 1 0 24656 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1364_
timestamp 1
transform -1 0 26036 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1365_
timestamp 1
transform 1 0 26404 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1366_
timestamp 1
transform -1 0 26404 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1367_
timestamp 1
transform 1 0 26312 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _1368_
timestamp 1
transform -1 0 27232 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1369_
timestamp 1
transform -1 0 20148 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _1370_
timestamp 1
transform -1 0 25760 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1371_
timestamp 1
transform -1 0 25300 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1372_
timestamp 1
transform 1 0 23644 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__or4b_1  _1373_
timestamp 1
transform -1 0 25116 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1374_
timestamp 1
transform -1 0 25484 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1375_
timestamp 1
transform 1 0 25484 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1376_
timestamp 1
transform -1 0 25668 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_1  _1377_
timestamp 1
transform 1 0 25024 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1378_
timestamp 1
transform -1 0 25024 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1379_
timestamp 1
transform 1 0 24380 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1380_
timestamp 1
transform -1 0 25208 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1381_
timestamp 1
transform 1 0 23828 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1382_
timestamp 1
transform -1 0 24288 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1383_
timestamp 1
transform -1 0 24380 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _1384_
timestamp 1
transform 1 0 24380 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1385_
timestamp 1
transform -1 0 23184 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _1386_
timestamp 1
transform -1 0 23460 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1387_
timestamp 1
transform 1 0 22540 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1388_
timestamp 1
transform -1 0 22540 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1389_
timestamp 1
transform -1 0 26496 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1390_
timestamp 1
transform -1 0 26220 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1391_
timestamp 1
transform -1 0 21896 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1392_
timestamp 1
transform -1 0 23460 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1393_
timestamp 1
transform -1 0 20884 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1394_
timestamp 1
transform -1 0 20240 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_2  _1395_
timestamp 1
transform 1 0 22540 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1396_
timestamp 1
transform 1 0 23276 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1397_
timestamp 1
transform -1 0 23552 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1398_
timestamp 1
transform 1 0 22632 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1399_
timestamp 1
transform 1 0 22540 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1400_
timestamp 1
transform -1 0 22632 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1401_
timestamp 1
transform -1 0 22448 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _1402_
timestamp 1
transform -1 0 23644 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1403_
timestamp 1
transform 1 0 20700 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1404_
timestamp 1
transform -1 0 21436 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1405_
timestamp 1
transform 1 0 20424 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a2111o_1  _1406_
timestamp 1
transform -1 0 21252 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _1407_
timestamp 1
transform -1 0 25300 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1408_
timestamp 1
transform 1 0 21252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1409_
timestamp 1
transform -1 0 20424 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1410_
timestamp 1
transform 1 0 19596 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1411_
timestamp 1
transform -1 0 21712 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1412_
timestamp 1
transform 1 0 20976 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1413_
timestamp 1
transform -1 0 19412 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1414_
timestamp 1
transform 1 0 21528 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1415_
timestamp 1
transform 1 0 20700 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_2  _1416_
timestamp 1
transform -1 0 24656 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1417_
timestamp 1
transform 1 0 25668 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1418_
timestamp 1
transform 1 0 25576 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1419_
timestamp 1
transform -1 0 20424 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_1  _1420_
timestamp 1
transform 1 0 19044 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a31oi_1  _1421_
timestamp 1
transform 1 0 20332 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1422_
timestamp 1
transform 1 0 20056 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _1423_
timestamp 1
transform 1 0 18492 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1424_
timestamp 1
transform 1 0 13432 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1425_
timestamp 1
transform -1 0 12880 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1426_
timestamp 1
transform -1 0 11040 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1427_
timestamp 1
transform 1 0 19228 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1428_
timestamp 1
transform 1 0 14536 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1429_
timestamp 1
transform -1 0 15364 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1430_
timestamp 1
transform 1 0 18492 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1431_
timestamp 1
transform 1 0 17940 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1432_
timestamp 1
transform -1 0 18768 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1433_
timestamp 1
transform 1 0 18308 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1434_
timestamp 1
transform -1 0 21712 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1435_
timestamp 1
transform -1 0 22448 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1436_
timestamp 1
transform 1 0 20700 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1437_
timestamp 1
transform 1 0 20792 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1438_
timestamp 1
transform -1 0 19596 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1439_
timestamp 1
transform 1 0 21804 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _1440_
timestamp 1
transform 1 0 16928 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1441_
timestamp 1
transform 1 0 17388 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1442_
timestamp 1
transform 1 0 14812 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1443_
timestamp 1
transform -1 0 16192 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1444_
timestamp 1
transform 1 0 17388 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1445_
timestamp 1
transform 1 0 16652 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1446_
timestamp 1
transform 1 0 16744 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1447_
timestamp 1
transform -1 0 20608 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1448_
timestamp 1
transform -1 0 15824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1449_
timestamp 1
transform -1 0 16376 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a311o_1  _1450_
timestamp 1
transform 1 0 19964 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o31ai_1  _1451_
timestamp 1
transform 1 0 15364 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1452_
timestamp 1
transform 1 0 15824 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1453_
timestamp 1
transform 1 0 19872 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1454_
timestamp 1
transform -1 0 19872 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1455_
timestamp 1
transform -1 0 18768 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1456_
timestamp 1
transform -1 0 15732 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1457_
timestamp 1
transform -1 0 15916 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1458_
timestamp 1
transform 1 0 15916 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _1459_
timestamp 1
transform 1 0 16652 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1460_
timestamp 1
transform -1 0 20516 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1461_
timestamp 1
transform 1 0 19872 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _1462_
timestamp 1
transform -1 0 20148 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1463_
timestamp 1
transform -1 0 15456 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1464_
timestamp 1
transform -1 0 15456 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1465_
timestamp 1
transform -1 0 15180 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _1466_
timestamp 1
transform 1 0 13800 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1467_
timestamp 1
transform 1 0 18676 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1468_
timestamp 1
transform 1 0 18860 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1469_
timestamp 1
transform 1 0 14628 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1470_
timestamp 1
transform 1 0 15824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1471_
timestamp 1
transform -1 0 15824 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _1472_
timestamp 1
transform 1 0 14720 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1473_
timestamp 1
transform -1 0 18492 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1474_
timestamp 1
transform 1 0 18400 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1475_
timestamp 1
transform 1 0 17756 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1476_
timestamp 1
transform -1 0 17112 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1477_
timestamp 1
transform -1 0 16560 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1478_
timestamp 1
transform 1 0 17848 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _1479_
timestamp 1
transform 1 0 16744 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__nand2b_1  _1480_
timestamp 1
transform -1 0 20976 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _1481_
timestamp 1
transform -1 0 20516 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1482_
timestamp 1
transform 1 0 19780 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1483_
timestamp 1
transform -1 0 19136 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1484_
timestamp 1
transform -1 0 16928 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1485_
timestamp 1
transform -1 0 15456 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1486_
timestamp 1
transform 1 0 16836 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _1487_
timestamp 1
transform 1 0 17204 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _1488_
timestamp 1
transform -1 0 21712 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1489_
timestamp 1
transform -1 0 19872 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1490_
timestamp 1
transform 1 0 17112 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1491_
timestamp 1
transform 1 0 18032 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1492_
timestamp 1
transform 1 0 17296 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1493_
timestamp 1
transform -1 0 20976 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a311o_1  _1494_
timestamp 1
transform -1 0 22540 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1495_
timestamp 1
transform -1 0 15364 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1496_
timestamp 1
transform 1 0 15916 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1497_
timestamp 1
transform -1 0 15272 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1498_
timestamp 1
transform 1 0 15916 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _1499_
timestamp 1
transform 1 0 14720 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1500_
timestamp 1
transform 1 0 18400 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1501_
timestamp 1
transform 1 0 17572 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1502_
timestamp 1
transform 1 0 16100 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1503_
timestamp 1
transform 1 0 16192 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _1504_
timestamp 1
transform 1 0 16652 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1505_
timestamp 1
transform -1 0 15916 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1506_
timestamp 1
transform -1 0 18400 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_2  _1507_
timestamp 1
transform 1 0 19228 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1508_
timestamp 1
transform -1 0 16744 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1509_
timestamp 1
transform -1 0 15272 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1510_
timestamp 1
transform -1 0 15548 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1511_
timestamp 1
transform 1 0 14536 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1512_
timestamp 1
transform -1 0 13800 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1513_
timestamp 1
transform -1 0 17940 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1514_
timestamp 1
transform -1 0 18308 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _1515_
timestamp 1
transform -1 0 17572 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1516_
timestamp 1
transform -1 0 14812 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1517_
timestamp 1
transform 1 0 13800 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1518_
timestamp 1
transform -1 0 14444 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _1519_
timestamp 1
transform 1 0 13616 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_1  _1520_
timestamp 1
transform 1 0 19504 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1521_
timestamp 1
transform -1 0 18676 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1522_
timestamp 1
transform -1 0 18400 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1523_
timestamp 1
transform 1 0 12604 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1524_
timestamp 1
transform 1 0 13984 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1525_
timestamp 1
transform -1 0 13984 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1526_
timestamp 1
transform 1 0 17848 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1527_
timestamp 1
transform -1 0 13248 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1528_
timestamp 1
transform 1 0 12144 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1529_
timestamp 1
transform 1 0 13064 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1530_
timestamp 1
transform 1 0 13064 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1531_
timestamp 1
transform 1 0 10764 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1532_
timestamp 1
transform -1 0 9476 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1533_
timestamp 1
transform -1 0 9844 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1534_
timestamp 1
transform 1 0 9844 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1535_
timestamp 1
transform -1 0 8188 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1536_
timestamp 1
transform -1 0 5980 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1537_
timestamp 1
transform -1 0 6256 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1538_
timestamp 1
transform 1 0 4784 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1539_
timestamp 1
transform 1 0 6808 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1540_
timestamp 1
transform -1 0 6808 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1541_
timestamp 1
transform 1 0 6624 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1542_
timestamp 1
transform 1 0 7360 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1543_
timestamp 1
transform -1 0 4140 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1544_
timestamp 1
transform -1 0 4416 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1545_
timestamp 1
transform 1 0 2760 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1546_
timestamp 1
transform 1 0 3588 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1547_
timestamp 1
transform -1 0 3404 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1548_
timestamp 1
transform -1 0 2944 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1549_
timestamp 1
transform 1 0 1932 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1550_
timestamp 1
transform -1 0 2944 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1551_
timestamp 1
transform 1 0 2944 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1552_
timestamp 1
transform 1 0 1748 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1553_
timestamp 1
transform -1 0 1748 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1554_
timestamp 1
transform -1 0 2300 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1555_
timestamp 1
transform 1 0 2024 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1556_
timestamp 1
transform 1 0 1748 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1557_
timestamp 1
transform 1 0 1380 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1558_
timestamp 1
transform 1 0 1932 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1559_
timestamp 1
transform -1 0 11040 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_2  _1560_
timestamp 1
transform 1 0 6072 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1561_
timestamp 1
transform -1 0 9660 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1562_
timestamp 1
transform -1 0 9568 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1563_
timestamp 1
transform 1 0 7820 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1564_
timestamp 1
transform 1 0 7820 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _1565_
timestamp 1
transform -1 0 8464 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1566_
timestamp 1
transform 1 0 8188 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1567_
timestamp 1
transform -1 0 8372 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1568_
timestamp 1
transform -1 0 8004 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a2111oi_1  _1569_
timestamp 1
transform 1 0 7084 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _1570_
timestamp 1
transform -1 0 7636 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1571_
timestamp 1
transform -1 0 3220 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1572_
timestamp 1
transform -1 0 4140 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1573_
timestamp 1
transform -1 0 2760 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1574_
timestamp 1
transform -1 0 3128 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1575_
timestamp 1
transform -1 0 3220 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1576_
timestamp 1
transform -1 0 2116 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1577_
timestamp 1
transform -1 0 2484 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1578_
timestamp 1
transform -1 0 2024 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1579_
timestamp 1
transform 1 0 1656 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1580_
timestamp 1
transform 1 0 2576 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1581_
timestamp 1
transform 1 0 2944 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _1582_
timestamp 1
transform 1 0 18584 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1583_
timestamp 1
transform 1 0 19688 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1584_
timestamp 1
transform 1 0 19688 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1585_
timestamp 1
transform 1 0 18584 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1586_
timestamp 1
transform 1 0 16652 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1587_
timestamp 1
transform -1 0 19596 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1588_
timestamp 1
transform -1 0 18768 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1589_
timestamp 1
transform -1 0 18584 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1590_
timestamp 1
transform 1 0 15088 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1591_
timestamp 1
transform 1 0 14076 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1592_
timestamp 1
transform 1 0 14076 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1593_
timestamp 1
transform 1 0 14444 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1594_
timestamp 1
transform 1 0 12604 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1595_
timestamp 1
transform 1 0 11684 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1596_
timestamp 1
transform 1 0 10764 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1597_
timestamp 1
transform 1 0 11224 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1598_
timestamp 1
transform 1 0 7360 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1599_
timestamp 1
transform 1 0 7728 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1600_
timestamp 1
transform 1 0 7452 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1601_
timestamp 1
transform -1 0 8188 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1602_
timestamp 1
transform 1 0 1380 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1603_
timestamp 1
transform 1 0 3772 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1604_
timestamp 1
transform 1 0 2208 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1605_
timestamp 1
transform 1 0 1380 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1606_
timestamp 1
transform 1 0 3772 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1607_
timestamp 1
transform 1 0 2208 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1608_
timestamp 1
transform 1 0 1380 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1609_
timestamp 1
transform 1 0 3772 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1610_
timestamp 1
transform 1 0 2300 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1611_
timestamp 1
transform 1 0 6624 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1612_
timestamp 1
transform 1 0 4784 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1613_
timestamp 1
transform 1 0 9384 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1614_
timestamp 1
transform 1 0 9384 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1615_
timestamp 1
transform 1 0 10120 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1616_
timestamp 1
transform -1 0 12420 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1617_
timestamp 1
transform 1 0 12512 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1618_
timestamp 1
transform 1 0 12420 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1619_
timestamp 1
transform -1 0 15824 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1620_
timestamp 1
transform 1 0 11500 0 -1 20672
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1621_
timestamp 1
transform 1 0 19228 0 1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1622_
timestamp 1
transform 1 0 19228 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1623_
timestamp 1
transform 1 0 17388 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1624_
timestamp 1
transform 1 0 16652 0 -1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1625_
timestamp 1
transform 1 0 16284 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1626_
timestamp 1
transform 1 0 12512 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1627_
timestamp 1
transform 1 0 14076 0 1 17408
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1628_
timestamp 1
transform 1 0 16652 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1629_
timestamp 1
transform 1 0 15732 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1630_
timestamp 1
transform 1 0 17940 0 -1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1631_
timestamp 1
transform 1 0 14444 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1632_
timestamp 1
transform 1 0 15456 0 1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1633_
timestamp 1
transform 1 0 13248 0 -1 11968
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1634_
timestamp 1
transform -1 0 13616 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1635_
timestamp 1
transform -1 0 13984 0 -1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1636_
timestamp 1
transform 1 0 11500 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1637_
timestamp 1
transform 1 0 8188 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1638_
timestamp 1
transform 1 0 3864 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1639_
timestamp 1
transform 1 0 7176 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1640_
timestamp 1
transform 1 0 2208 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1641_
timestamp 1
transform 1 0 1380 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1642_
timestamp 1
transform 1 0 1380 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1643_
timestamp 1
transform 1 0 2392 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1644_
timestamp 1
transform 1 0 1932 0 1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1645_
timestamp 1
transform -1 0 10764 0 -1 28288
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1646_
timestamp 1
transform -1 0 10764 0 1 26112
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1647_
timestamp 1
transform -1 0 10120 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1648_
timestamp 1
transform 1 0 7360 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1649_
timestamp 1
transform -1 0 6256 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1650_
timestamp 1
transform -1 0 4784 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1651_
timestamp 1
transform 1 0 1380 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1652_
timestamp 1
transform 1 0 1380 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1653_
timestamp 1
transform 1 0 2484 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_CLK_10MHZ
timestamp 1
transform 1 0 10580 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_CLK_10MHZ
timestamp 1
transform 1 0 5428 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_CLK_10MHZ
timestamp 1
transform -1 0 6072 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_CLK_10MHZ
timestamp 1
transform -1 0 7084 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_CLK_10MHZ
timestamp 1
transform 1 0 8924 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_CLK_10MHZ
timestamp 1
transform -1 0 14168 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_CLK_10MHZ
timestamp 1
transform 1 0 14720 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_CLK_10MHZ
timestamp 1
transform -1 0 14720 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_CLK_10MHZ
timestamp 1
transform 1 0 15364 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_6  clkload0
timestamp 1
transform 1 0 5520 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__clkinvlp_4  clkload1
timestamp 1
transform 1 0 4600 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__bufinv_16  clkload2
timestamp 1
transform 1 0 5244 0 1 22848
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinv_2  clkload3
timestamp 1
transform 1 0 8464 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_4  clkload4
timestamp 1
transform 1 0 12328 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__bufinv_16  clkload5
timestamp 1
transform 1 0 15088 0 1 18496
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinv_2  clkload6
timestamp 1
transform 1 0 12512 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout14
timestamp 1
transform 1 0 21712 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout15
timestamp 1
transform -1 0 20424 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout16
timestamp 1
transform -1 0 25944 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout17
timestamp 1
transform -1 0 26220 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout18
timestamp 1
transform 1 0 24380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout19
timestamp 1
transform 1 0 25484 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout20
timestamp 1
transform -1 0 25300 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout22
timestamp 1
transform 1 0 22172 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout23
timestamp 1
transform 1 0 21804 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout24
timestamp 1
transform 1 0 15824 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout25
timestamp 1
transform 1 0 14812 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout26
timestamp 1
transform 1 0 14628 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout27
timestamp 1
transform -1 0 6072 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout28
timestamp 1
transform 1 0 4692 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout30
timestamp 1
transform -1 0 9292 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout31
timestamp 1
transform 1 0 14076 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout32
timestamp 1
transform -1 0 12512 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout33
timestamp 1
transform 1 0 12512 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout34
timestamp 1
transform -1 0 14628 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout35
timestamp 1
transform 1 0 15824 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout36
timestamp 1
transform -1 0 9292 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout37
timestamp 1
transform -1 0 5244 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout39
timestamp 1
transform -1 0 9292 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout40
timestamp 1
transform 1 0 14076 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout41
timestamp 1
transform 1 0 12696 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout42
timestamp 1
transform 1 0 8096 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout43
timestamp 1
transform 1 0 3312 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout44
timestamp 1
transform 1 0 3220 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout45
timestamp 1
transform 1 0 8740 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout46
timestamp 1
transform -1 0 17296 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout47
timestamp 1
transform -1 0 17848 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout48
timestamp 1
transform 1 0 14444 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout49
timestamp 1
transform -1 0 16192 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout50
timestamp 1
transform -1 0 18308 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout51
timestamp 1
transform 1 0 21344 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3
timestamp 1636968456
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1636968456
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp 1
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1636968456
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1636968456
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp 1
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1636968456
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1636968456
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1636968456
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_97
timestamp 1
transform 1 0 10028 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_102
timestamp 1
transform 1 0 10488 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113
timestamp 1
transform 1 0 11500 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_120
timestamp 1636968456
transform 1 0 12144 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_132
timestamp 1
transform 1 0 13248 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_141
timestamp 1
transform 1 0 14076 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_149
timestamp 1
transform 1 0 14812 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_161
timestamp 1
transform 1 0 15916 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_169
timestamp 1
transform 1 0 16652 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_177
timestamp 1
transform 1 0 17388 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_183
timestamp 1636968456
transform 1 0 17940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1636968456
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1636968456
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1636968456
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1636968456
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1636968456
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1636968456
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_281
timestamp 1
transform 1 0 26956 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_287
timestamp 1
transform 1 0 27508 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_6
timestamp 1636968456
transform 1 0 1656 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_18
timestamp 1636968456
transform 1 0 2760 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_30
timestamp 1636968456
transform 1 0 3864 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_42
timestamp 1636968456
transform 1 0 4968 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1636968456
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1636968456
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_81
timestamp 1
transform 1 0 8556 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_89
timestamp 1
transform 1 0 9292 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_113
timestamp 1
transform 1 0 11500 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_126
timestamp 1
transform 1 0 12696 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_169
timestamp 1
transform 1 0 16652 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_189
timestamp 1
transform 1 0 18492 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_215
timestamp 1
transform 1 0 20884 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_234
timestamp 1636968456
transform 1 0 22632 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_246
timestamp 1636968456
transform 1 0 23736 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_258
timestamp 1636968456
transform 1 0 24840 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_270
timestamp 1
transform 1 0 25944 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_278
timestamp 1
transform 1 0 26680 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_281
timestamp 1
transform 1 0 26956 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1636968456
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1636968456
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1636968456
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1636968456
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1636968456
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1636968456
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_98
timestamp 1636968456
transform 1 0 10120 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_118
timestamp 1636968456
transform 1 0 11960 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_130
timestamp 1
transform 1 0 13064 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_134
timestamp 1
transform 1 0 13432 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_163
timestamp 1
transform 1 0 16100 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_190
timestamp 1
transform 1 0 18584 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_197
timestamp 1
transform 1 0 19228 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_220
timestamp 1
transform 1 0 21344 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_248
timestamp 1
transform 1 0 23920 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_253
timestamp 1
transform 1 0 24380 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_263
timestamp 1636968456
transform 1 0 25300 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_275
timestamp 1636968456
transform 1 0 26404 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_287
timestamp 1
transform 1 0 27508 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1636968456
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1636968456
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1636968456
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1636968456
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1636968456
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1636968456
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1636968456
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_93
timestamp 1
transform 1 0 9660 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_121
timestamp 1636968456
transform 1 0 12236 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_133
timestamp 1636968456
transform 1 0 13340 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_145
timestamp 1
transform 1 0 14444 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_169
timestamp 1
transform 1 0 16652 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_177
timestamp 1636968456
transform 1 0 17388 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_189
timestamp 1636968456
transform 1 0 18492 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_201
timestamp 1
transform 1 0 19596 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_244
timestamp 1
transform 1 0 23552 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_250
timestamp 1
transform 1 0 24104 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_269
timestamp 1
transform 1 0 25852 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_277
timestamp 1
transform 1 0 26588 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_281
timestamp 1
transform 1 0 26956 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_287
timestamp 1
transform 1 0 27508 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1636968456
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1636968456
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_29
timestamp 1
transform 1 0 3772 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_37
timestamp 1
transform 1 0 4508 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_50
timestamp 1
transform 1 0 5704 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_60
timestamp 1
transform 1 0 6624 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_4_92
timestamp 1
transform 1 0 9568 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_100
timestamp 1
transform 1 0 10304 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_105
timestamp 1636968456
transform 1 0 10764 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_117
timestamp 1
transform 1 0 11868 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_121
timestamp 1
transform 1 0 12236 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_134
timestamp 1
transform 1 0 13432 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_4_148
timestamp 1
transform 1 0 14720 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_161
timestamp 1
transform 1 0 15916 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_168
timestamp 1636968456
transform 1 0 16560 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_180
timestamp 1
transform 1 0 17664 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_190
timestamp 1
transform 1 0 18584 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_4_197
timestamp 1
transform 1 0 19228 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_205
timestamp 1
transform 1 0 19964 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_212
timestamp 1636968456
transform 1 0 20608 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_224
timestamp 1
transform 1 0 21712 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1636968456
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_264
timestamp 1636968456
transform 1 0 25392 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_276
timestamp 1636968456
transform 1 0 26496 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1636968456
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1636968456
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_27
timestamp 1
transform 1 0 3588 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_35
timestamp 1
transform 1 0 4324 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_48
timestamp 1
transform 1 0 5520 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_64
timestamp 1
transform 1 0 6992 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_72
timestamp 1
transform 1 0 7728 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_97
timestamp 1636968456
transform 1 0 10028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_109
timestamp 1
transform 1 0 11132 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_122
timestamp 1636968456
transform 1 0 12328 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_134
timestamp 1
transform 1 0 13432 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_141
timestamp 1
transform 1 0 14076 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_162
timestamp 1
transform 1 0 16008 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_196
timestamp 1
transform 1 0 19136 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_202
timestamp 1
transform 1 0 19688 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_206
timestamp 1636968456
transform 1 0 20056 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_218
timestamp 1
transform 1 0 21160 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_225
timestamp 1
transform 1 0 21804 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_238
timestamp 1
transform 1 0 23000 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_246
timestamp 1
transform 1 0 23736 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_254
timestamp 1
transform 1 0 24472 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_264
timestamp 1636968456
transform 1 0 25392 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_276
timestamp 1
transform 1 0 26496 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_281
timestamp 1
transform 1 0 26956 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_287
timestamp 1
transform 1 0 27508 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1636968456
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1636968456
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1636968456
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_41
timestamp 1
transform 1 0 4876 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_49
timestamp 1
transform 1 0 5612 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_55
timestamp 1
transform 1 0 6164 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_63
timestamp 1
transform 1 0 6900 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_73
timestamp 1
transform 1 0 7820 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_81
timestamp 1
transform 1 0 8556 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_85
timestamp 1
transform 1 0 8924 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_89
timestamp 1
transform 1 0 9292 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_97
timestamp 1
transform 1 0 10028 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_6_111
timestamp 1
transform 1 0 11316 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_128
timestamp 1
transform 1 0 12880 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_135
timestamp 1
transform 1 0 13524 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_141
timestamp 1
transform 1 0 14076 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_150
timestamp 1636968456
transform 1 0 14904 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_162
timestamp 1
transform 1 0 16008 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_168
timestamp 1
transform 1 0 16560 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_189
timestamp 1
transform 1 0 18492 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_197
timestamp 1
transform 1 0 19228 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_232
timestamp 1636968456
transform 1 0 22448 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_253
timestamp 1
transform 1 0 24380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_257
timestamp 1
transform 1 0 24748 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_266
timestamp 1636968456
transform 1 0 25576 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_278
timestamp 1
transform 1 0 26680 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_286
timestamp 1
transform 1 0 27416 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1636968456
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1636968456
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1636968456
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_39
timestamp 1
transform 1 0 4692 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_52
timestamp 1
transform 1 0 5888 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_64
timestamp 1
transform 1 0 6992 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_79
timestamp 1636968456
transform 1 0 8372 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_91
timestamp 1
transform 1 0 9476 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_97
timestamp 1
transform 1 0 10028 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_113
timestamp 1
transform 1 0 11500 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_164
timestamp 1
transform 1 0 16192 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1636968456
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_181
timestamp 1
transform 1 0 17756 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_195
timestamp 1636968456
transform 1 0 19044 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_207
timestamp 1
transform 1 0 20148 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_211
timestamp 1
transform 1 0 20516 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_221
timestamp 1
transform 1 0 21436 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1636968456
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_237
timestamp 1
transform 1 0 22908 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1636968456
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_261
timestamp 1
transform 1 0 25116 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_266
timestamp 1636968456
transform 1 0 25576 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_278
timestamp 1
transform 1 0 26680 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_281
timestamp 1
transform 1 0 26956 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_287
timestamp 1
transform 1 0 27508 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1636968456
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1636968456
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1636968456
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1636968456
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_59
timestamp 1636968456
transform 1 0 6532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_71
timestamp 1636968456
transform 1 0 7636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1636968456
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1636968456
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1636968456
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_153
timestamp 1
transform 1 0 15180 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_169
timestamp 1
transform 1 0 16652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_180
timestamp 1636968456
transform 1 0 17664 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_192
timestamp 1
transform 1 0 18768 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_200
timestamp 1
transform 1 0 19504 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_210
timestamp 1
transform 1 0 20424 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_218
timestamp 1
transform 1 0 21160 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_232
timestamp 1
transform 1 0 22448 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_240
timestamp 1
transform 1 0 23184 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_249
timestamp 1
transform 1 0 24012 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_253
timestamp 1
transform 1 0 24380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_257
timestamp 1
transform 1 0 24748 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_275
timestamp 1636968456
transform 1 0 26404 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_287
timestamp 1
transform 1 0 27508 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1636968456
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1636968456
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_27
timestamp 1
transform 1 0 3588 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_35
timestamp 1
transform 1 0 4324 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_43
timestamp 1
transform 1 0 5060 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_47
timestamp 1
transform 1 0 5428 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_63
timestamp 1
transform 1 0 6900 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_75
timestamp 1
transform 1 0 8004 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_85
timestamp 1
transform 1 0 8924 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_93
timestamp 1
transform 1 0 9660 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_99
timestamp 1
transform 1 0 10212 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_103
timestamp 1
transform 1 0 10580 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_129
timestamp 1
transform 1 0 12972 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_137
timestamp 1
transform 1 0 13708 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_9_150
timestamp 1
transform 1 0 14904 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_165
timestamp 1
transform 1 0 16284 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_169
timestamp 1
transform 1 0 16652 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_225
timestamp 1
transform 1 0 21804 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_233
timestamp 1
transform 1 0 22540 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_243
timestamp 1
transform 1 0 23460 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_255
timestamp 1
transform 1 0 24564 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_270
timestamp 1
transform 1 0 25944 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_278
timestamp 1
transform 1 0 26680 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_281
timestamp 1
transform 1 0 26956 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_287
timestamp 1
transform 1 0 27508 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1636968456
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1636968456
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_29
timestamp 1
transform 1 0 3772 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_54
timestamp 1636968456
transform 1 0 6072 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_66
timestamp 1
transform 1 0 7176 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_88
timestamp 1
transform 1 0 9200 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_99
timestamp 1
transform 1 0 10212 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_120
timestamp 1
transform 1 0 12144 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_141
timestamp 1
transform 1 0 14076 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_155
timestamp 1636968456
transform 1 0 15364 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_167
timestamp 1636968456
transform 1 0 16468 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_185
timestamp 1
transform 1 0 18124 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_193
timestamp 1
transform 1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_208
timestamp 1636968456
transform 1 0 20240 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_220
timestamp 1
transform 1 0 21344 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_10_236
timestamp 1
transform 1 0 22816 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1636968456
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1636968456
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_277
timestamp 1
transform 1 0 26588 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_285
timestamp 1
transform 1 0 27324 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1636968456
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_15
timestamp 1
transform 1 0 2484 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_23
timestamp 1
transform 1 0 3220 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_31
timestamp 1
transform 1 0 3956 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_37
timestamp 1
transform 1 0 4508 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_42
timestamp 1636968456
transform 1 0 4968 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_63
timestamp 1636968456
transform 1 0 6900 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_75
timestamp 1636968456
transform 1 0 8004 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_87
timestamp 1
transform 1 0 9108 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_103
timestamp 1
transform 1 0 10580 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_107
timestamp 1
transform 1 0 10948 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_113
timestamp 1
transform 1 0 11500 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_117
timestamp 1
transform 1 0 11868 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_143
timestamp 1
transform 1 0 14260 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_11_162
timestamp 1
transform 1 0 16008 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_176
timestamp 1
transform 1 0 17296 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_263
timestamp 1636968456
transform 1 0 25300 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_275
timestamp 1
transform 1 0 26404 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_281
timestamp 1
transform 1 0 26956 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_287
timestamp 1
transform 1 0 27508 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1636968456
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1636968456
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_34
timestamp 1
transform 1 0 4232 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_42
timestamp 1
transform 1 0 4968 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_53
timestamp 1
transform 1 0 5980 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_70
timestamp 1
transform 1 0 7544 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_85
timestamp 1
transform 1 0 8924 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_93
timestamp 1
transform 1 0 9660 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_107
timestamp 1
transform 1 0 10948 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_112
timestamp 1
transform 1 0 11408 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_120
timestamp 1
transform 1 0 12144 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_128
timestamp 1
transform 1 0 12880 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_132
timestamp 1
transform 1 0 13248 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_141
timestamp 1
transform 1 0 14076 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_155
timestamp 1
transform 1 0 15364 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_161
timestamp 1
transform 1 0 15916 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_186
timestamp 1
transform 1 0 18216 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_197
timestamp 1
transform 1 0 19228 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_218
timestamp 1
transform 1 0 21160 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_237
timestamp 1636968456
transform 1 0 22908 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_270
timestamp 1636968456
transform 1 0 25944 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_282
timestamp 1
transform 1 0 27048 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1636968456
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_15
timestamp 1
transform 1 0 2484 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_23
timestamp 1
transform 1 0 3220 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_50
timestamp 1
transform 1 0 5704 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_13_63
timestamp 1
transform 1 0 6900 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_92
timestamp 1636968456
transform 1 0 9568 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_104
timestamp 1
transform 1 0 10672 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_120
timestamp 1
transform 1 0 12144 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_163
timestamp 1
transform 1 0 16100 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_178
timestamp 1636968456
transform 1 0 17480 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_190
timestamp 1
transform 1 0 18584 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_198
timestamp 1
transform 1 0 19320 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_206
timestamp 1636968456
transform 1 0 20056 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_218
timestamp 1
transform 1 0 21160 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1636968456
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_237
timestamp 1
transform 1 0 22908 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_250
timestamp 1636968456
transform 1 0 24104 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_262
timestamp 1636968456
transform 1 0 25208 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_274
timestamp 1
transform 1 0 26312 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_13_281
timestamp 1
transform 1 0 26956 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_287
timestamp 1
transform 1 0 27508 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1636968456
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1636968456
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1636968456
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_41
timestamp 1
transform 1 0 4876 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_53
timestamp 1
transform 1 0 5980 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_63
timestamp 1
transform 1 0 6900 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_71
timestamp 1
transform 1 0 7636 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_78
timestamp 1
transform 1 0 8280 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_98
timestamp 1
transform 1 0 10120 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_122
timestamp 1636968456
transform 1 0 12328 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_134
timestamp 1
transform 1 0 13432 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_167
timestamp 1
transform 1 0 16468 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_182
timestamp 1
transform 1 0 17848 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_190
timestamp 1
transform 1 0 18584 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_197
timestamp 1
transform 1 0 19228 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_211
timestamp 1
transform 1 0 20516 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_14_234
timestamp 1
transform 1 0 22632 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_240
timestamp 1
transform 1 0 23184 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1636968456
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_279
timestamp 1
transform 1 0 26772 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_287
timestamp 1
transform 1 0 27508 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1636968456
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_15
timestamp 1
transform 1 0 2484 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_44
timestamp 1636968456
transform 1 0 5152 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_74
timestamp 1636968456
transform 1 0 7912 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_86
timestamp 1
transform 1 0 9016 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_94
timestamp 1636968456
transform 1 0 9752 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_106
timestamp 1
transform 1 0 10856 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_15_113
timestamp 1
transform 1 0 11500 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_119
timestamp 1
transform 1 0 12052 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_131
timestamp 1636968456
transform 1 0 13156 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_143
timestamp 1636968456
transform 1 0 14260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_155
timestamp 1
transform 1 0 15364 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_186
timestamp 1636968456
transform 1 0 18216 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_198
timestamp 1
transform 1 0 19320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_204
timestamp 1
transform 1 0 19872 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_219
timestamp 1
transform 1 0 21252 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_239
timestamp 1636968456
transform 1 0 23092 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_251
timestamp 1
transform 1 0 24196 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_268
timestamp 1636968456
transform 1 0 25760 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_281
timestamp 1
transform 1 0 26956 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_287
timestamp 1
transform 1 0 27508 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1636968456
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1636968456
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_29
timestamp 1
transform 1 0 3772 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_37
timestamp 1
transform 1 0 4508 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_42
timestamp 1
transform 1 0 4968 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_51
timestamp 1636968456
transform 1 0 5796 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_63
timestamp 1
transform 1 0 6900 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_67
timestamp 1
transform 1 0 7268 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_80
timestamp 1
transform 1 0 8464 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_90
timestamp 1
transform 1 0 9384 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_112
timestamp 1636968456
transform 1 0 11408 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_163
timestamp 1636968456
transform 1 0 16100 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_182
timestamp 1
transform 1 0 17848 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_202
timestamp 1636968456
transform 1 0 19688 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_214
timestamp 1636968456
transform 1 0 20792 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_226
timestamp 1
transform 1 0 21896 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_232
timestamp 1636968456
transform 1 0 22448 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_244
timestamp 1
transform 1 0 23552 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_253
timestamp 1
transform 1 0 24380 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_257
timestamp 1636968456
transform 1 0 24748 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_269
timestamp 1
transform 1 0 25852 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_274
timestamp 1636968456
transform 1 0 26312 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_286
timestamp 1
transform 1 0 27416 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_19
timestamp 1
transform 1 0 2852 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_27
timestamp 1
transform 1 0 3588 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_31
timestamp 1
transform 1 0 3956 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_17_78
timestamp 1
transform 1 0 8280 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_84
timestamp 1
transform 1 0 8832 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_88
timestamp 1
transform 1 0 9200 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_96
timestamp 1
transform 1 0 9936 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_113
timestamp 1
transform 1 0 11500 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_126
timestamp 1
transform 1 0 12696 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1636968456
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1636968456
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_181
timestamp 1
transform 1 0 17756 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_189
timestamp 1
transform 1 0 18492 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_195
timestamp 1636968456
transform 1 0 19044 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_207
timestamp 1
transform 1 0 20148 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_211
timestamp 1
transform 1 0 20516 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_219
timestamp 1
transform 1 0 21252 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1636968456
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_237
timestamp 1
transform 1 0 22908 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_258
timestamp 1
transform 1 0 24840 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_17_277
timestamp 1
transform 1 0 26588 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_286
timestamp 1
transform 1 0 27416 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_3
timestamp 1
transform 1 0 1380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_23
timestamp 1
transform 1 0 3220 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_58
timestamp 1
transform 1 0 6440 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_85
timestamp 1
transform 1 0 8924 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1636968456
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_109
timestamp 1
transform 1 0 11132 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_113
timestamp 1
transform 1 0 11500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_117
timestamp 1
transform 1 0 11868 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_126
timestamp 1636968456
transform 1 0 12696 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1636968456
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_153
timestamp 1
transform 1 0 15180 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_173
timestamp 1
transform 1 0 17020 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_183
timestamp 1636968456
transform 1 0 17940 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_197
timestamp 1
transform 1 0 19228 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_215
timestamp 1
transform 1 0 20884 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_221
timestamp 1
transform 1 0 21436 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_243
timestamp 1
transform 1 0 23460 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_253
timestamp 1
transform 1 0 24380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_259
timestamp 1
transform 1 0 24932 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_270
timestamp 1636968456
transform 1 0 25944 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_282
timestamp 1
transform 1 0 27048 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1636968456
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_15
timestamp 1
transform 1 0 2484 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_23
timestamp 1
transform 1 0 3220 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_33
timestamp 1636968456
transform 1 0 4140 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_45
timestamp 1
transform 1 0 5244 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_53
timestamp 1
transform 1 0 5980 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_70
timestamp 1
transform 1 0 7544 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_80
timestamp 1636968456
transform 1 0 8464 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_92
timestamp 1
transform 1 0 9568 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1636968456
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_125
timestamp 1
transform 1 0 12604 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_19_138
timestamp 1
transform 1 0 13800 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_161
timestamp 1
transform 1 0 15916 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_177
timestamp 1
transform 1 0 17388 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_199
timestamp 1
transform 1 0 19412 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_207
timestamp 1
transform 1 0 20148 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_214
timestamp 1
transform 1 0 20792 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1636968456
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_237
timestamp 1
transform 1 0 22908 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_278
timestamp 1
transform 1 0 26680 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_281
timestamp 1
transform 1 0 26956 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_287
timestamp 1
transform 1 0 27508 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_3
timestamp 1
transform 1 0 1380 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_7
timestamp 1
transform 1 0 1748 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_13
timestamp 1636968456
transform 1 0 2300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_25
timestamp 1
transform 1 0 3404 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_34
timestamp 1
transform 1 0 4232 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_42
timestamp 1
transform 1 0 4968 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_49
timestamp 1636968456
transform 1 0 5612 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_61
timestamp 1
transform 1 0 6716 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_88
timestamp 1
transform 1 0 9200 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_96
timestamp 1
transform 1 0 9936 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_101
timestamp 1
transform 1 0 10396 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_105
timestamp 1
transform 1 0 10764 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_117
timestamp 1636968456
transform 1 0 11868 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_129
timestamp 1
transform 1 0 12972 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_137
timestamp 1
transform 1 0 13708 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_145
timestamp 1
transform 1 0 14444 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_157
timestamp 1
transform 1 0 15548 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_168
timestamp 1636968456
transform 1 0 16560 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_180
timestamp 1636968456
transform 1 0 17664 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_192
timestamp 1
transform 1 0 18768 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_204
timestamp 1
transform 1 0 19872 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_227
timestamp 1
transform 1 0 21988 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_240
timestamp 1636968456
transform 1 0 23184 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_261
timestamp 1
transform 1 0 25116 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_274
timestamp 1636968456
transform 1 0 26312 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_286
timestamp 1
transform 1 0 27416 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_30
timestamp 1
transform 1 0 3864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_65
timestamp 1
transform 1 0 7084 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_21_80
timestamp 1
transform 1 0 8464 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_88
timestamp 1
transform 1 0 9200 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_98
timestamp 1
transform 1 0 10120 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_103
timestamp 1
transform 1 0 10580 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_113
timestamp 1
transform 1 0 11500 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_119
timestamp 1
transform 1 0 12052 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1636968456
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_169
timestamp 1
transform 1 0 16652 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_187
timestamp 1
transform 1 0 18308 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_21_210
timestamp 1
transform 1 0 20424 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_225
timestamp 1
transform 1 0 21804 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_21_243
timestamp 1636968456
transform 1 0 23460 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_255
timestamp 1
transform 1 0 24564 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_259
timestamp 1
transform 1 0 24932 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_263
timestamp 1
transform 1 0 25300 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_281
timestamp 1
transform 1 0 26956 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_287
timestamp 1
transform 1 0 27508 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_13
timestamp 1
transform 1 0 2300 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_19
timestamp 1
transform 1 0 2852 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_37
timestamp 1636968456
transform 1 0 4508 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_49
timestamp 1
transform 1 0 5612 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_57
timestamp 1
transform 1 0 6348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1636968456
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_85
timestamp 1
transform 1 0 8924 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_22_94
timestamp 1
transform 1 0 9752 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_106
timestamp 1636968456
transform 1 0 10856 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_118
timestamp 1
transform 1 0 11960 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_141
timestamp 1
transform 1 0 14076 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_154
timestamp 1
transform 1 0 15272 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_22_170
timestamp 1636968456
transform 1 0 16744 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_191
timestamp 1
transform 1 0 18676 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1636968456
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1636968456
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_226
timestamp 1
transform 1 0 21896 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_233
timestamp 1
transform 1 0 22540 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_237
timestamp 1
transform 1 0 22908 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_244
timestamp 1
transform 1 0 23552 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_22_256
timestamp 1636968456
transform 1 0 24656 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_268
timestamp 1
transform 1 0 25760 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_284
timestamp 1
transform 1 0 27232 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_3
timestamp 1
transform 1 0 1380 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_16
timestamp 1
transform 1 0 2576 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_20
timestamp 1
transform 1 0 2944 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_26
timestamp 1
transform 1 0 3496 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_44
timestamp 1
transform 1 0 5152 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_98
timestamp 1
transform 1 0 10120 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_104
timestamp 1
transform 1 0 10672 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_145
timestamp 1
transform 1 0 14444 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_165
timestamp 1
transform 1 0 16284 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_176
timestamp 1
transform 1 0 17296 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_180
timestamp 1
transform 1 0 17664 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_188
timestamp 1636968456
transform 1 0 18400 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_200
timestamp 1
transform 1 0 19504 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_207
timestamp 1
transform 1 0 20148 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_211
timestamp 1
transform 1 0 20516 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_233
timestamp 1636968456
transform 1 0 22540 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_245
timestamp 1
transform 1 0 23644 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_249
timestamp 1
transform 1 0 24012 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_263
timestamp 1636968456
transform 1 0 25300 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_275
timestamp 1
transform 1 0 26404 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_281
timestamp 1
transform 1 0 26956 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_287
timestamp 1
transform 1 0 27508 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_3
timestamp 1
transform 1 0 1380 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_26
timestamp 1
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_29
timestamp 1
transform 1 0 3772 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_45
timestamp 1
transform 1 0 5244 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_60
timestamp 1636968456
transform 1 0 6624 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_72
timestamp 1
transform 1 0 7728 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_81
timestamp 1
transform 1 0 8556 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1636968456
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1636968456
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1636968456
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_121
timestamp 1
transform 1 0 12236 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_129
timestamp 1
transform 1 0 12972 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_141
timestamp 1
transform 1 0 14076 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_149
timestamp 1
transform 1 0 14812 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_155
timestamp 1
transform 1 0 15364 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_191
timestamp 1
transform 1 0 18676 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_216
timestamp 1
transform 1 0 20976 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_228
timestamp 1
transform 1 0 22080 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_263
timestamp 1
transform 1 0 25300 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_276
timestamp 1636968456
transform 1 0 26496 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1636968456
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1636968456
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_27
timestamp 1
transform 1 0 3588 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_57
timestamp 1
transform 1 0 6348 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_65
timestamp 1
transform 1 0 7084 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_73
timestamp 1
transform 1 0 7820 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_88
timestamp 1
transform 1 0 9200 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_113
timestamp 1
transform 1 0 11500 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_119
timestamp 1
transform 1 0 12052 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_143
timestamp 1
transform 1 0 14260 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_156
timestamp 1636968456
transform 1 0 15456 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_175
timestamp 1636968456
transform 1 0 17204 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_187
timestamp 1636968456
transform 1 0 18308 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_199
timestamp 1636968456
transform 1 0 19412 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_211
timestamp 1636968456
transform 1 0 20516 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1636968456
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1636968456
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_249
timestamp 1
transform 1 0 24012 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_25_266
timestamp 1636968456
transform 1 0 25576 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_278
timestamp 1
transform 1 0 26680 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_281
timestamp 1
transform 1 0 26956 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_287
timestamp 1
transform 1 0 27508 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_3
timestamp 1
transform 1 0 1380 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_26_25
timestamp 1
transform 1 0 3404 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_29
timestamp 1
transform 1 0 3772 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_35
timestamp 1
transform 1 0 4324 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_39
timestamp 1
transform 1 0 4692 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_47
timestamp 1
transform 1 0 5428 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_63
timestamp 1636968456
transform 1 0 6900 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_75
timestamp 1
transform 1 0 8004 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_88
timestamp 1
transform 1 0 9200 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_100
timestamp 1
transform 1 0 10304 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_106
timestamp 1
transform 1 0 10856 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_126
timestamp 1
transform 1 0 12696 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_137
timestamp 1
transform 1 0 13708 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_161
timestamp 1636968456
transform 1 0 15916 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_173
timestamp 1
transform 1 0 17020 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_181
timestamp 1
transform 1 0 17756 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_193
timestamp 1
transform 1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_197
timestamp 1
transform 1 0 19228 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_212
timestamp 1
transform 1 0 20608 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_225
timestamp 1636968456
transform 1 0 21804 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_250
timestamp 1
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1636968456
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1636968456
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_277
timestamp 1
transform 1 0 26588 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_285
timestamp 1
transform 1 0 27324 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_33
timestamp 1
transform 1 0 4140 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_62
timestamp 1
transform 1 0 6808 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_77
timestamp 1
transform 1 0 8188 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_83
timestamp 1636968456
transform 1 0 8740 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_103
timestamp 1
transform 1 0 10580 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_120
timestamp 1
transform 1 0 12144 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_140
timestamp 1
transform 1 0 13984 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_163
timestamp 1
transform 1 0 16100 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_174
timestamp 1
transform 1 0 17112 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_200
timestamp 1
transform 1 0 19504 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_208
timestamp 1
transform 1 0 20240 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_245
timestamp 1636968456
transform 1 0 23644 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_281
timestamp 1
transform 1 0 26956 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_287
timestamp 1
transform 1 0 27508 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1636968456
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_15
timestamp 1
transform 1 0 2484 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_26
timestamp 1
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_29
timestamp 1
transform 1 0 3772 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_37
timestamp 1
transform 1 0 4508 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_42
timestamp 1
transform 1 0 4968 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_56
timestamp 1
transform 1 0 6256 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_63
timestamp 1
transform 1 0 6900 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_67
timestamp 1
transform 1 0 7268 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_76
timestamp 1
transform 1 0 8096 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_85
timestamp 1
transform 1 0 8924 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_91
timestamp 1
transform 1 0 9476 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_110
timestamp 1
transform 1 0 11224 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_114
timestamp 1
transform 1 0 11592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_119
timestamp 1
transform 1 0 12052 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_136
timestamp 1
transform 1 0 13616 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_197
timestamp 1
transform 1 0 19228 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_203
timestamp 1
transform 1 0 19780 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_208
timestamp 1636968456
transform 1 0 20240 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_220
timestamp 1636968456
transform 1 0 21344 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_232
timestamp 1
transform 1 0 22448 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_239
timestamp 1636968456
transform 1 0 23092 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_266
timestamp 1636968456
transform 1 0 25576 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_278
timestamp 1
transform 1 0 26680 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_286
timestamp 1
transform 1 0 27416 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_3
timestamp 1
transform 1 0 1380 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_11
timestamp 1
transform 1 0 2116 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_36
timestamp 1
transform 1 0 4416 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_98
timestamp 1
transform 1 0 10120 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_102
timestamp 1
transform 1 0 10488 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_113
timestamp 1
transform 1 0 11500 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_142
timestamp 1
transform 1 0 14168 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_225
timestamp 1
transform 1 0 21804 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_229
timestamp 1
transform 1 0 22172 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_250
timestamp 1
transform 1 0 24104 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_267
timestamp 1636968456
transform 1 0 25668 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_281
timestamp 1
transform 1 0 26956 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_287
timestamp 1
transform 1 0 27508 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1636968456
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1636968456
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_29
timestamp 1
transform 1 0 3772 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_67
timestamp 1636968456
transform 1 0 7268 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_79
timestamp 1
transform 1 0 8372 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_89
timestamp 1
transform 1 0 9292 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_93
timestamp 1
transform 1 0 9660 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_125
timestamp 1
transform 1 0 12604 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_141
timestamp 1
transform 1 0 14076 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_176
timestamp 1
transform 1 0 17296 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_180
timestamp 1
transform 1 0 17664 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_197
timestamp 1
transform 1 0 19228 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_205
timestamp 1
transform 1 0 19964 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_210
timestamp 1
transform 1 0 20424 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_218
timestamp 1
transform 1 0 21160 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_225
timestamp 1
transform 1 0 21804 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_233
timestamp 1
transform 1 0 22540 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_239
timestamp 1636968456
transform 1 0 23092 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1636968456
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_265
timestamp 1636968456
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_277
timestamp 1
transform 1 0 26588 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_285
timestamp 1
transform 1 0 27324 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_19
timestamp 1
transform 1 0 2852 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_27
timestamp 1
transform 1 0 3588 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_45
timestamp 1
transform 1 0 5244 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_65
timestamp 1
transform 1 0 7084 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_94
timestamp 1
transform 1 0 9752 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_108
timestamp 1
transform 1 0 11040 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_136
timestamp 1
transform 1 0 13616 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_146
timestamp 1
transform 1 0 14536 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_159
timestamp 1
transform 1 0 15732 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_177
timestamp 1636968456
transform 1 0 17388 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_195
timestamp 1
transform 1 0 19044 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_31_216
timestamp 1
transform 1 0 20976 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1636968456
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_242
timestamp 1
transform 1 0 23368 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_255
timestamp 1
transform 1 0 24564 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_263
timestamp 1636968456
transform 1 0 25300 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_275
timestamp 1
transform 1 0 26404 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_281
timestamp 1
transform 1 0 26956 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_287
timestamp 1
transform 1 0 27508 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_6
timestamp 1
transform 1 0 1656 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_29
timestamp 1
transform 1 0 3772 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_33
timestamp 1
transform 1 0 4140 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_89
timestamp 1
transform 1 0 9292 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_95
timestamp 1
transform 1 0 9844 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_99
timestamp 1
transform 1 0 10212 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_123
timestamp 1
transform 1 0 12420 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_207
timestamp 1
transform 1 0 20148 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_32_232
timestamp 1
transform 1 0 22448 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_260
timestamp 1636968456
transform 1 0 25024 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_272
timestamp 1636968456
transform 1 0 26128 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_284
timestamp 1
transform 1 0 27232 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1636968456
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_15
timestamp 1
transform 1 0 2484 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_25
timestamp 1
transform 1 0 3404 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_29
timestamp 1
transform 1 0 3772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_52
timestamp 1
transform 1 0 5888 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_57
timestamp 1
transform 1 0 6348 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_64
timestamp 1636968456
transform 1 0 6992 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_76
timestamp 1
transform 1 0 8096 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_82
timestamp 1
transform 1 0 8648 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_90
timestamp 1
transform 1 0 9384 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_108
timestamp 1
transform 1 0 11040 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_130
timestamp 1
transform 1 0 13064 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_142
timestamp 1
transform 1 0 14168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_147
timestamp 1
transform 1 0 14628 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_155
timestamp 1
transform 1 0 15364 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_164
timestamp 1
transform 1 0 16192 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1636968456
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1636968456
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_193
timestamp 1636968456
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_205
timestamp 1
transform 1 0 19964 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_212
timestamp 1636968456
transform 1 0 20608 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1636968456
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_237
timestamp 1
transform 1 0 22908 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_245
timestamp 1
transform 1 0 23644 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_253
timestamp 1636968456
transform 1 0 24380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_265
timestamp 1636968456
transform 1 0 25484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_277
timestamp 1
transform 1 0 26588 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_33_281
timestamp 1
transform 1 0 26956 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_287
timestamp 1
transform 1 0 27508 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_53
timestamp 1
transform 1 0 5980 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_64
timestamp 1
transform 1 0 6992 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_74
timestamp 1
transform 1 0 7912 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_82
timestamp 1
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_88
timestamp 1
transform 1 0 9200 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_106
timestamp 1636968456
transform 1 0 10856 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_118
timestamp 1636968456
transform 1 0 11960 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_130
timestamp 1
transform 1 0 13064 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_138
timestamp 1
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_141
timestamp 1
transform 1 0 14076 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_154
timestamp 1
transform 1 0 15272 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_158
timestamp 1
transform 1 0 15640 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_164
timestamp 1
transform 1 0 16192 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_34_180
timestamp 1
transform 1 0 17664 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_201
timestamp 1
transform 1 0 19596 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_224
timestamp 1
transform 1 0 21712 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_34_244
timestamp 1
transform 1 0 23552 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1636968456
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1636968456
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_277
timestamp 1
transform 1 0 26588 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_285
timestamp 1
transform 1 0 27324 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_35_6
timestamp 1
transform 1 0 1656 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_12
timestamp 1
transform 1 0 2208 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_29
timestamp 1
transform 1 0 3772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_38
timestamp 1
transform 1 0 4600 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_57
timestamp 1
transform 1 0 6348 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_68
timestamp 1
transform 1 0 7360 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_88
timestamp 1636968456
transform 1 0 9200 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_100
timestamp 1636968456
transform 1 0 10304 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_113
timestamp 1
transform 1 0 11500 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_140
timestamp 1
transform 1 0 13984 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_180
timestamp 1
transform 1 0 17664 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_35_192
timestamp 1
transform 1 0 18768 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_200
timestamp 1
transform 1 0 19504 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_209
timestamp 1636968456
transform 1 0 20332 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_221
timestamp 1
transform 1 0 21436 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_236
timestamp 1
transform 1 0 22816 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_248
timestamp 1636968456
transform 1 0 23920 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_260
timestamp 1636968456
transform 1 0 25024 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_272
timestamp 1
transform 1 0 26128 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_35_281
timestamp 1
transform 1 0 26956 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_287
timestamp 1
transform 1 0 27508 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_19
timestamp 1
transform 1 0 2852 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_71
timestamp 1
transform 1 0 7636 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_76
timestamp 1
transform 1 0 8096 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_81
timestamp 1
transform 1 0 8556 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_85
timestamp 1
transform 1 0 8924 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_93
timestamp 1
transform 1 0 9660 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_102
timestamp 1
transform 1 0 10488 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_110
timestamp 1
transform 1 0 11224 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_119
timestamp 1
transform 1 0 12052 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_148
timestamp 1
transform 1 0 14720 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_156
timestamp 1
transform 1 0 15456 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_160
timestamp 1
transform 1 0 15824 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_168
timestamp 1
transform 1 0 16560 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_194
timestamp 1
transform 1 0 18952 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_217
timestamp 1636968456
transform 1 0 21068 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_229
timestamp 1636968456
transform 1 0 22172 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_241
timestamp 1
transform 1 0 23276 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_249
timestamp 1
transform 1 0 24012 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1636968456
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1636968456
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_277
timestamp 1
transform 1 0 26588 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_285
timestamp 1
transform 1 0 27324 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_3
timestamp 1
transform 1 0 1380 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_11
timestamp 1
transform 1 0 2116 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_28
timestamp 1
transform 1 0 3680 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_38
timestamp 1
transform 1 0 4600 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_57
timestamp 1
transform 1 0 6348 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_63
timestamp 1
transform 1 0 6900 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_67
timestamp 1
transform 1 0 7268 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_128
timestamp 1
transform 1 0 12880 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_138
timestamp 1
transform 1 0 13800 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_209
timestamp 1
transform 1 0 20332 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_213
timestamp 1
transform 1 0 20700 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_232
timestamp 1636968456
transform 1 0 22448 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_244
timestamp 1636968456
transform 1 0 23552 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_256
timestamp 1636968456
transform 1 0 24656 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_268
timestamp 1636968456
transform 1 0 25760 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_281
timestamp 1
transform 1 0 26956 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_287
timestamp 1
transform 1 0 27508 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1636968456
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_15
timestamp 1
transform 1 0 2484 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_25
timestamp 1
transform 1 0 3404 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_33
timestamp 1636968456
transform 1 0 4140 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_74
timestamp 1
transform 1 0 7912 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_82
timestamp 1
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_89
timestamp 1
transform 1 0 9292 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1636968456
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1636968456
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_121
timestamp 1
transform 1 0 12236 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_38_149
timestamp 1
transform 1 0 14812 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_38_175
timestamp 1
transform 1 0 17204 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_193
timestamp 1
transform 1 0 18860 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_38_224
timestamp 1636968456
transform 1 0 21712 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_236
timestamp 1636968456
transform 1 0 22816 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_248
timestamp 1
transform 1 0 23920 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1636968456
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_265
timestamp 1636968456
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_277
timestamp 1
transform 1 0 26588 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_285
timestamp 1
transform 1 0 27324 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_10
timestamp 1
transform 1 0 2024 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_14
timestamp 1
transform 1 0 2392 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_23
timestamp 1
transform 1 0 3220 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_57
timestamp 1
transform 1 0 6348 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_63
timestamp 1
transform 1 0 6900 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_71
timestamp 1
transform 1 0 7636 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_75
timestamp 1
transform 1 0 8004 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_80
timestamp 1636968456
transform 1 0 8464 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_92
timestamp 1
transform 1 0 9568 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_121
timestamp 1
transform 1 0 12236 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_153
timestamp 1
transform 1 0 15180 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_165
timestamp 1
transform 1 0 16284 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1636968456
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1636968456
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_193
timestamp 1
transform 1 0 18860 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_204
timestamp 1636968456
transform 1 0 19872 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_216
timestamp 1
transform 1 0 20976 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1636968456
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_237
timestamp 1636968456
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_249
timestamp 1636968456
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_261
timestamp 1636968456
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_281
timestamp 1
transform 1 0 26956 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_287
timestamp 1
transform 1 0 27508 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1636968456
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_41
timestamp 1
transform 1 0 4876 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_49
timestamp 1
transform 1 0 5612 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_63
timestamp 1
transform 1 0 6900 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_71
timestamp 1
transform 1 0 7636 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_105
timestamp 1
transform 1 0 10764 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_136
timestamp 1
transform 1 0 13616 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_180
timestamp 1
transform 1 0 17664 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_188
timestamp 1
transform 1 0 18400 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_193
timestamp 1
transform 1 0 18860 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_197
timestamp 1
transform 1 0 19228 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_201
timestamp 1
transform 1 0 19596 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_226
timestamp 1636968456
transform 1 0 21896 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_238
timestamp 1636968456
transform 1 0 23000 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_250
timestamp 1
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_253
timestamp 1636968456
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_265
timestamp 1636968456
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_277
timestamp 1
transform 1 0 26588 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_285
timestamp 1
transform 1 0 27324 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_41_7
timestamp 1
transform 1 0 1748 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_11
timestamp 1
transform 1 0 2116 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_41_22
timestamp 1
transform 1 0 3128 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_41_39
timestamp 1
transform 1 0 4692 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_45
timestamp 1
transform 1 0 5244 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_41_50
timestamp 1
transform 1 0 5704 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_54
timestamp 1
transform 1 0 6072 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_98
timestamp 1
transform 1 0 10120 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_102
timestamp 1
transform 1 0 10488 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_110
timestamp 1
transform 1 0 11224 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_121
timestamp 1
transform 1 0 12236 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_148
timestamp 1
transform 1 0 14720 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_169
timestamp 1
transform 1 0 16652 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_173
timestamp 1
transform 1 0 17020 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_214
timestamp 1
transform 1 0 20792 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_222
timestamp 1
transform 1 0 21528 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1636968456
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1636968456
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1636968456
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_261
timestamp 1636968456
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_281
timestamp 1
transform 1 0 26956 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_287
timestamp 1
transform 1 0 27508 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_10
timestamp 1636968456
transform 1 0 2024 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_22
timestamp 1
transform 1 0 3128 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_63
timestamp 1
transform 1 0 6900 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_75
timestamp 1
transform 1 0 8004 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_79
timestamp 1
transform 1 0 8372 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_85
timestamp 1
transform 1 0 8924 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_95
timestamp 1
transform 1 0 9844 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_42_114
timestamp 1
transform 1 0 11592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1636968456
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_153
timestamp 1
transform 1 0 15180 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_158
timestamp 1
transform 1 0 15640 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_162
timestamp 1
transform 1 0 16008 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_168
timestamp 1636968456
transform 1 0 16560 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_180
timestamp 1636968456
transform 1 0 17664 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_192
timestamp 1
transform 1 0 18768 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_197
timestamp 1
transform 1 0 19228 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_226
timestamp 1636968456
transform 1 0 21896 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_238
timestamp 1636968456
transform 1 0 23000 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_250
timestamp 1
transform 1 0 24104 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1636968456
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1636968456
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_277
timestamp 1
transform 1 0 26588 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_285
timestamp 1
transform 1 0 27324 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_43_3
timestamp 1
transform 1 0 1380 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_43_20
timestamp 1
transform 1 0 2944 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_43_39
timestamp 1
transform 1 0 4692 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_43_49
timestamp 1
transform 1 0 5612 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_43_62
timestamp 1
transform 1 0 6808 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_69
timestamp 1
transform 1 0 7452 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_81
timestamp 1
transform 1 0 8556 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_87
timestamp 1
transform 1 0 9108 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1636968456
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_105
timestamp 1
transform 1 0 10764 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_113
timestamp 1
transform 1 0 11500 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_43_139
timestamp 1
transform 1 0 13892 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_147
timestamp 1
transform 1 0 14628 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_155
timestamp 1
transform 1 0 15364 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_43_169
timestamp 1
transform 1 0 16652 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_187
timestamp 1636968456
transform 1 0 18308 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_199
timestamp 1
transform 1 0 19412 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_43_221
timestamp 1
transform 1 0 21436 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1636968456
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1636968456
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1636968456
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1636968456
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_281
timestamp 1
transform 1 0 26956 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_287
timestamp 1
transform 1 0 27508 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_11
timestamp 1
transform 1 0 2116 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_44_22
timestamp 1
transform 1 0 3128 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_44_29
timestamp 1
transform 1 0 3772 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_46
timestamp 1
transform 1 0 5336 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_71
timestamp 1
transform 1 0 7636 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_44_85
timestamp 1
transform 1 0 8924 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_121
timestamp 1
transform 1 0 12236 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_157
timestamp 1
transform 1 0 15548 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_168
timestamp 1
transform 1 0 16560 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_192
timestamp 1
transform 1 0 18768 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_197
timestamp 1
transform 1 0 19228 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_204
timestamp 1636968456
transform 1 0 19872 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_216
timestamp 1636968456
transform 1 0 20976 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_228
timestamp 1636968456
transform 1 0 22080 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_240
timestamp 1636968456
transform 1 0 23184 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1636968456
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1636968456
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_277
timestamp 1
transform 1 0 26588 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_285
timestamp 1
transform 1 0 27324 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_45_3
timestamp 1
transform 1 0 1380 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_45_15
timestamp 1
transform 1 0 2484 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_24
timestamp 1636968456
transform 1 0 3312 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_36
timestamp 1
transform 1 0 4416 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_45_42
timestamp 1
transform 1 0 4968 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_46
timestamp 1
transform 1 0 5336 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_54
timestamp 1
transform 1 0 6072 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_57
timestamp 1
transform 1 0 6348 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_63
timestamp 1
transform 1 0 6900 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_67
timestamp 1
transform 1 0 7268 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_73
timestamp 1
transform 1 0 7820 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_79
timestamp 1
transform 1 0 8372 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_87
timestamp 1
transform 1 0 9108 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_92
timestamp 1
transform 1 0 9568 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_104
timestamp 1
transform 1 0 10672 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_45_113
timestamp 1
transform 1 0 11500 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_121
timestamp 1
transform 1 0 12236 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_148
timestamp 1
transform 1 0 14720 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_45_165
timestamp 1
transform 1 0 16284 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_169
timestamp 1
transform 1 0 16652 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_173
timestamp 1
transform 1 0 17020 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_180
timestamp 1
transform 1 0 17664 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_186
timestamp 1
transform 1 0 18216 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_219
timestamp 1
transform 1 0 21252 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1636968456
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1636968456
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1636968456
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1636968456
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_281
timestamp 1
transform 1 0 26956 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_287
timestamp 1
transform 1 0 27508 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_46_19
timestamp 1
transform 1 0 2852 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_43
timestamp 1
transform 1 0 5060 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_51
timestamp 1
transform 1 0 5796 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_60
timestamp 1
transform 1 0 6624 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_46_85
timestamp 1
transform 1 0 8924 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_108
timestamp 1
transform 1 0 11040 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_126
timestamp 1
transform 1 0 12696 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_149
timestamp 1
transform 1 0 14812 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_160
timestamp 1
transform 1 0 15824 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_167
timestamp 1
transform 1 0 16468 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_173
timestamp 1
transform 1 0 17020 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1636968456
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1636968456
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_221
timestamp 1636968456
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_233
timestamp 1636968456
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1636968456
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1636968456
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_277
timestamp 1
transform 1 0 26588 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_285
timestamp 1
transform 1 0 27324 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_47_3
timestamp 1
transform 1 0 1380 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_47_9
timestamp 1
transform 1 0 1932 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_47_45
timestamp 1
transform 1 0 5244 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_64
timestamp 1
transform 1 0 6992 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_70
timestamp 1
transform 1 0 7544 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_47_113
timestamp 1
transform 1 0 11500 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_47_124
timestamp 1
transform 1 0 12512 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_141
timestamp 1
transform 1 0 14076 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_161
timestamp 1
transform 1 0 15916 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_209
timestamp 1636968456
transform 1 0 20332 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_221
timestamp 1
transform 1 0 21436 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1636968456
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_237
timestamp 1636968456
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_249
timestamp 1636968456
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_261
timestamp 1636968456
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_281
timestamp 1
transform 1 0 26956 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_287
timestamp 1
transform 1 0 27508 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1636968456
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_15
timestamp 1
transform 1 0 2484 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_23
timestamp 1
transform 1 0 3220 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_29
timestamp 1
transform 1 0 3772 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_37
timestamp 1
transform 1 0 4508 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_44
timestamp 1
transform 1 0 5152 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_77
timestamp 1
transform 1 0 8188 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1636968456
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_109
timestamp 1
transform 1 0 11132 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_48_113
timestamp 1
transform 1 0 11500 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_121
timestamp 1
transform 1 0 12236 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_125
timestamp 1636968456
transform 1 0 12604 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_137
timestamp 1
transform 1 0 13708 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1636968456
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_153
timestamp 1636968456
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_165
timestamp 1
transform 1 0 16284 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_169
timestamp 1
transform 1 0 16652 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_176
timestamp 1636968456
transform 1 0 17296 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_188
timestamp 1
transform 1 0 18400 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1636968456
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_209
timestamp 1636968456
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_221
timestamp 1
transform 1 0 21436 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_225
timestamp 1636968456
transform 1 0 21804 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_237
timestamp 1636968456
transform 1 0 22908 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_249
timestamp 1
transform 1 0 24012 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1636968456
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1636968456
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_277
timestamp 1
transform 1 0 26588 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_48_281
timestamp 1
transform 1 0 26956 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_287
timestamp 1
transform 1 0 27508 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 1
transform -1 0 9660 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1
transform -1 0 3588 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1
transform -1 0 3404 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1
transform -1 0 3404 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1
transform -1 0 4600 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1
transform -1 0 4600 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1
transform 1 0 3864 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1
transform 1 0 7268 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1
transform -1 0 20792 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1
transform -1 0 18676 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1
transform -1 0 20792 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1
transform -1 0 12512 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1
transform -1 0 21896 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1
transform 1 0 19964 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1
transform -1 0 20332 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1
transform -1 0 14812 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1
transform -1 0 13616 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1
transform -1 0 18492 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1
transform 1 0 12420 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1
transform -1 0 12788 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1
transform -1 0 18860 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1
transform -1 0 21896 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1
transform -1 0 12236 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1
transform 1 0 11500 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1
transform -1 0 14812 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1
transform 1 0 13156 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1
transform -1 0 18952 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1
transform -1 0 17664 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1
transform -1 0 15824 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1
transform -1 0 18492 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1
transform -1 0 20332 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1
transform -1 0 14628 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1
transform -1 0 3588 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1
transform -1 0 10672 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1
transform -1 0 9844 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 1
transform 1 0 9936 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 1
transform -1 0 3680 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 1
transform -1 0 13800 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 1
transform -1 0 16284 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 1
transform 1 0 12972 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 1
transform -1 0 4508 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 1
transform -1 0 20332 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 1
transform -1 0 14812 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 1
transform 1 0 9660 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 1
transform -1 0 18308 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 1
transform 1 0 13248 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 1
transform -1 0 9384 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 1
transform -1 0 15640 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1
transform 1 0 8464 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1
transform 1 0 1748 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1
transform -1 0 1656 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1
transform -1 0 1656 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  intro_2_stopwatch_52
timestamp 1
transform 1 0 1380 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  intro_2_stopwatch_53
timestamp 1
transform 1 0 3312 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  intro_2_stopwatch_54
timestamp 1
transform -1 0 27600 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  max_cap21
timestamp 1
transform -1 0 20240 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  max_cap29
timestamp 1
transform 1 0 7544 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output5
timestamp 1
transform -1 0 2116 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp 1
transform 1 0 9660 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp 1
transform -1 0 1748 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp 1
transform -1 0 1748 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 1
transform 1 0 5888 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1
transform -1 0 1748 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 1
transform -1 0 1748 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1
transform 1 0 6348 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 1
transform 1 0 7176 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_49
timestamp 1
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1
transform -1 0 27876 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_50
timestamp 1
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1
transform -1 0 27876 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_51
timestamp 1
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1
transform -1 0 27876 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_52
timestamp 1
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1
transform -1 0 27876 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_53
timestamp 1
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1
transform -1 0 27876 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_54
timestamp 1
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1
transform -1 0 27876 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_55
timestamp 1
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1
transform -1 0 27876 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_56
timestamp 1
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1
transform -1 0 27876 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_57
timestamp 1
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1
transform -1 0 27876 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_58
timestamp 1
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1
transform -1 0 27876 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_59
timestamp 1
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1
transform -1 0 27876 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_60
timestamp 1
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1
transform -1 0 27876 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_61
timestamp 1
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1
transform -1 0 27876 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_62
timestamp 1
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1
transform -1 0 27876 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_63
timestamp 1
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1
transform -1 0 27876 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_64
timestamp 1
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1
transform -1 0 27876 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_65
timestamp 1
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1
transform -1 0 27876 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_66
timestamp 1
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1
transform -1 0 27876 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_67
timestamp 1
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1
transform -1 0 27876 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_68
timestamp 1
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1
transform -1 0 27876 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_69
timestamp 1
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1
transform -1 0 27876 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_70
timestamp 1
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1
transform -1 0 27876 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_71
timestamp 1
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1
transform -1 0 27876 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_72
timestamp 1
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1
transform -1 0 27876 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_73
timestamp 1
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1
transform -1 0 27876 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_74
timestamp 1
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1
transform -1 0 27876 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_75
timestamp 1
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1
transform -1 0 27876 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_76
timestamp 1
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1
transform -1 0 27876 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_77
timestamp 1
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1
transform -1 0 27876 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_78
timestamp 1
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1
transform -1 0 27876 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_79
timestamp 1
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1
transform -1 0 27876 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_80
timestamp 1
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1
transform -1 0 27876 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_81
timestamp 1
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1
transform -1 0 27876 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_82
timestamp 1
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1
transform -1 0 27876 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_83
timestamp 1
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 1
transform -1 0 27876 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_84
timestamp 1
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 1
transform -1 0 27876 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_85
timestamp 1
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 1
transform -1 0 27876 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_86
timestamp 1
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 1
transform -1 0 27876 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_87
timestamp 1
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 1
transform -1 0 27876 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_88
timestamp 1
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp 1
transform -1 0 27876 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_89
timestamp 1
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp 1
transform -1 0 27876 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_90
timestamp 1
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp 1
transform -1 0 27876 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Left_91
timestamp 1
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Right_42
timestamp 1
transform -1 0 27876 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Left_92
timestamp 1
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Right_43
timestamp 1
transform -1 0 27876 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Left_93
timestamp 1
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Right_44
timestamp 1
transform -1 0 27876 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Left_94
timestamp 1
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Right_45
timestamp 1
transform -1 0 27876 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Left_95
timestamp 1
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Right_46
timestamp 1
transform -1 0 27876 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Left_96
timestamp 1
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Right_47
timestamp 1
transform -1 0 27876 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Left_97
timestamp 1
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Right_48
timestamp 1
transform -1 0 27876 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_98
timestamp 1
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_99
timestamp 1
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_100
timestamp 1
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_101
timestamp 1
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_102
timestamp 1
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_103
timestamp 1
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_104
timestamp 1
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_105
timestamp 1
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_106
timestamp 1
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_107
timestamp 1
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_108
timestamp 1
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_109
timestamp 1
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_110
timestamp 1
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_111
timestamp 1
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_112
timestamp 1
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_113
timestamp 1
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_114
timestamp 1
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_115
timestamp 1
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_116
timestamp 1
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_117
timestamp 1
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_118
timestamp 1
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_119
timestamp 1
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_120
timestamp 1
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_121
timestamp 1
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_122
timestamp 1
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_123
timestamp 1
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_124
timestamp 1
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_125
timestamp 1
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_126
timestamp 1
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_127
timestamp 1
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_128
timestamp 1
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_129
timestamp 1
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_130
timestamp 1
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_131
timestamp 1
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_132
timestamp 1
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_133
timestamp 1
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_134
timestamp 1
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_135
timestamp 1
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_136
timestamp 1
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_137
timestamp 1
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_138
timestamp 1
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_139
timestamp 1
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_140
timestamp 1
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_141
timestamp 1
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_142
timestamp 1
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_143
timestamp 1
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_144
timestamp 1
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_145
timestamp 1
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_146
timestamp 1
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_147
timestamp 1
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_148
timestamp 1
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_149
timestamp 1
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_150
timestamp 1
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_151
timestamp 1
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_152
timestamp 1
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_153
timestamp 1
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_154
timestamp 1
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_155
timestamp 1
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_156
timestamp 1
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_157
timestamp 1
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_158
timestamp 1
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_159
timestamp 1
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_160
timestamp 1
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_161
timestamp 1
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_162
timestamp 1
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_163
timestamp 1
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_164
timestamp 1
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_165
timestamp 1
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_166
timestamp 1
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_167
timestamp 1
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_168
timestamp 1
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_169
timestamp 1
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_170
timestamp 1
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_171
timestamp 1
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_172
timestamp 1
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_173
timestamp 1
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_174
timestamp 1
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_175
timestamp 1
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_176
timestamp 1
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_177
timestamp 1
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_178
timestamp 1
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_179
timestamp 1
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_180
timestamp 1
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_181
timestamp 1
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_182
timestamp 1
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_183
timestamp 1
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_184
timestamp 1
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_185
timestamp 1
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_186
timestamp 1
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_187
timestamp 1
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_188
timestamp 1
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_189
timestamp 1
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_190
timestamp 1
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_191
timestamp 1
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_192
timestamp 1
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_193
timestamp 1
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_194
timestamp 1
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_195
timestamp 1
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_196
timestamp 1
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_197
timestamp 1
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_198
timestamp 1
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_199
timestamp 1
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_200
timestamp 1
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_201
timestamp 1
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_202
timestamp 1
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_203
timestamp 1
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_204
timestamp 1
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_205
timestamp 1
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_206
timestamp 1
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_207
timestamp 1
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_208
timestamp 1
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_209
timestamp 1
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_210
timestamp 1
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_211
timestamp 1
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_212
timestamp 1
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_213
timestamp 1
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_214
timestamp 1
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_215
timestamp 1
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_216
timestamp 1
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_217
timestamp 1
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_218
timestamp 1
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_219
timestamp 1
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_220
timestamp 1
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_221
timestamp 1
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_222
timestamp 1
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_223
timestamp 1
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_224
timestamp 1
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_225
timestamp 1
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_226
timestamp 1
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_227
timestamp 1
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_228
timestamp 1
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_229
timestamp 1
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_230
timestamp 1
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_231
timestamp 1
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_232
timestamp 1
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_233
timestamp 1
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_234
timestamp 1
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_235
timestamp 1
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_236
timestamp 1
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_237
timestamp 1
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_238
timestamp 1
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_239
timestamp 1
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_240
timestamp 1
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_241
timestamp 1
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_242
timestamp 1
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_243
timestamp 1
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_244
timestamp 1
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_245
timestamp 1
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_246
timestamp 1
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_247
timestamp 1
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_248
timestamp 1
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_249
timestamp 1
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_250
timestamp 1
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_251
timestamp 1
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_252
timestamp 1
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_253
timestamp 1
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_254
timestamp 1
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_255
timestamp 1
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_256
timestamp 1
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_257
timestamp 1
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_258
timestamp 1
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_259
timestamp 1
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_260
timestamp 1
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_261
timestamp 1
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_262
timestamp 1
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_263
timestamp 1
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_264
timestamp 1
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_265
timestamp 1
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_266
timestamp 1
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_267
timestamp 1
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_268
timestamp 1
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_269
timestamp 1
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_270
timestamp 1
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_271
timestamp 1
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_272
timestamp 1
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_273
timestamp 1
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_274
timestamp 1
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_275
timestamp 1
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_276
timestamp 1
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_277
timestamp 1
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_278
timestamp 1
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_279
timestamp 1
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_280
timestamp 1
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_281
timestamp 1
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_282
timestamp 1
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_283
timestamp 1
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_284
timestamp 1
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_285
timestamp 1
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_286
timestamp 1
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_287
timestamp 1
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_288
timestamp 1
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_289
timestamp 1
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_290
timestamp 1
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_291
timestamp 1
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_292
timestamp 1
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_293
timestamp 1
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_294
timestamp 1
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_295
timestamp 1
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_296
timestamp 1
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_297
timestamp 1
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_298
timestamp 1
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_299
timestamp 1
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_300
timestamp 1
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_301
timestamp 1
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_302
timestamp 1
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_303
timestamp 1
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_304
timestamp 1
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_305
timestamp 1
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_306
timestamp 1
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_307
timestamp 1
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_308
timestamp 1
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_309
timestamp 1
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_310
timestamp 1
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_311
timestamp 1
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_312
timestamp 1
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_313
timestamp 1
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_314
timestamp 1
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_315
timestamp 1
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_316
timestamp 1
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_317
timestamp 1
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_318
timestamp 1
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_319
timestamp 1
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_320
timestamp 1
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_321
timestamp 1
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_322
timestamp 1
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_323
timestamp 1
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_324
timestamp 1
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_325
timestamp 1
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_326
timestamp 1
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_327
timestamp 1
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_328
timestamp 1
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_329
timestamp 1
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_330
timestamp 1
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_331
timestamp 1
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_332
timestamp 1
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_333
timestamp 1
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_334
timestamp 1
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_335
timestamp 1
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_336
timestamp 1
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_337
timestamp 1
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_338
timestamp 1
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_339
timestamp 1
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_340
timestamp 1
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_341
timestamp 1
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_342
timestamp 1
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_343
timestamp 1
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_344
timestamp 1
transform 1 0 6256 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_345
timestamp 1
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_346
timestamp 1
transform 1 0 11408 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_347
timestamp 1
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_348
timestamp 1
transform 1 0 16560 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_349
timestamp 1
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_350
timestamp 1
transform 1 0 21712 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_351
timestamp 1
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_352
timestamp 1
transform 1 0 26864 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  wire38
timestamp 1
transform -1 0 6072 0 1 23936
box -38 -48 314 592
<< labels >>
flabel metal2 s 8390 30364 8446 31164 0 FreeSans 224 90 0 0 BTN[0]
port 0 nsew signal input
flabel metal3 s 0 23128 800 23248 0 FreeSans 480 0 0 0 BTN[1]
port 1 nsew signal input
flabel metal3 s 0 19728 800 19848 0 FreeSans 480 0 0 0 BTN[2]
port 2 nsew signal input
flabel metal3 s 0 21088 800 21208 0 FreeSans 480 0 0 0 BTN[3]
port 3 nsew signal input
flabel metal3 s 0 27888 800 28008 0 FreeSans 480 0 0 0 CLK_10MHZ
port 4 nsew signal input
flabel metal3 s 0 26528 800 26648 0 FreeSans 480 0 0 0 D0_AN_0
port 5 nsew signal output
flabel metal2 s 9034 30364 9090 31164 0 FreeSans 224 90 0 0 D0_AN_1
port 6 nsew signal output
flabel metal3 s 0 2728 800 2848 0 FreeSans 480 0 0 0 D0_AN_2
port 7 nsew signal output
flabel metal2 s 3238 30364 3294 31164 0 FreeSans 224 90 0 0 D0_AN_3
port 8 nsew signal output
flabel metal3 s 0 25168 800 25288 0 FreeSans 480 0 0 0 D0_SEG[0]
port 9 nsew signal output
flabel metal3 s 0 23808 800 23928 0 FreeSans 480 0 0 0 D0_SEG[1]
port 10 nsew signal output
flabel metal2 s 5814 30364 5870 31164 0 FreeSans 224 90 0 0 D0_SEG[2]
port 11 nsew signal output
flabel metal3 s 0 25848 800 25968 0 FreeSans 480 0 0 0 D0_SEG[3]
port 12 nsew signal output
flabel metal3 s 0 24488 800 24608 0 FreeSans 480 0 0 0 D0_SEG[4]
port 13 nsew signal output
flabel metal2 s 6458 30364 6514 31164 0 FreeSans 224 90 0 0 D0_SEG[5]
port 14 nsew signal output
flabel metal2 s 7102 30364 7158 31164 0 FreeSans 224 90 0 0 D0_SEG[6]
port 15 nsew signal output
flabel metal3 s 28220 2728 29020 2848 0 FreeSans 480 0 0 0 D0_SEG[7]
port 16 nsew signal output
flabel metal4 s 4868 2128 5188 28880 0 FreeSans 1920 90 0 0 VGND
port 17 nsew ground bidirectional
flabel metal4 s 4208 2128 4528 28880 0 FreeSans 1920 90 0 0 VPWR
port 18 nsew power bidirectional
rlabel metal1 14490 28288 14490 28288 0 VGND
rlabel metal1 14490 28832 14490 28832 0 VPWR
rlabel metal1 8556 28526 8556 28526 0 BTN[0]
rlabel metal3 1326 23188 1326 23188 0 BTN[1]
rlabel metal3 751 19788 751 19788 0 BTN[2]
rlabel metal3 751 21148 751 21148 0 BTN[3]
rlabel metal3 1004 27948 1004 27948 0 CLK_10MHZ
rlabel metal1 1564 26554 1564 26554 0 D0_AN_0
rlabel metal1 9476 28730 9476 28730 0 D0_AN_1
rlabel metal3 751 25228 751 25228 0 D0_SEG[0]
rlabel metal1 1380 23834 1380 23834 0 D0_SEG[1]
rlabel metal1 5980 28730 5980 28730 0 D0_SEG[2]
rlabel metal3 1096 25908 1096 25908 0 D0_SEG[3]
rlabel metal3 751 24548 751 24548 0 D0_SEG[4]
rlabel metal1 6532 28730 6532 28730 0 D0_SEG[5]
rlabel metal1 7268 28186 7268 28186 0 D0_SEG[6]
rlabel metal2 18722 24582 18722 24582 0 _0000_
rlabel metal2 19826 23868 19826 23868 0 _0001_
rlabel metal1 20511 25194 20511 25194 0 _0002_
rlabel metal1 18660 27030 18660 27030 0 _0003_
rlabel metal2 16790 27812 16790 27812 0 _0004_
rlabel metal1 17986 27574 17986 27574 0 _0005_
rlabel metal1 18036 26350 18036 26350 0 _0006_
rlabel metal2 16882 24582 16882 24582 0 _0007_
rlabel via1 15318 23851 15318 23851 0 _0008_
rlabel metal2 14674 23970 14674 23970 0 _0009_
rlabel metal1 14152 26282 14152 26282 0 _0010_
rlabel metal1 14720 26894 14720 26894 0 _0011_
rlabel metal1 12824 28050 12824 28050 0 _0012_
rlabel metal2 12466 24786 12466 24786 0 _0013_
rlabel metal2 11270 26146 11270 26146 0 _0014_
rlabel metal1 11444 27438 11444 27438 0 _0015_
rlabel metal1 7728 22202 7728 22202 0 _0016_
rlabel metal2 7038 19618 7038 19618 0 _0017_
rlabel metal1 5285 22610 5285 22610 0 _0018_
rlabel metal1 9522 20570 9522 20570 0 _0019_
rlabel metal1 9598 22678 9598 22678 0 _0020_
rlabel metal2 10994 24446 10994 24446 0 _0021_
rlabel metal2 10810 24106 10810 24106 0 _0022_
rlabel metal1 12642 21590 12642 21590 0 _0023_
rlabel metal1 12829 23766 12829 23766 0 _0024_
rlabel metal1 14724 22678 14724 22678 0 _0025_
rlabel metal1 11720 20434 11720 20434 0 _0026_
rlabel metal1 18906 21896 18906 21896 0 _0027_
rlabel metal2 18998 22882 18998 22882 0 _0028_
rlabel metal2 17342 22610 17342 22610 0 _0029_
rlabel metal1 16751 22678 16751 22678 0 _0030_
rlabel metal2 16698 19618 16698 19618 0 _0031_
rlabel metal2 13846 19618 13846 19618 0 _0032_
rlabel metal2 14766 17476 14766 17476 0 _0033_
rlabel metal2 16790 18054 16790 18054 0 _0034_
rlabel metal1 16647 15402 16647 15402 0 _0035_
rlabel metal1 18062 17238 18062 17238 0 _0036_
rlabel metal2 14766 15810 14766 15810 0 _0037_
rlabel metal1 15538 12206 15538 12206 0 _0038_
rlabel metal1 13370 11798 13370 11798 0 _0039_
rlabel metal1 13493 13974 13493 13974 0 _0040_
rlabel metal1 13892 16218 13892 16218 0 _0041_
rlabel metal1 11576 15062 11576 15062 0 _0042_
rlabel metal1 8310 19414 8310 19414 0 _0043_
rlabel metal2 4830 18530 4830 18530 0 _0044_
rlabel metal1 7452 17850 7452 17850 0 _0045_
rlabel metal1 2852 17850 2852 17850 0 _0046_
rlabel metal2 1978 16966 1978 16966 0 _0047_
rlabel via1 1697 11730 1697 11730 0 _0048_
rlabel metal1 2514 13974 2514 13974 0 _0049_
rlabel metal2 2530 15266 2530 15266 0 _0050_
rlabel metal2 10442 27812 10442 27812 0 _0051_
rlabel metal1 9982 26860 9982 26860 0 _0052_
rlabel metal1 9204 24786 9204 24786 0 _0053_
rlabel metal1 7820 27098 7820 27098 0 _0054_
rlabel metal1 6501 23766 6501 23766 0 _0055_
rlabel metal1 3546 23766 3546 23766 0 _0056_
rlabel metal1 1881 24174 1881 24174 0 _0057_
rlabel via1 1697 27438 1697 27438 0 _0058_
rlabel metal2 2990 27438 2990 27438 0 _0059_
rlabel metal1 8188 21930 8188 21930 0 _0060_
rlabel metal2 6946 25602 6946 25602 0 _0061_
rlabel metal2 8326 24752 8326 24752 0 _0062_
rlabel metal1 7038 26316 7038 26316 0 _0063_
rlabel metal2 7866 21114 7866 21114 0 _0064_
rlabel metal1 5382 20978 5382 20978 0 _0065_
rlabel metal1 18630 20978 18630 20978 0 _0066_
rlabel metal1 20838 23086 20838 23086 0 _0067_
rlabel via1 23414 21522 23414 21522 0 _0068_
rlabel metal2 9982 16796 9982 16796 0 _0069_
rlabel metal1 14674 13940 14674 13940 0 _0070_
rlabel metal2 8694 14620 8694 14620 0 _0071_
rlabel metal1 2162 26010 2162 26010 0 _0072_
rlabel metal1 3358 27642 3358 27642 0 _0073_
rlabel metal1 2162 25908 2162 25908 0 _0074_
rlabel metal2 1794 25466 1794 25466 0 _0075_
rlabel metal1 6348 26010 6348 26010 0 _0076_
rlabel metal1 7452 24786 7452 24786 0 _0077_
rlabel metal1 2369 25262 2369 25262 0 _0078_
rlabel metal2 6394 25534 6394 25534 0 _0079_
rlabel metal1 7682 26554 7682 26554 0 _0080_
rlabel metal2 5382 24956 5382 24956 0 _0081_
rlabel metal1 4462 25772 4462 25772 0 _0082_
rlabel metal1 5382 25262 5382 25262 0 _0083_
rlabel metal1 4416 24582 4416 24582 0 _0084_
rlabel metal1 4600 26554 4600 26554 0 _0085_
rlabel via1 4817 26350 4817 26350 0 _0086_
rlabel metal1 5796 25806 5796 25806 0 _0087_
rlabel metal1 5658 24752 5658 24752 0 _0088_
rlabel metal1 5336 24650 5336 24650 0 _0089_
rlabel metal1 4278 25908 4278 25908 0 _0090_
rlabel metal2 5014 26401 5014 26401 0 _0091_
rlabel metal1 5612 26554 5612 26554 0 _0092_
rlabel metal1 6440 27642 6440 27642 0 _0093_
rlabel metal1 4692 28186 4692 28186 0 _0094_
rlabel metal1 5382 27574 5382 27574 0 _0095_
rlabel metal1 6072 28050 6072 28050 0 _0096_
rlabel metal1 6670 26554 6670 26554 0 _0097_
rlabel metal2 6578 28254 6578 28254 0 _0098_
rlabel metal2 21068 26010 21068 26010 0 _0099_
rlabel metal2 20010 25636 20010 25636 0 _0100_
rlabel metal1 18354 27030 18354 27030 0 _0101_
rlabel metal1 16192 25942 16192 25942 0 _0102_
rlabel metal1 19090 26554 19090 26554 0 _0103_
rlabel metal1 15962 26792 15962 26792 0 _0104_
rlabel metal2 16146 26452 16146 26452 0 _0105_
rlabel metal2 16514 26758 16514 26758 0 _0106_
rlabel metal2 13110 23936 13110 23936 0 _0107_
rlabel metal1 17204 27506 17204 27506 0 _0108_
rlabel metal1 16200 27370 16200 27370 0 _0109_
rlabel metal2 16698 24684 16698 24684 0 _0110_
rlabel metal2 17526 26418 17526 26418 0 _0111_
rlabel metal1 15640 23494 15640 23494 0 _0112_
rlabel metal1 14582 25908 14582 25908 0 _0113_
rlabel via1 15494 23834 15494 23834 0 _0114_
rlabel metal1 14858 23732 14858 23732 0 _0115_
rlabel metal2 14122 26115 14122 26115 0 _0116_
rlabel metal1 13424 27030 13424 27030 0 _0117_
rlabel metal2 13754 26112 13754 26112 0 _0118_
rlabel metal2 13478 24956 13478 24956 0 _0119_
rlabel metal1 13570 27540 13570 27540 0 _0120_
rlabel metal1 12834 24106 12834 24106 0 _0121_
rlabel metal1 12834 25772 12834 25772 0 _0122_
rlabel metal1 12972 26486 12972 26486 0 _0123_
rlabel metal1 6900 22746 6900 22746 0 _0124_
rlabel metal1 8970 20876 8970 20876 0 _0125_
rlabel metal2 11822 15742 11822 15742 0 _0126_
rlabel metal2 8510 16983 8510 16983 0 _0127_
rlabel metal2 11638 18292 11638 18292 0 _0128_
rlabel metal1 10166 18700 10166 18700 0 _0129_
rlabel metal1 10534 17850 10534 17850 0 _0130_
rlabel via1 6486 19346 6486 19346 0 _0131_
rlabel metal1 12466 22168 12466 22168 0 _0132_
rlabel metal1 13570 20434 13570 20434 0 _0133_
rlabel metal2 5290 15334 5290 15334 0 _0134_
rlabel metal1 4876 17306 4876 17306 0 _0135_
rlabel metal1 10074 18700 10074 18700 0 _0136_
rlabel metal2 12650 18190 12650 18190 0 _0137_
rlabel metal1 10442 17612 10442 17612 0 _0138_
rlabel metal1 10534 17782 10534 17782 0 _0139_
rlabel metal1 11684 17306 11684 17306 0 _0140_
rlabel metal1 10762 18734 10762 18734 0 _0141_
rlabel metal1 12466 16626 12466 16626 0 _0142_
rlabel metal1 11546 16456 11546 16456 0 _0143_
rlabel metal2 11086 17680 11086 17680 0 _0144_
rlabel metal1 11546 18836 11546 18836 0 _0145_
rlabel metal1 11178 18734 11178 18734 0 _0146_
rlabel metal2 10442 19074 10442 19074 0 _0147_
rlabel metal1 10258 19822 10258 19822 0 _0148_
rlabel metal1 9476 18734 9476 18734 0 _0149_
rlabel metal1 5796 21114 5796 21114 0 _0150_
rlabel metal2 6762 21454 6762 21454 0 _0151_
rlabel metal1 7130 20910 7130 20910 0 _0152_
rlabel metal2 7222 21828 7222 21828 0 _0153_
rlabel metal1 5658 20944 5658 20944 0 _0154_
rlabel metal1 6348 19346 6348 19346 0 _0155_
rlabel metal2 6578 20196 6578 20196 0 _0156_
rlabel via1 6856 19346 6856 19346 0 _0157_
rlabel metal2 5658 19788 5658 19788 0 _0158_
rlabel metal1 6808 21590 6808 21590 0 _0159_
rlabel metal1 6532 19210 6532 19210 0 _0160_
rlabel metal1 6210 21454 6210 21454 0 _0161_
rlabel metal2 9614 17238 9614 17238 0 _0162_
rlabel metal1 13202 22134 13202 22134 0 _0163_
rlabel metal2 13202 20604 13202 20604 0 _0164_
rlabel metal1 13524 17850 13524 17850 0 _0165_
rlabel metal2 13018 18020 13018 18020 0 _0166_
rlabel metal1 10594 17646 10594 17646 0 _0167_
rlabel metal1 8326 17238 8326 17238 0 _0168_
rlabel metal1 9890 17714 9890 17714 0 _0169_
rlabel metal1 9844 17850 9844 17850 0 _0170_
rlabel metal1 5106 17136 5106 17136 0 _0171_
rlabel via1 4738 16082 4738 16082 0 _0172_
rlabel metal1 12558 22644 12558 22644 0 _0173_
rlabel metal1 16514 14382 16514 14382 0 _0174_
rlabel metal2 9062 20570 9062 20570 0 _0175_
rlabel metal1 9936 21998 9936 21998 0 _0176_
rlabel metal2 9246 22712 9246 22712 0 _0177_
rlabel metal2 10442 24106 10442 24106 0 _0178_
rlabel metal1 11178 23732 11178 23732 0 _0179_
rlabel metal1 11454 21964 11454 21964 0 _0180_
rlabel metal1 12604 23086 12604 23086 0 _0181_
rlabel metal1 11730 21522 11730 21522 0 _0182_
rlabel metal2 12834 23732 12834 23732 0 _0183_
rlabel metal1 12972 23290 12972 23290 0 _0184_
rlabel metal1 5290 16116 5290 16116 0 _0185_
rlabel metal2 5474 16796 5474 16796 0 _0186_
rlabel metal2 4278 16252 4278 16252 0 _0187_
rlabel metal1 5980 16082 5980 16082 0 _0188_
rlabel metal1 10161 16048 10161 16048 0 _0189_
rlabel metal1 15226 14348 15226 14348 0 _0190_
rlabel metal2 8142 17238 8142 17238 0 _0191_
rlabel metal1 7268 16558 7268 16558 0 _0192_
rlabel metal1 4600 12682 4600 12682 0 _0193_
rlabel metal1 10626 14416 10626 14416 0 _0194_
rlabel metal1 12466 12172 12466 12172 0 _0195_
rlabel metal1 10166 13702 10166 13702 0 _0196_
rlabel metal1 9982 14994 9982 14994 0 _0197_
rlabel metal2 10442 13532 10442 13532 0 _0198_
rlabel metal2 8970 14076 8970 14076 0 _0199_
rlabel metal2 9154 13498 9154 13498 0 _0200_
rlabel metal1 9246 10710 9246 10710 0 _0201_
rlabel metal2 10166 12988 10166 12988 0 _0202_
rlabel metal1 9614 12206 9614 12206 0 _0203_
rlabel metal1 8694 12308 8694 12308 0 _0204_
rlabel metal1 8786 12274 8786 12274 0 _0205_
rlabel metal2 8234 10778 8234 10778 0 _0206_
rlabel metal1 8740 16082 8740 16082 0 _0207_
rlabel metal1 7958 15674 7958 15674 0 _0208_
rlabel metal1 8188 13430 8188 13430 0 _0209_
rlabel metal1 8510 12240 8510 12240 0 _0210_
rlabel metal2 8418 14212 8418 14212 0 _0211_
rlabel metal1 7038 12410 7038 12410 0 _0212_
rlabel metal1 6992 11662 6992 11662 0 _0213_
rlabel metal1 8096 12818 8096 12818 0 _0214_
rlabel metal2 7222 15436 7222 15436 0 _0215_
rlabel metal1 7222 14450 7222 14450 0 _0216_
rlabel metal1 6624 11730 6624 11730 0 _0217_
rlabel metal1 8326 15504 8326 15504 0 _0218_
rlabel metal1 8694 15130 8694 15130 0 _0219_
rlabel metal1 8510 13498 8510 13498 0 _0220_
rlabel metal1 8050 13498 8050 13498 0 _0221_
rlabel metal2 7590 7055 7590 7055 0 _0222_
rlabel metal2 7590 11696 7590 11696 0 _0223_
rlabel metal2 8142 12886 8142 12886 0 _0224_
rlabel metal1 5566 11764 5566 11764 0 _0225_
rlabel metal1 8418 12716 8418 12716 0 _0226_
rlabel metal1 10902 12886 10902 12886 0 _0227_
rlabel metal1 10672 9010 10672 9010 0 _0228_
rlabel metal2 10718 12988 10718 12988 0 _0229_
rlabel metal1 10764 11118 10764 11118 0 _0230_
rlabel metal1 9154 12818 9154 12818 0 _0231_
rlabel metal1 6118 11730 6118 11730 0 _0232_
rlabel metal1 5474 11050 5474 11050 0 _0233_
rlabel metal1 6210 16558 6210 16558 0 _0234_
rlabel metal1 4462 14484 4462 14484 0 _0235_
rlabel metal2 3266 11866 3266 11866 0 _0236_
rlabel metal2 3542 10030 3542 10030 0 _0237_
rlabel metal2 4094 14620 4094 14620 0 _0238_
rlabel metal1 3864 14246 3864 14246 0 _0239_
rlabel metal1 5290 11764 5290 11764 0 _0240_
rlabel metal2 6210 15708 6210 15708 0 _0241_
rlabel metal2 6394 14416 6394 14416 0 _0242_
rlabel metal1 5473 13328 5473 13328 0 _0243_
rlabel metal1 5244 13158 5244 13158 0 _0244_
rlabel metal1 4094 12614 4094 12614 0 _0245_
rlabel metal1 4738 13702 4738 13702 0 _0246_
rlabel metal1 5566 14042 5566 14042 0 _0247_
rlabel metal1 5704 7310 5704 7310 0 _0248_
rlabel metal1 6302 16456 6302 16456 0 _0249_
rlabel metal2 4830 14110 4830 14110 0 _0250_
rlabel metal1 4876 14042 4876 14042 0 _0251_
rlabel metal2 4830 11492 4830 11492 0 _0252_
rlabel metal1 10120 11118 10120 11118 0 _0253_
rlabel metal1 4508 12206 4508 12206 0 _0254_
rlabel metal1 5106 10030 5106 10030 0 _0255_
rlabel metal2 9522 10336 9522 10336 0 _0256_
rlabel metal2 5566 9146 5566 9146 0 _0257_
rlabel metal1 12650 12240 12650 12240 0 _0258_
rlabel metal2 12650 11900 12650 11900 0 _0259_
rlabel metal2 12466 11900 12466 11900 0 _0260_
rlabel metal2 12650 11084 12650 11084 0 _0261_
rlabel metal1 13018 9588 13018 9588 0 _0262_
rlabel metal2 12742 10812 12742 10812 0 _0263_
rlabel metal1 8050 9996 8050 9996 0 _0264_
rlabel metal1 8004 9894 8004 9894 0 _0265_
rlabel metal2 6670 9758 6670 9758 0 _0266_
rlabel metal2 6302 10404 6302 10404 0 _0267_
rlabel metal2 6946 12240 6946 12240 0 _0268_
rlabel metal1 6670 7310 6670 7310 0 _0269_
rlabel metal1 6302 7514 6302 7514 0 _0270_
rlabel metal1 7958 7412 7958 7412 0 _0271_
rlabel metal2 6578 9180 6578 9180 0 _0272_
rlabel metal1 7636 7378 7636 7378 0 _0273_
rlabel metal1 7406 7412 7406 7412 0 _0274_
rlabel metal1 7774 9452 7774 9452 0 _0275_
rlabel metal2 7774 7548 7774 7548 0 _0276_
rlabel metal1 8004 6426 8004 6426 0 _0277_
rlabel metal2 7958 5474 7958 5474 0 _0278_
rlabel metal2 9338 10370 9338 10370 0 _0279_
rlabel metal1 10120 8262 10120 8262 0 _0280_
rlabel metal2 10718 6970 10718 6970 0 _0281_
rlabel metal1 10718 11220 10718 11220 0 _0282_
rlabel metal1 9982 8983 9982 8983 0 _0283_
rlabel metal2 11270 8670 11270 8670 0 _0284_
rlabel metal2 9798 8058 9798 8058 0 _0285_
rlabel metal2 9154 10812 9154 10812 0 _0286_
rlabel metal2 9890 9146 9890 9146 0 _0287_
rlabel metal2 8602 8670 8602 8670 0 _0288_
rlabel metal1 8924 5134 8924 5134 0 _0289_
rlabel metal1 8096 7786 8096 7786 0 _0290_
rlabel metal1 9062 7446 9062 7446 0 _0291_
rlabel metal1 6394 7412 6394 7412 0 _0292_
rlabel metal1 11316 11322 11316 11322 0 _0293_
rlabel metal1 11500 8942 11500 8942 0 _0294_
rlabel metal1 9154 7888 9154 7888 0 _0295_
rlabel metal2 8694 7548 8694 7548 0 _0296_
rlabel metal2 6578 7548 6578 7548 0 _0297_
rlabel metal1 6486 6800 6486 6800 0 _0298_
rlabel metal1 6578 6630 6578 6630 0 _0299_
rlabel metal2 5014 9282 5014 9282 0 _0300_
rlabel metal1 5612 9010 5612 9010 0 _0301_
rlabel metal2 5934 7242 5934 7242 0 _0302_
rlabel metal1 5842 13947 5842 13947 0 _0303_
rlabel metal1 5980 5338 5980 5338 0 _0304_
rlabel metal1 6348 5542 6348 5542 0 _0305_
rlabel metal1 4738 7820 4738 7820 0 _0306_
rlabel metal1 4646 9554 4646 9554 0 _0307_
rlabel metal1 4462 10540 4462 10540 0 _0308_
rlabel metal2 4462 7548 4462 7548 0 _0309_
rlabel metal1 4002 8976 4002 8976 0 _0310_
rlabel metal2 3818 9146 3818 9146 0 _0311_
rlabel metal2 4646 5984 4646 5984 0 _0312_
rlabel metal1 4738 7922 4738 7922 0 _0313_
rlabel metal1 4370 7956 4370 7956 0 _0314_
rlabel metal2 12466 9316 12466 9316 0 _0315_
rlabel metal1 4055 10642 4055 10642 0 _0316_
rlabel metal1 4738 7412 4738 7412 0 _0317_
rlabel metal1 9430 8534 9430 8534 0 _0318_
rlabel metal1 13064 10506 13064 10506 0 _0319_
rlabel metal2 11822 9962 11822 9962 0 _0320_
rlabel metal1 14122 10030 14122 10030 0 _0321_
rlabel metal2 12834 9350 12834 9350 0 _0322_
rlabel metal1 14812 9486 14812 9486 0 _0323_
rlabel metal1 14030 8432 14030 8432 0 _0324_
rlabel metal1 13938 7922 13938 7922 0 _0325_
rlabel metal2 5290 8058 5290 8058 0 _0326_
rlabel via2 12558 7803 12558 7803 0 _0327_
rlabel metal1 4646 5270 4646 5270 0 _0328_
rlabel metal2 5474 4794 5474 4794 0 _0329_
rlabel metal1 10074 4080 10074 4080 0 _0330_
rlabel metal1 6210 6154 6210 6154 0 _0331_
rlabel metal1 6348 5202 6348 5202 0 _0332_
rlabel metal2 10534 4964 10534 4964 0 _0333_
rlabel metal1 5106 4590 5106 4590 0 _0334_
rlabel viali 13662 3502 13662 3502 0 _0335_
rlabel metal2 11178 4284 11178 4284 0 _0336_
rlabel metal2 11270 7854 11270 7854 0 _0337_
rlabel metal1 10856 6766 10856 6766 0 _0338_
rlabel metal2 10442 6426 10442 6426 0 _0339_
rlabel metal1 9660 5746 9660 5746 0 _0340_
rlabel metal1 11040 5678 11040 5678 0 _0341_
rlabel metal1 14490 5270 14490 5270 0 _0342_
rlabel metal1 11408 9078 11408 9078 0 _0343_
rlabel metal2 13294 6766 13294 6766 0 _0344_
rlabel metal2 12098 8398 12098 8398 0 _0345_
rlabel metal1 13156 6290 13156 6290 0 _0346_
rlabel metal2 13662 9214 13662 9214 0 _0347_
rlabel metal1 13708 5678 13708 5678 0 _0348_
rlabel metal1 11500 7310 11500 7310 0 _0349_
rlabel metal2 12742 6562 12742 6562 0 _0350_
rlabel metal1 12742 6154 12742 6154 0 _0351_
rlabel metal1 8786 4556 8786 4556 0 _0352_
rlabel metal1 8878 4658 8878 4658 0 _0353_
rlabel metal1 12489 4590 12489 4590 0 _0354_
rlabel metal2 8878 6970 8878 6970 0 _0355_
rlabel metal1 13386 4692 13386 4692 0 _0356_
rlabel metal1 11638 5882 11638 5882 0 _0357_
rlabel metal2 12650 6086 12650 6086 0 _0358_
rlabel metal2 11914 5440 11914 5440 0 _0359_
rlabel metal1 12374 6154 12374 6154 0 _0360_
rlabel metal2 12926 5644 12926 5644 0 _0361_
rlabel metal1 11822 2278 11822 2278 0 _0362_
rlabel metal1 10626 2482 10626 2482 0 _0363_
rlabel metal1 9798 4182 9798 4182 0 _0364_
rlabel metal1 6302 6290 6302 6290 0 _0365_
rlabel metal2 9982 5134 9982 5134 0 _0366_
rlabel metal2 10534 3502 10534 3502 0 _0367_
rlabel metal1 10672 4046 10672 4046 0 _0368_
rlabel metal2 13478 3553 13478 3553 0 _0369_
rlabel metal1 11638 4250 11638 4250 0 _0370_
rlabel metal2 12834 4352 12834 4352 0 _0371_
rlabel viali 15044 7854 15044 7854 0 _0372_
rlabel metal2 14306 8466 14306 8466 0 _0373_
rlabel metal1 14030 8942 14030 8942 0 _0374_
rlabel metal1 14950 8874 14950 8874 0 _0375_
rlabel metal1 14122 3536 14122 3536 0 _0376_
rlabel metal1 12650 2992 12650 2992 0 _0377_
rlabel metal1 13018 3094 13018 3094 0 _0378_
rlabel metal1 13662 2380 13662 2380 0 _0379_
rlabel metal1 10626 2992 10626 2992 0 _0380_
rlabel metal1 10442 3128 10442 3128 0 _0381_
rlabel metal1 16422 2822 16422 2822 0 _0382_
rlabel metal2 13570 3434 13570 3434 0 _0383_
rlabel metal1 15732 3502 15732 3502 0 _0384_
rlabel metal1 15548 3638 15548 3638 0 _0385_
rlabel metal1 13386 6256 13386 6256 0 _0386_
rlabel metal1 14674 6154 14674 6154 0 _0387_
rlabel metal2 14858 6154 14858 6154 0 _0388_
rlabel metal1 13754 5134 13754 5134 0 _0389_
rlabel metal1 15870 6324 15870 6324 0 _0390_
rlabel metal1 14352 7514 14352 7514 0 _0391_
rlabel metal1 17158 11186 17158 11186 0 _0392_
rlabel metal2 15502 10744 15502 10744 0 _0393_
rlabel metal2 15594 9554 15594 9554 0 _0394_
rlabel metal2 16054 9282 16054 9282 0 _0395_
rlabel metal2 16790 10404 16790 10404 0 _0396_
rlabel metal1 16330 9146 16330 9146 0 _0397_
rlabel metal1 15410 9962 15410 9962 0 _0398_
rlabel via1 16246 8874 16246 8874 0 _0399_
rlabel metal1 17986 8908 17986 8908 0 _0400_
rlabel metal1 14996 7378 14996 7378 0 _0401_
rlabel metal1 14628 7854 14628 7854 0 _0402_
rlabel metal2 17158 8228 17158 8228 0 _0403_
rlabel metal1 17986 7854 17986 7854 0 _0404_
rlabel metal2 16330 7548 16330 7548 0 _0405_
rlabel metal2 15962 6596 15962 6596 0 _0406_
rlabel metal1 17526 7344 17526 7344 0 _0407_
rlabel metal1 16422 6732 16422 6732 0 _0408_
rlabel metal1 17250 6732 17250 6732 0 _0409_
rlabel metal2 16698 5372 16698 5372 0 _0410_
rlabel metal2 15594 5338 15594 5338 0 _0411_
rlabel metal1 13202 4556 13202 4556 0 _0412_
rlabel metal1 12834 4658 12834 4658 0 _0413_
rlabel metal1 16054 4590 16054 4590 0 _0414_
rlabel metal1 14904 5134 14904 5134 0 _0415_
rlabel metal1 16514 5236 16514 5236 0 _0416_
rlabel metal2 16330 4998 16330 4998 0 _0417_
rlabel metal1 16790 5168 16790 5168 0 _0418_
rlabel metal1 15686 4624 15686 4624 0 _0419_
rlabel metal2 16238 3774 16238 3774 0 _0420_
rlabel metal2 15870 2587 15870 2587 0 _0421_
rlabel metal2 9522 3978 9522 3978 0 _0422_
rlabel metal1 15318 2550 15318 2550 0 _0423_
rlabel metal1 15686 3094 15686 3094 0 _0424_
rlabel metal1 16882 3502 16882 3502 0 _0425_
rlabel metal1 14582 3638 14582 3638 0 _0426_
rlabel metal2 17940 8942 17940 8942 0 _0427_
rlabel metal1 17342 2414 17342 2414 0 _0428_
rlabel metal1 17204 5678 17204 5678 0 _0429_
rlabel metal2 17342 10268 17342 10268 0 _0430_
rlabel metal2 16882 9180 16882 9180 0 _0431_
rlabel metal1 20056 8942 20056 8942 0 _0432_
rlabel metal1 17848 2414 17848 2414 0 _0433_
rlabel metal1 18308 2618 18308 2618 0 _0434_
rlabel metal2 20102 3332 20102 3332 0 _0435_
rlabel metal1 21298 3060 21298 3060 0 _0436_
rlabel metal1 17986 3570 17986 3570 0 _0437_
rlabel metal1 17940 2958 17940 2958 0 _0438_
rlabel metal1 20838 2958 20838 2958 0 _0439_
rlabel metal1 17940 5338 17940 5338 0 _0440_
rlabel metal1 18308 4658 18308 4658 0 _0441_
rlabel metal2 19826 4998 19826 4998 0 _0442_
rlabel metal1 22264 5202 22264 5202 0 _0443_
rlabel metal1 15272 2414 15272 2414 0 _0444_
rlabel metal1 16008 2618 16008 2618 0 _0445_
rlabel metal2 20010 4607 20010 4607 0 _0446_
rlabel metal1 19826 5644 19826 5644 0 _0447_
rlabel metal1 17480 5542 17480 5542 0 _0448_
rlabel metal1 18400 5610 18400 5610 0 _0449_
rlabel via1 19826 6630 19826 6630 0 _0450_
rlabel metal2 18722 6528 18722 6528 0 _0451_
rlabel metal1 20470 5746 20470 5746 0 _0452_
rlabel metal2 18078 7514 18078 7514 0 _0453_
rlabel metal2 17066 6970 17066 6970 0 _0454_
rlabel metal1 19642 7888 19642 7888 0 _0455_
rlabel metal1 18124 8466 18124 8466 0 _0456_
rlabel metal1 21850 8432 21850 8432 0 _0457_
rlabel metal1 20424 8466 20424 8466 0 _0458_
rlabel metal1 20194 6834 20194 6834 0 _0459_
rlabel metal1 21574 5610 21574 5610 0 _0460_
rlabel metal2 20378 6154 20378 6154 0 _0461_
rlabel metal2 20286 5168 20286 5168 0 _0462_
rlabel metal1 17802 10166 17802 10166 0 _0463_
rlabel metal1 16974 10234 16974 10234 0 _0464_
rlabel metal2 19734 10370 19734 10370 0 _0465_
rlabel metal1 18032 11118 18032 11118 0 _0466_
rlabel metal1 20746 10642 20746 10642 0 _0467_
rlabel metal2 18630 11254 18630 11254 0 _0468_
rlabel metal1 20056 16762 20056 16762 0 _0469_
rlabel metal1 19734 10642 19734 10642 0 _0470_
rlabel metal2 20010 10268 20010 10268 0 _0471_
rlabel metal2 22310 10506 22310 10506 0 _0472_
rlabel metal2 19550 9996 19550 9996 0 _0473_
rlabel metal2 19550 9112 19550 9112 0 _0474_
rlabel metal2 22034 8704 22034 8704 0 _0475_
rlabel metal2 20562 6562 20562 6562 0 _0476_
rlabel metal2 20470 5168 20470 5168 0 _0477_
rlabel metal2 20654 4012 20654 4012 0 _0478_
rlabel metal2 21298 3570 21298 3570 0 _0479_
rlabel metal1 17779 3366 17779 3366 0 _0480_
rlabel viali 20838 3503 20838 3503 0 _0481_
rlabel metal1 21390 3400 21390 3400 0 _0482_
rlabel metal1 21850 16558 21850 16558 0 _0483_
rlabel metal1 19964 9146 19964 9146 0 _0484_
rlabel metal1 20194 16490 20194 16490 0 _0485_
rlabel via1 19742 8806 19742 8806 0 _0486_
rlabel metal1 21850 7310 21850 7310 0 _0487_
rlabel metal1 22862 8976 22862 8976 0 _0488_
rlabel metal1 19918 9044 19918 9044 0 _0489_
rlabel metal1 22356 15470 22356 15470 0 _0490_
rlabel metal2 21850 10404 21850 10404 0 _0491_
rlabel metal1 22035 10098 22035 10098 0 _0492_
rlabel metal1 24426 15470 24426 15470 0 _0493_
rlabel metal1 20884 10778 20884 10778 0 _0494_
rlabel metal2 21206 10268 21206 10268 0 _0495_
rlabel metal1 23506 14994 23506 14994 0 _0496_
rlabel metal1 20838 17136 20838 17136 0 _0497_
rlabel metal1 21252 16694 21252 16694 0 _0498_
rlabel metal2 22402 17714 22402 17714 0 _0499_
rlabel metal2 21206 16898 21206 16898 0 _0500_
rlabel metal1 20470 17204 20470 17204 0 _0501_
rlabel metal1 21022 17306 21022 17306 0 _0502_
rlabel metal1 21597 17034 21597 17034 0 _0503_
rlabel metal1 23046 14518 23046 14518 0 _0504_
rlabel metal1 21850 10506 21850 10506 0 _0505_
rlabel metal1 24426 14416 24426 14416 0 _0506_
rlabel metal1 24012 15130 24012 15130 0 _0507_
rlabel metal2 22586 10438 22586 10438 0 _0508_
rlabel metal1 24518 10676 24518 10676 0 _0509_
rlabel metal2 20746 7514 20746 7514 0 _0510_
rlabel metal2 21022 6562 21022 6562 0 _0511_
rlabel metal1 19964 6086 19964 6086 0 _0512_
rlabel metal1 21850 6834 21850 6834 0 _0513_
rlabel metal2 18446 6086 18446 6086 0 _0514_
rlabel metal1 21206 6290 21206 6290 0 _0515_
rlabel metal1 21942 5712 21942 5712 0 _0516_
rlabel metal2 23230 6086 23230 6086 0 _0517_
rlabel metal1 25254 7378 25254 7378 0 _0518_
rlabel metal1 25438 6800 25438 6800 0 _0519_
rlabel metal1 22678 5678 22678 5678 0 _0520_
rlabel metal2 23230 5338 23230 5338 0 _0521_
rlabel metal2 23506 6222 23506 6222 0 _0522_
rlabel metal1 23644 6426 23644 6426 0 _0523_
rlabel metal1 25622 6426 25622 6426 0 _0524_
rlabel metal2 24702 9792 24702 9792 0 _0525_
rlabel metal1 22494 8602 22494 8602 0 _0526_
rlabel metal1 22770 7446 22770 7446 0 _0527_
rlabel metal2 24150 8092 24150 8092 0 _0528_
rlabel metal1 23598 7854 23598 7854 0 _0529_
rlabel metal1 20654 12138 20654 12138 0 _0530_
rlabel metal1 21160 6970 21160 6970 0 _0531_
rlabel metal1 21666 7208 21666 7208 0 _0532_
rlabel metal2 24058 9724 24058 9724 0 _0533_
rlabel metal1 23368 6766 23368 6766 0 _0534_
rlabel metal2 23690 5338 23690 5338 0 _0535_
rlabel metal1 23414 8058 23414 8058 0 _0536_
rlabel metal2 24334 7582 24334 7582 0 _0537_
rlabel metal2 24058 5508 24058 5508 0 _0538_
rlabel metal2 23506 4828 23506 4828 0 _0539_
rlabel metal1 24610 4080 24610 4080 0 _0540_
rlabel metal1 23138 3162 23138 3162 0 _0541_
rlabel metal1 22540 4046 22540 4046 0 _0542_
rlabel metal2 22402 3808 22402 3808 0 _0543_
rlabel metal2 24702 4352 24702 4352 0 _0544_
rlabel metal1 23552 3638 23552 3638 0 _0545_
rlabel metal1 23874 3536 23874 3536 0 _0546_
rlabel metal3 25461 15300 25461 15300 0 _0547_
rlabel metal1 23368 3706 23368 3706 0 _0548_
rlabel metal1 23452 17238 23452 17238 0 _0549_
rlabel metal1 24472 11322 24472 11322 0 _0550_
rlabel metal1 25116 4658 25116 4658 0 _0551_
rlabel metal1 23920 9554 23920 9554 0 _0552_
rlabel metal1 25300 6766 25300 6766 0 _0553_
rlabel metal2 24886 5372 24886 5372 0 _0554_
rlabel metal2 26174 13362 26174 13362 0 _0555_
rlabel metal1 25898 7276 25898 7276 0 _0556_
rlabel metal1 25300 6698 25300 6698 0 _0557_
rlabel metal1 26082 13260 26082 13260 0 _0558_
rlabel metal1 26450 12886 26450 12886 0 _0559_
rlabel metal1 25024 13226 25024 13226 0 _0560_
rlabel metal2 23046 12002 23046 12002 0 _0561_
rlabel metal1 23552 9690 23552 9690 0 _0562_
rlabel metal1 25070 12852 25070 12852 0 _0563_
rlabel metal1 24748 12750 24748 12750 0 _0564_
rlabel metal2 25162 8602 25162 8602 0 _0565_
rlabel metal1 24058 8330 24058 8330 0 _0566_
rlabel metal2 23230 12036 23230 12036 0 _0567_
rlabel metal2 22034 14654 22034 14654 0 _0568_
rlabel metal1 26082 11220 26082 11220 0 _0569_
rlabel metal1 23138 15395 23138 15395 0 _0570_
rlabel metal1 24610 10574 24610 10574 0 _0571_
rlabel metal2 25070 14722 25070 14722 0 _0572_
rlabel via1 24703 14994 24703 14994 0 _0573_
rlabel metal2 25530 15878 25530 15878 0 _0574_
rlabel metal1 25346 16116 25346 16116 0 _0575_
rlabel metal1 25070 16048 25070 16048 0 _0576_
rlabel metal2 24518 14858 24518 14858 0 _0577_
rlabel metal2 24886 15606 24886 15606 0 _0578_
rlabel metal2 22862 18462 22862 18462 0 _0579_
rlabel metal1 22678 17612 22678 17612 0 _0580_
rlabel metal2 22862 19924 22862 19924 0 _0581_
rlabel metal1 22954 19380 22954 19380 0 _0582_
rlabel metal2 21850 17782 21850 17782 0 _0583_
rlabel metal1 23414 16626 23414 16626 0 _0584_
rlabel metal2 23138 19040 23138 19040 0 _0585_
rlabel metal1 23292 19414 23292 19414 0 _0586_
rlabel metal1 24334 19380 24334 19380 0 _0587_
rlabel metal1 24150 19482 24150 19482 0 _0588_
rlabel metal2 24058 19686 24058 19686 0 _0589_
rlabel metal2 24610 17952 24610 17952 0 _0590_
rlabel metal1 25254 17000 25254 17000 0 _0591_
rlabel metal1 25300 15878 25300 15878 0 _0592_
rlabel metal1 24058 13974 24058 13974 0 _0593_
rlabel metal1 25760 12818 25760 12818 0 _0594_
rlabel metal1 26174 13362 26174 13362 0 _0595_
rlabel metal1 26634 11730 26634 11730 0 _0596_
rlabel metal1 26128 11322 26128 11322 0 _0597_
rlabel metal1 26358 11628 26358 11628 0 _0598_
rlabel metal1 26588 10030 26588 10030 0 _0599_
rlabel metal2 25530 7378 25530 7378 0 _0600_
rlabel metal1 24932 3570 24932 3570 0 _0601_
rlabel metal1 25760 10030 25760 10030 0 _0602_
rlabel metal1 25990 17170 25990 17170 0 _0603_
rlabel metal1 26404 10030 26404 10030 0 _0604_
rlabel metal2 21298 13566 21298 13566 0 _0605_
rlabel metal1 26680 14042 26680 14042 0 _0606_
rlabel metal1 20148 13906 20148 13906 0 _0607_
rlabel metal1 19772 13896 19772 13896 0 _0608_
rlabel metal1 24104 12818 24104 12818 0 _0609_
rlabel metal1 19688 13294 19688 13294 0 _0610_
rlabel metal1 24012 12886 24012 12886 0 _0611_
rlabel metal1 21758 13328 21758 13328 0 _0612_
rlabel metal1 24932 18258 24932 18258 0 _0613_
rlabel metal2 25622 17612 25622 17612 0 _0614_
rlabel metal1 19182 18190 19182 18190 0 _0615_
rlabel metal2 25070 18020 25070 18020 0 _0616_
rlabel metal1 24426 18292 24426 18292 0 _0617_
rlabel metal1 20470 18360 20470 18360 0 _0618_
rlabel metal1 21298 19822 21298 19822 0 _0619_
rlabel metal2 24242 20196 24242 20196 0 _0620_
rlabel metal2 24426 20060 24426 20060 0 _0621_
rlabel metal2 21666 19584 21666 19584 0 _0622_
rlabel metal1 22954 19958 22954 19958 0 _0623_
rlabel metal1 23230 13158 23230 13158 0 _0624_
rlabel metal2 22310 14076 22310 14076 0 _0625_
rlabel metal2 22586 14212 22586 14212 0 _0626_
rlabel metal2 21206 15198 21206 15198 0 _0627_
rlabel metal1 26220 15538 26220 15538 0 _0628_
rlabel metal1 20930 14790 20930 14790 0 _0629_
rlabel metal2 21206 14076 21206 14076 0 _0630_
rlabel metal1 20562 12308 20562 12308 0 _0631_
rlabel metal1 21114 13226 21114 13226 0 _0632_
rlabel metal1 20424 13498 20424 13498 0 _0633_
rlabel metal1 22540 21046 22540 21046 0 _0634_
rlabel metal2 22402 20264 22402 20264 0 _0635_
rlabel metal1 22402 20842 22402 20842 0 _0636_
rlabel metal2 22678 21318 22678 21318 0 _0637_
rlabel metal1 22310 21522 22310 21522 0 _0638_
rlabel metal1 21206 20944 21206 20944 0 _0639_
rlabel metal1 20516 20502 20516 20502 0 _0640_
rlabel metal1 20792 20910 20792 20910 0 _0641_
rlabel metal1 20470 19788 20470 19788 0 _0642_
rlabel metal1 20286 20978 20286 20978 0 _0643_
rlabel metal2 20102 19584 20102 19584 0 _0644_
rlabel metal2 21574 17578 21574 17578 0 _0645_
rlabel metal2 21482 18972 21482 18972 0 _0646_
rlabel metal2 21482 17034 21482 17034 0 _0647_
rlabel metal2 20286 18768 20286 18768 0 _0648_
rlabel metal2 18722 18972 18722 18972 0 _0649_
rlabel metal1 20930 15504 20930 15504 0 _0650_
rlabel metal1 19182 12852 19182 12852 0 _0651_
rlabel viali 17994 12750 17994 12750 0 _0652_
rlabel metal1 20470 13226 20470 13226 0 _0653_
rlabel metal1 20562 13362 20562 13362 0 _0654_
rlabel metal1 19090 13940 19090 13940 0 _0655_
rlabel metal1 25668 13498 25668 13498 0 _0656_
rlabel metal1 20750 13906 20750 13906 0 _0657_
rlabel metal2 19504 13940 19504 13940 0 _0658_
rlabel metal1 19872 13362 19872 13362 0 _0659_
rlabel metal1 20608 12614 20608 12614 0 _0660_
rlabel metal1 21758 15402 21758 15402 0 _0661_
rlabel metal1 18860 18258 18860 18258 0 _0662_
rlabel metal1 13110 19278 13110 19278 0 _0663_
rlabel metal1 11868 19482 11868 19482 0 _0664_
rlabel metal2 18722 21318 18722 21318 0 _0665_
rlabel metal2 20838 22304 20838 22304 0 _0666_
rlabel metal1 17848 21522 17848 21522 0 _0667_
rlabel metal1 18584 21114 18584 21114 0 _0668_
rlabel metal1 18400 21454 18400 21454 0 _0669_
rlabel metal2 18446 21828 18446 21828 0 _0670_
rlabel metal2 22126 21318 22126 21318 0 _0671_
rlabel metal1 21850 22576 21850 22576 0 _0672_
rlabel metal2 21298 22848 21298 22848 0 _0673_
rlabel metal1 20194 22610 20194 22610 0 _0674_
rlabel metal1 21850 21624 21850 21624 0 _0675_
rlabel metal2 17618 21284 17618 21284 0 _0676_
rlabel metal1 17158 21590 17158 21590 0 _0677_
rlabel metal1 15624 19754 15624 19754 0 _0678_
rlabel metal1 16468 21522 16468 21522 0 _0679_
rlabel metal1 16882 21454 16882 21454 0 _0680_
rlabel metal2 16698 21828 16698 21828 0 _0681_
rlabel metal2 20562 20604 20562 20604 0 _0682_
rlabel metal1 15617 21522 15617 21522 0 _0683_
rlabel metal1 15824 21318 15824 21318 0 _0684_
rlabel metal1 17250 20842 17250 20842 0 _0685_
rlabel metal2 15870 22134 15870 22134 0 _0686_
rlabel metal1 19872 19890 19872 19890 0 _0687_
rlabel metal2 18722 19618 18722 19618 0 _0688_
rlabel metal1 17802 19414 17802 19414 0 _0689_
rlabel metal1 15778 19482 15778 19482 0 _0690_
rlabel metal2 15410 19006 15410 19006 0 _0691_
rlabel metal2 16882 19516 16882 19516 0 _0692_
rlabel metal1 20240 18054 20240 18054 0 _0693_
rlabel metal2 20102 18054 20102 18054 0 _0694_
rlabel metal2 19550 18938 19550 18938 0 _0695_
rlabel metal1 15134 19380 15134 19380 0 _0696_
rlabel metal1 14996 19346 14996 19346 0 _0697_
rlabel metal1 14030 19312 14030 19312 0 _0698_
rlabel metal2 19090 18462 19090 18462 0 _0699_
rlabel metal1 15042 17136 15042 17136 0 _0700_
rlabel metal2 15778 17884 15778 17884 0 _0701_
rlabel metal1 15778 16966 15778 16966 0 _0702_
rlabel metal1 14950 17204 14950 17204 0 _0703_
rlabel metal2 18446 18292 18446 18292 0 _0704_
rlabel metal1 18262 18700 18262 18700 0 _0705_
rlabel metal2 17066 18122 17066 18122 0 _0706_
rlabel metal2 16698 17289 16698 17289 0 _0707_
rlabel metal1 16928 17306 16928 17306 0 _0708_
rlabel metal1 16974 17714 16974 17714 0 _0709_
rlabel metal2 20102 15164 20102 15164 0 _0710_
rlabel metal1 19734 15572 19734 15572 0 _0711_
rlabel metal1 19642 14858 19642 14858 0 _0712_
rlabel metal1 17526 15538 17526 15538 0 _0713_
rlabel metal1 16836 15130 16836 15130 0 _0714_
rlabel metal1 17112 16082 17112 16082 0 _0715_
rlabel metal2 17434 15674 17434 15674 0 _0716_
rlabel metal1 20654 15062 20654 15062 0 _0717_
rlabel metal2 19274 16014 19274 16014 0 _0718_
rlabel metal1 18124 16626 18124 16626 0 _0719_
rlabel metal1 18032 16762 18032 16762 0 _0720_
rlabel metal1 21942 14926 21942 14926 0 _0721_
rlabel metal1 15042 14960 15042 14960 0 _0722_
rlabel metal1 15870 14994 15870 14994 0 _0723_
rlabel metal2 16330 13498 16330 13498 0 _0724_
rlabel metal1 15456 14586 15456 14586 0 _0725_
rlabel metal1 14950 15062 14950 15062 0 _0726_
rlabel metal1 17848 12818 17848 12818 0 _0727_
rlabel metal1 17480 12410 17480 12410 0 _0728_
rlabel metal1 16744 13158 16744 13158 0 _0729_
rlabel metal1 16698 12818 16698 12818 0 _0730_
rlabel metal1 15870 12886 15870 12886 0 _0731_
rlabel metal1 16422 12682 16422 12682 0 _0732_
rlabel metal2 17618 14110 17618 14110 0 _0733_
rlabel metal1 15640 13362 15640 13362 0 _0734_
rlabel metal2 14858 13090 14858 13090 0 _0735_
rlabel metal1 14674 13294 14674 13294 0 _0736_
rlabel metal1 14168 12818 14168 12818 0 _0737_
rlabel metal1 17664 13702 17664 13702 0 _0738_
rlabel metal2 17986 14518 17986 14518 0 _0739_
rlabel metal2 13938 13804 13938 13804 0 _0740_
rlabel metal2 14398 13498 14398 13498 0 _0741_
rlabel metal2 14398 14297 14398 14297 0 _0742_
rlabel metal1 14030 13498 14030 13498 0 _0743_
rlabel metal2 18630 14212 18630 14212 0 _0744_
rlabel metal1 18354 14586 18354 14586 0 _0745_
rlabel metal2 17802 15538 17802 15538 0 _0746_
rlabel metal1 14030 16116 14030 16116 0 _0747_
rlabel viali 13754 16081 13754 16081 0 _0748_
rlabel metal1 15824 14518 15824 14518 0 _0749_
rlabel metal2 13202 14756 13202 14756 0 _0750_
rlabel via1 12558 16235 12558 16235 0 _0751_
rlabel metal2 13294 15164 13294 15164 0 _0752_
rlabel metal1 10810 15028 10810 15028 0 _0753_
rlabel metal1 9752 17782 9752 17782 0 _0754_
rlabel metal1 9660 18326 9660 18326 0 _0755_
rlabel metal1 9890 18394 9890 18394 0 _0756_
rlabel metal2 5566 17986 5566 17986 0 _0757_
rlabel metal2 6118 17952 6118 17952 0 _0758_
rlabel metal1 6900 17646 6900 17646 0 _0759_
rlabel metal2 4094 17119 4094 17119 0 _0760_
rlabel metal1 7590 17680 7590 17680 0 _0761_
rlabel metal2 3082 17952 3082 17952 0 _0762_
rlabel metal1 2990 17680 2990 17680 0 _0763_
rlabel metal1 2254 16456 2254 16456 0 _0764_
rlabel metal2 1426 14110 1426 14110 0 _0765_
rlabel metal1 2714 16592 2714 16592 0 _0766_
rlabel metal1 2070 12104 2070 12104 0 _0767_
rlabel metal1 1978 12240 1978 12240 0 _0768_
rlabel metal1 1882 14042 1882 14042 0 _0769_
rlabel metal1 1978 14382 1978 14382 0 _0770_
rlabel metal2 1794 14076 1794 14076 0 _0771_
rlabel metal2 1978 14790 1978 14790 0 _0772_
rlabel metal1 2530 26860 2530 26860 0 _0773_
rlabel metal1 9430 26010 9430 26010 0 _0774_
rlabel metal2 8050 25228 8050 25228 0 _0775_
rlabel metal1 7958 24378 7958 24378 0 _0776_
rlabel metal1 8188 26554 8188 26554 0 _0777_
rlabel metal2 7222 23936 7222 23936 0 _0778_
rlabel metal2 7130 24072 7130 24072 0 _0779_
rlabel metal1 2530 23766 2530 23766 0 _0780_
rlabel metal1 3404 23290 3404 23290 0 _0781_
rlabel metal1 1932 24786 1932 24786 0 _0782_
rlabel metal2 2990 24582 2990 24582 0 _0783_
rlabel metal1 1978 27098 1978 27098 0 _0784_
rlabel metal1 1748 27098 1748 27098 0 _0785_
rlabel metal1 2898 26826 2898 26826 0 _0786_
rlabel metal1 9384 26214 9384 26214 0 bcd_num\[0\]
rlabel metal1 6440 25874 6440 25874 0 bcd_num\[1\]
rlabel metal2 8786 26588 8786 26588 0 bcd_num\[2\]
rlabel metal2 5842 24310 5842 24310 0 bcd_num\[3\]
rlabel metal1 3312 24174 3312 24174 0 bcd_num\[4\]
rlabel metal1 4600 27982 4600 27982 0 bcd_num\[5\]
rlabel metal2 3450 27370 3450 27370 0 bcd_num\[6\]
rlabel metal2 2622 27166 2622 27166 0 bcd_num\[7\]
rlabel metal1 15226 23086 15226 23086 0 clknet_0_CLK_10MHZ
rlabel metal1 1426 11764 1426 11764 0 clknet_3_0__leaf_CLK_10MHZ
rlabel metal1 1426 20842 1426 20842 0 clknet_3_1__leaf_CLK_10MHZ
rlabel via1 2438 22073 2438 22073 0 clknet_3_2__leaf_CLK_10MHZ
rlabel metal2 10074 24378 10074 24378 0 clknet_3_3__leaf_CLK_10MHZ
rlabel metal1 13524 13906 13524 13906 0 clknet_3_4__leaf_CLK_10MHZ
rlabel metal1 14674 24174 14674 24174 0 clknet_3_5__leaf_CLK_10MHZ
rlabel metal1 13386 24684 13386 24684 0 clknet_3_6__leaf_CLK_10MHZ
rlabel metal1 18584 24786 18584 24786 0 clknet_3_7__leaf_CLK_10MHZ
rlabel metal1 10902 21114 10902 21114 0 clock_div.cycles\[0\]
rlabel metal1 18492 22542 18492 22542 0 clock_div.cycles\[10\]
rlabel metal2 16100 22610 16100 22610 0 clock_div.cycles\[11\]
rlabel metal1 15732 20434 15732 20434 0 clock_div.cycles\[12\]
rlabel metal1 14260 19754 14260 19754 0 clock_div.cycles\[13\]
rlabel metal1 10672 11730 10672 11730 0 clock_div.cycles\[14\]
rlabel metal1 17756 17646 17756 17646 0 clock_div.cycles\[15\]
rlabel metal1 17434 15674 17434 15674 0 clock_div.cycles\[16\]
rlabel metal1 17710 16558 17710 16558 0 clock_div.cycles\[17\]
rlabel metal2 10258 16558 10258 16558 0 clock_div.cycles\[18\]
rlabel metal2 10626 16422 10626 16422 0 clock_div.cycles\[19\]
rlabel metal1 10534 21998 10534 21998 0 clock_div.cycles\[1\]
rlabel metal2 14030 14790 14030 14790 0 clock_div.cycles\[20\]
rlabel metal1 13294 14348 13294 14348 0 clock_div.cycles\[21\]
rlabel metal2 12834 15232 12834 15232 0 clock_div.cycles\[22\]
rlabel via1 13018 14586 13018 14586 0 clock_div.cycles\[23\]
rlabel metal2 6118 15232 6118 15232 0 clock_div.cycles\[24\]
rlabel metal1 5520 13838 5520 13838 0 clock_div.cycles\[25\]
rlabel metal1 10810 18258 10810 18258 0 clock_div.cycles\[26\]
rlabel metal1 4554 15028 4554 15028 0 clock_div.cycles\[27\]
rlabel metal2 3266 14722 3266 14722 0 clock_div.cycles\[28\]
rlabel metal1 2484 12206 2484 12206 0 clock_div.cycles\[29\]
rlabel metal1 10488 24786 10488 24786 0 clock_div.cycles\[2\]
rlabel metal1 1886 13498 1886 13498 0 clock_div.cycles\[30\]
rlabel metal1 1610 14450 1610 14450 0 clock_div.cycles\[31\]
rlabel metal2 12098 23868 12098 23868 0 clock_div.cycles\[3\]
rlabel metal1 13110 22202 13110 22202 0 clock_div.cycles\[4\]
rlabel metal1 13846 23596 13846 23596 0 clock_div.cycles\[5\]
rlabel metal1 14536 22746 14536 22746 0 clock_div.cycles\[6\]
rlabel metal1 18400 20910 18400 20910 0 clock_div.cycles\[7\]
rlabel metal1 13340 19346 13340 19346 0 clock_div.cycles\[8\]
rlabel metal1 21022 23222 21022 23222 0 clock_div.cycles\[9\]
rlabel metal1 8556 25874 8556 25874 0 clock_div.second_tick
rlabel metal1 20608 24786 20608 24786 0 digit_scanner.period_counter\[0\]
rlabel metal1 14950 26962 14950 26962 0 digit_scanner.period_counter\[10\]
rlabel metal1 15824 27846 15824 27846 0 digit_scanner.period_counter\[11\]
rlabel metal2 14030 27676 14030 27676 0 digit_scanner.period_counter\[12\]
rlabel metal1 12926 26214 12926 26214 0 digit_scanner.period_counter\[13\]
rlabel metal1 12558 26316 12558 26316 0 digit_scanner.period_counter\[14\]
rlabel metal2 12650 27030 12650 27030 0 digit_scanner.period_counter\[15\]
rlabel metal1 20148 25670 20148 25670 0 digit_scanner.period_counter\[1\]
rlabel metal1 21022 25466 21022 25466 0 digit_scanner.period_counter\[2\]
rlabel metal1 20654 26860 20654 26860 0 digit_scanner.period_counter\[3\]
rlabel metal1 16836 26214 16836 26214 0 digit_scanner.period_counter\[4\]
rlabel metal1 17250 25908 17250 25908 0 digit_scanner.period_counter\[5\]
rlabel metal1 17250 26214 17250 26214 0 digit_scanner.period_counter\[6\]
rlabel metal1 17526 24276 17526 24276 0 digit_scanner.period_counter\[7\]
rlabel metal1 16146 25466 16146 25466 0 digit_scanner.period_counter\[8\]
rlabel metal1 14352 26010 14352 26010 0 digit_scanner.period_counter\[9\]
rlabel metal1 7406 20298 7406 20298 0 fsm_inst1.currentState\[0\]
rlabel metal1 6670 21080 6670 21080 0 fsm_inst1.currentState\[1\]
rlabel metal1 8275 28118 8275 28118 0 net1
rlabel metal1 1702 26316 1702 26316 0 net10
rlabel metal2 14306 14076 14306 14076 0 net100
rlabel metal1 8372 17714 8372 17714 0 net101
rlabel metal1 14352 25874 14352 25874 0 net102
rlabel metal1 1702 24752 1702 24752 0 net11
rlabel metal2 6210 28356 6210 28356 0 net12
rlabel metal1 7084 28050 7084 28050 0 net13
rlabel metal1 21988 15674 21988 15674 0 net14
rlabel metal1 19182 17646 19182 17646 0 net15
rlabel metal1 23506 20978 23506 20978 0 net16
rlabel metal2 23230 20638 23230 20638 0 net17
rlabel metal1 25254 14892 25254 14892 0 net18
rlabel metal1 23660 15470 23660 15470 0 net19
rlabel via1 1697 21998 1697 21998 0 net2
rlabel metal1 25116 15334 25116 15334 0 net20
rlabel metal2 20010 7548 20010 7548 0 net21
rlabel metal2 21114 9945 21114 9945 0 net22
rlabel metal1 21160 16762 21160 16762 0 net23
rlabel metal2 17112 10030 17112 10030 0 net24
rlabel metal1 17710 8432 17710 8432 0 net25
rlabel metal1 10856 2414 10856 2414 0 net26
rlabel metal2 11086 8160 11086 8160 0 net27
rlabel metal1 11730 6766 11730 6766 0 net28
rlabel metal1 7038 9554 7038 9554 0 net29
rlabel via1 1697 19346 1697 19346 0 net3
rlabel metal2 2116 12206 2116 12206 0 net30
rlabel metal2 21850 13906 21850 13906 0 net31
rlabel metal2 20654 21012 20654 21012 0 net32
rlabel metal1 13570 22474 13570 22474 0 net33
rlabel metal1 14306 20230 14306 20230 0 net34
rlabel metal1 15686 17646 15686 17646 0 net35
rlabel metal1 12696 22950 12696 22950 0 net36
rlabel metal1 9982 13294 9982 13294 0 net37
rlabel metal2 4002 23664 4002 23664 0 net38
rlabel via1 2323 12206 2323 12206 0 net39
rlabel viali 1697 20910 1697 20910 0 net4
rlabel via1 14319 19414 14319 19414 0 net40
rlabel metal2 18722 22304 18722 22304 0 net41
rlabel metal2 14122 20434 14122 20434 0 net42
rlabel metal1 4002 25228 4002 25228 0 net43
rlabel metal1 4784 27030 4784 27030 0 net44
rlabel metal1 6624 26418 6624 26418 0 net45
rlabel metal1 16698 15028 16698 15028 0 net46
rlabel metal1 13570 17578 13570 17578 0 net47
rlabel metal1 15226 19992 15226 19992 0 net48
rlabel metal1 15502 19312 15502 19312 0 net49
rlabel metal2 1886 26112 1886 26112 0 net5
rlabel metal1 19642 16558 19642 16558 0 net50
rlabel metal1 21252 23290 21252 23290 0 net51
rlabel metal3 751 2788 751 2788 0 net52
rlabel metal1 3312 28594 3312 28594 0 net53
rlabel metal2 27554 2873 27554 2873 0 net54
rlabel metal1 8433 28458 8433 28458 0 net55
rlabel metal2 2898 21318 2898 21318 0 net56
rlabel metal1 2617 19754 2617 19754 0 net57
rlabel metal1 2617 22678 2617 22678 0 net58
rlabel via1 4089 19346 4089 19346 0 net59
rlabel metal1 9522 28186 9522 28186 0 net6
rlabel metal1 3992 21998 3992 21998 0 net60
rlabel metal1 4917 20842 4917 20842 0 net61
rlabel metal1 7861 21590 7861 21590 0 net62
rlabel metal1 19458 23732 19458 23732 0 net63
rlabel metal1 17940 15470 17940 15470 0 net64
rlabel metal1 19964 26350 19964 26350 0 net65
rlabel metal1 11408 28050 11408 28050 0 net66
rlabel metal1 20424 25262 20424 25262 0 net67
rlabel metal1 20930 25874 20930 25874 0 net68
rlabel metal1 19458 22678 19458 22678 0 net69
rlabel metal1 1702 25296 1702 25296 0 net7
rlabel metal1 14030 27370 14030 27370 0 net70
rlabel metal1 12742 27642 12742 27642 0 net71
rlabel metal1 17572 19346 17572 19346 0 net72
rlabel metal1 13156 26282 13156 26282 0 net73
rlabel metal1 11730 25874 11730 25874 0 net74
rlabel metal1 17756 17714 17756 17714 0 net75
rlabel metal1 19550 23664 19550 23664 0 net76
rlabel metal1 10534 23630 10534 23630 0 net77
rlabel via1 12102 24174 12102 24174 0 net78
rlabel metal1 13846 23086 13846 23086 0 net79
rlabel metal2 2254 24174 2254 24174 0 net8
rlabel metal1 13248 25126 13248 25126 0 net80
rlabel metal1 17664 22678 17664 22678 0 net81
rlabel metal1 16744 24174 16744 24174 0 net82
rlabel metal2 14306 27132 14306 27132 0 net83
rlabel metal1 17572 27438 17572 27438 0 net84
rlabel metal1 19376 28050 19376 28050 0 net85
rlabel metal1 12834 23018 12834 23018 0 net86
rlabel metal2 2622 16626 2622 16626 0 net87
rlabel metal1 9476 20434 9476 20434 0 net88
rlabel metal1 8832 25126 8832 25126 0 net89
rlabel metal2 5566 27268 5566 27268 0 net9
rlabel metal1 10544 26350 10544 26350 0 net90
rlabel metal2 2254 14110 2254 14110 0 net91
rlabel metal2 12190 21641 12190 21641 0 net92
rlabel metal1 15364 23698 15364 23698 0 net93
rlabel metal2 13294 16252 13294 16252 0 net94
rlabel metal1 3496 27098 3496 27098 0 net95
rlabel metal1 19136 21658 19136 21658 0 net96
rlabel metal1 13800 12886 13800 12886 0 net97
rlabel metal1 10810 27506 10810 27506 0 net98
rlabel metal1 17066 25772 17066 25772 0 net99
rlabel metal1 5244 20434 5244 20434 0 sync_clear.q
rlabel metal1 3450 20978 3450 20978 0 sync_clear.sync_1
rlabel metal1 4002 21420 4002 21420 0 sync_clear.sync_2
rlabel metal1 8924 21522 8924 21522 0 sync_one.q
rlabel metal2 9154 28356 9154 28356 0 sync_one.sync_1
rlabel metal1 6854 21420 6854 21420 0 sync_one.sync_2
rlabel metal1 5658 19482 5658 19482 0 sync_pause.q
rlabel metal1 2806 19278 2806 19278 0 sync_pause.sync_1
rlabel metal1 5474 20366 5474 20366 0 sync_pause.sync_2
rlabel metal1 5244 21862 5244 21862 0 sync_ten.q
rlabel metal1 3036 22202 3036 22202 0 sync_ten.sync_1
rlabel metal1 4968 21454 4968 21454 0 sync_ten.sync_2
<< properties >>
string FIXED_BBOX 0 0 29020 31164
<< end >>
