VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fpgacell
  CLASS BLOCK ;
  FOREIGN fpgacell ;
  ORIGIN 0.000 0.000 ;
  SIZE 185.000 BY 185.000 ;
  PIN CBeast_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 181.000 93.880 185.000 94.480 ;
    END
  END CBeast_in[0]
  PIN CBeast_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.028400 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 181.000 148.280 185.000 148.880 ;
    END
  END CBeast_in[10]
  PIN CBeast_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 181.000 153.720 185.000 154.320 ;
    END
  END CBeast_in[11]
  PIN CBeast_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 181.000 159.160 185.000 159.760 ;
    END
  END CBeast_in[12]
  PIN CBeast_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 181.000 164.600 185.000 165.200 ;
    END
  END CBeast_in[13]
  PIN CBeast_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 181.000 99.320 185.000 99.920 ;
    END
  END CBeast_in[1]
  PIN CBeast_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 181.000 104.760 185.000 105.360 ;
    END
  END CBeast_in[2]
  PIN CBeast_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 181.000 110.200 185.000 110.800 ;
    END
  END CBeast_in[3]
  PIN CBeast_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 181.000 115.640 185.000 116.240 ;
    END
  END CBeast_in[4]
  PIN CBeast_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 181.000 121.080 185.000 121.680 ;
    END
  END CBeast_in[5]
  PIN CBeast_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 181.000 126.520 185.000 127.120 ;
    END
  END CBeast_in[6]
  PIN CBeast_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 181.000 131.960 185.000 132.560 ;
    END
  END CBeast_in[7]
  PIN CBeast_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 181.000 137.400 185.000 138.000 ;
    END
  END CBeast_in[8]
  PIN CBeast_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.028400 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met3 ;
        RECT 181.000 142.840 185.000 143.440 ;
    END
  END CBeast_in[9]
  PIN CBeast_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 181.000 17.720 185.000 18.320 ;
    END
  END CBeast_out[0]
  PIN CBeast_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 181.000 72.120 185.000 72.720 ;
    END
  END CBeast_out[10]
  PIN CBeast_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 181.000 77.560 185.000 78.160 ;
    END
  END CBeast_out[11]
  PIN CBeast_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 181.000 83.000 185.000 83.600 ;
    END
  END CBeast_out[12]
  PIN CBeast_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 181.000 88.440 185.000 89.040 ;
    END
  END CBeast_out[13]
  PIN CBeast_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 181.000 23.160 185.000 23.760 ;
    END
  END CBeast_out[1]
  PIN CBeast_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 181.000 28.600 185.000 29.200 ;
    END
  END CBeast_out[2]
  PIN CBeast_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 181.000 34.040 185.000 34.640 ;
    END
  END CBeast_out[3]
  PIN CBeast_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 181.000 39.480 185.000 40.080 ;
    END
  END CBeast_out[4]
  PIN CBeast_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 181.000 44.920 185.000 45.520 ;
    END
  END CBeast_out[5]
  PIN CBeast_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 181.000 50.360 185.000 50.960 ;
    END
  END CBeast_out[6]
  PIN CBeast_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 181.000 55.800 185.000 56.400 ;
    END
  END CBeast_out[7]
  PIN CBeast_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 181.000 61.240 185.000 61.840 ;
    END
  END CBeast_out[8]
  PIN CBeast_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 181.000 66.680 185.000 67.280 ;
    END
  END CBeast_out[9]
  PIN CBnorth_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.028400 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 27.690 181.000 27.970 185.000 ;
    END
  END CBnorth_in[0]
  PIN CBnorth_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 82.890 181.000 83.170 185.000 ;
    END
  END CBnorth_in[10]
  PIN CBnorth_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 88.410 181.000 88.690 185.000 ;
    END
  END CBnorth_in[11]
  PIN CBnorth_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.028400 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 93.930 181.000 94.210 185.000 ;
    END
  END CBnorth_in[12]
  PIN CBnorth_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 99.450 181.000 99.730 185.000 ;
    END
  END CBnorth_in[13]
  PIN CBnorth_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.028400 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 33.210 181.000 33.490 185.000 ;
    END
  END CBnorth_in[1]
  PIN CBnorth_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 38.730 181.000 39.010 185.000 ;
    END
  END CBnorth_in[2]
  PIN CBnorth_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 44.250 181.000 44.530 185.000 ;
    END
  END CBnorth_in[3]
  PIN CBnorth_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 49.770 181.000 50.050 185.000 ;
    END
  END CBnorth_in[4]
  PIN CBnorth_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 55.290 181.000 55.570 185.000 ;
    END
  END CBnorth_in[5]
  PIN CBnorth_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 60.810 181.000 61.090 185.000 ;
    END
  END CBnorth_in[6]
  PIN CBnorth_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 66.330 181.000 66.610 185.000 ;
    END
  END CBnorth_in[7]
  PIN CBnorth_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 71.850 181.000 72.130 185.000 ;
    END
  END CBnorth_in[8]
  PIN CBnorth_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 77.370 181.000 77.650 185.000 ;
    END
  END CBnorth_in[9]
  PIN CBnorth_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 104.970 181.000 105.250 185.000 ;
    END
  END CBnorth_out[0]
  PIN CBnorth_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 160.170 181.000 160.450 185.000 ;
    END
  END CBnorth_out[10]
  PIN CBnorth_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 165.690 181.000 165.970 185.000 ;
    END
  END CBnorth_out[11]
  PIN CBnorth_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 171.210 181.000 171.490 185.000 ;
    END
  END CBnorth_out[12]
  PIN CBnorth_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 176.730 181.000 177.010 185.000 ;
    END
  END CBnorth_out[13]
  PIN CBnorth_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 110.490 181.000 110.770 185.000 ;
    END
  END CBnorth_out[1]
  PIN CBnorth_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 116.010 181.000 116.290 185.000 ;
    END
  END CBnorth_out[2]
  PIN CBnorth_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 121.530 181.000 121.810 185.000 ;
    END
  END CBnorth_out[3]
  PIN CBnorth_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 127.050 181.000 127.330 185.000 ;
    END
  END CBnorth_out[4]
  PIN CBnorth_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 132.570 181.000 132.850 185.000 ;
    END
  END CBnorth_out[5]
  PIN CBnorth_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 138.090 181.000 138.370 185.000 ;
    END
  END CBnorth_out[6]
  PIN CBnorth_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 143.610 181.000 143.890 185.000 ;
    END
  END CBnorth_out[7]
  PIN CBnorth_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 149.130 181.000 149.410 185.000 ;
    END
  END CBnorth_out[8]
  PIN CBnorth_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 154.650 181.000 154.930 185.000 ;
    END
  END CBnorth_out[9]
  PIN SBsouth_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 107.730 0.000 108.010 4.000 ;
    END
  END SBsouth_in[0]
  PIN SBsouth_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 162.930 0.000 163.210 4.000 ;
    END
  END SBsouth_in[10]
  PIN SBsouth_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 168.450 0.000 168.730 4.000 ;
    END
  END SBsouth_in[11]
  PIN SBsouth_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END SBsouth_in[12]
  PIN SBsouth_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 179.490 0.000 179.770 4.000 ;
    END
  END SBsouth_in[13]
  PIN SBsouth_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 113.250 0.000 113.530 4.000 ;
    END
  END SBsouth_in[1]
  PIN SBsouth_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 118.770 0.000 119.050 4.000 ;
    END
  END SBsouth_in[2]
  PIN SBsouth_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 124.290 0.000 124.570 4.000 ;
    END
  END SBsouth_in[3]
  PIN SBsouth_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 130.090 4.000 ;
    END
  END SBsouth_in[4]
  PIN SBsouth_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END SBsouth_in[5]
  PIN SBsouth_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 140.850 0.000 141.130 4.000 ;
    END
  END SBsouth_in[6]
  PIN SBsouth_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 146.370 0.000 146.650 4.000 ;
    END
  END SBsouth_in[7]
  PIN SBsouth_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 151.890 0.000 152.170 4.000 ;
    END
  END SBsouth_in[8]
  PIN SBsouth_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 157.410 0.000 157.690 4.000 ;
    END
  END SBsouth_in[9]
  PIN SBsouth_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 30.450 0.000 30.730 4.000 ;
    END
  END SBsouth_out[0]
  PIN SBsouth_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 85.650 0.000 85.930 4.000 ;
    END
  END SBsouth_out[10]
  PIN SBsouth_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 91.170 0.000 91.450 4.000 ;
    END
  END SBsouth_out[11]
  PIN SBsouth_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END SBsouth_out[12]
  PIN SBsouth_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 4.000 ;
    END
  END SBsouth_out[13]
  PIN SBsouth_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 35.970 0.000 36.250 4.000 ;
    END
  END SBsouth_out[1]
  PIN SBsouth_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 41.490 0.000 41.770 4.000 ;
    END
  END SBsouth_out[2]
  PIN SBsouth_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 4.000 ;
    END
  END SBsouth_out[3]
  PIN SBsouth_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 52.530 0.000 52.810 4.000 ;
    END
  END SBsouth_out[4]
  PIN SBsouth_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END SBsouth_out[5]
  PIN SBsouth_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 63.570 0.000 63.850 4.000 ;
    END
  END SBsouth_out[6]
  PIN SBsouth_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END SBsouth_out[7]
  PIN SBsouth_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 4.000 ;
    END
  END SBsouth_out[8]
  PIN SBsouth_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 80.130 0.000 80.410 4.000 ;
    END
  END SBsouth_out[9]
  PIN SBwest_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 4.000 18.320 ;
    END
  END SBwest_in[0]
  PIN SBwest_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 4.000 72.720 ;
    END
  END SBwest_in[10]
  PIN SBwest_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.560 4.000 78.160 ;
    END
  END SBwest_in[11]
  PIN SBwest_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 4.000 83.600 ;
    END
  END SBwest_in[12]
  PIN SBwest_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END SBwest_in[13]
  PIN SBwest_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.160 4.000 23.760 ;
    END
  END SBwest_in[1]
  PIN SBwest_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 4.000 29.200 ;
    END
  END SBwest_in[2]
  PIN SBwest_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END SBwest_in[3]
  PIN SBwest_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END SBwest_in[4]
  PIN SBwest_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 4.000 45.520 ;
    END
  END SBwest_in[5]
  PIN SBwest_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 4.000 50.960 ;
    END
  END SBwest_in[6]
  PIN SBwest_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 4.000 56.400 ;
    END
  END SBwest_in[7]
  PIN SBwest_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END SBwest_in[8]
  PIN SBwest_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.680 4.000 67.280 ;
    END
  END SBwest_in[9]
  PIN SBwest_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 4.000 94.480 ;
    END
  END SBwest_out[0]
  PIN SBwest_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.280 4.000 148.880 ;
    END
  END SBwest_out[10]
  PIN SBwest_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.720 4.000 154.320 ;
    END
  END SBwest_out[11]
  PIN SBwest_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.160 4.000 159.760 ;
    END
  END SBwest_out[12]
  PIN SBwest_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.600 4.000 165.200 ;
    END
  END SBwest_out[13]
  PIN SBwest_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.320 4.000 99.920 ;
    END
  END SBwest_out[1]
  PIN SBwest_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.760 4.000 105.360 ;
    END
  END SBwest_out[2]
  PIN SBwest_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 4.000 110.800 ;
    END
  END SBwest_out[3]
  PIN SBwest_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END SBwest_out[4]
  PIN SBwest_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 4.000 121.680 ;
    END
  END SBwest_out[5]
  PIN SBwest_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 4.000 127.120 ;
    END
  END SBwest_out[6]
  PIN SBwest_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.960 4.000 132.560 ;
    END
  END SBwest_out[7]
  PIN SBwest_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END SBwest_out[8]
  PIN SBwest_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END SBwest_out[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 5.610 181.000 5.890 185.000 ;
    END
  END clk
  PIN config_data_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 22.170 181.000 22.450 185.000 ;
    END
  END config_data_in
  PIN config_data_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END config_data_out
  PIN config_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 16.650 181.000 16.930 185.000 ;
    END
  END config_en
  PIN le_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 8.370 0.000 8.650 4.000 ;
    END
  END le_clk
  PIN le_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 13.890 0.000 14.170 4.000 ;
    END
  END le_en
  PIN le_nrst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END le_nrst
  PIN nrst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 11.130 181.000 11.410 185.000 ;
    END
  END nrst
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2.420 4.640 4.020 179.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 172.420 4.640 174.020 179.760 ;
    END
    PORT
      LAYER met5 ;
        RECT 2.420 4.640 181.940 6.240 ;
    END
    PORT
      LAYER met5 ;
        RECT 2.420 174.640 181.940 176.240 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 5.720 5.200 7.320 179.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 175.720 5.200 177.320 179.760 ;
    END
    PORT
      LAYER met5 ;
        RECT 2.980 7.940 181.940 9.540 ;
    END
    PORT
      LAYER met5 ;
        RECT 2.980 177.940 181.940 179.540 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 3.030 5.355 181.890 179.605 ;
      LAYER li1 ;
        RECT 3.220 5.355 181.700 179.605 ;
      LAYER met1 ;
        RECT 0.070 1.400 183.930 184.240 ;
      LAYER met2 ;
        RECT 0.090 180.720 5.330 184.270 ;
        RECT 6.170 180.720 10.850 184.270 ;
        RECT 11.690 180.720 16.370 184.270 ;
        RECT 17.210 180.720 21.890 184.270 ;
        RECT 22.730 180.720 27.410 184.270 ;
        RECT 28.250 180.720 32.930 184.270 ;
        RECT 33.770 180.720 38.450 184.270 ;
        RECT 39.290 180.720 43.970 184.270 ;
        RECT 44.810 180.720 49.490 184.270 ;
        RECT 50.330 180.720 55.010 184.270 ;
        RECT 55.850 180.720 60.530 184.270 ;
        RECT 61.370 180.720 66.050 184.270 ;
        RECT 66.890 180.720 71.570 184.270 ;
        RECT 72.410 180.720 77.090 184.270 ;
        RECT 77.930 180.720 82.610 184.270 ;
        RECT 83.450 180.720 88.130 184.270 ;
        RECT 88.970 180.720 93.650 184.270 ;
        RECT 94.490 180.720 99.170 184.270 ;
        RECT 100.010 180.720 104.690 184.270 ;
        RECT 105.530 180.720 110.210 184.270 ;
        RECT 111.050 180.720 115.730 184.270 ;
        RECT 116.570 180.720 121.250 184.270 ;
        RECT 122.090 180.720 126.770 184.270 ;
        RECT 127.610 180.720 132.290 184.270 ;
        RECT 133.130 180.720 137.810 184.270 ;
        RECT 138.650 180.720 143.330 184.270 ;
        RECT 144.170 180.720 148.850 184.270 ;
        RECT 149.690 180.720 154.370 184.270 ;
        RECT 155.210 180.720 159.890 184.270 ;
        RECT 160.730 180.720 165.410 184.270 ;
        RECT 166.250 180.720 170.930 184.270 ;
        RECT 171.770 180.720 176.450 184.270 ;
        RECT 177.290 180.720 183.900 184.270 ;
        RECT 0.090 4.280 183.900 180.720 ;
        RECT 0.090 1.370 2.570 4.280 ;
        RECT 3.410 1.370 8.090 4.280 ;
        RECT 8.930 1.370 13.610 4.280 ;
        RECT 14.450 1.370 19.130 4.280 ;
        RECT 19.970 1.370 30.170 4.280 ;
        RECT 31.010 1.370 35.690 4.280 ;
        RECT 36.530 1.370 41.210 4.280 ;
        RECT 42.050 1.370 46.730 4.280 ;
        RECT 47.570 1.370 52.250 4.280 ;
        RECT 53.090 1.370 57.770 4.280 ;
        RECT 58.610 1.370 63.290 4.280 ;
        RECT 64.130 1.370 68.810 4.280 ;
        RECT 69.650 1.370 74.330 4.280 ;
        RECT 75.170 1.370 79.850 4.280 ;
        RECT 80.690 1.370 85.370 4.280 ;
        RECT 86.210 1.370 90.890 4.280 ;
        RECT 91.730 1.370 96.410 4.280 ;
        RECT 97.250 1.370 101.930 4.280 ;
        RECT 102.770 1.370 107.450 4.280 ;
        RECT 108.290 1.370 112.970 4.280 ;
        RECT 113.810 1.370 118.490 4.280 ;
        RECT 119.330 1.370 124.010 4.280 ;
        RECT 124.850 1.370 129.530 4.280 ;
        RECT 130.370 1.370 135.050 4.280 ;
        RECT 135.890 1.370 140.570 4.280 ;
        RECT 141.410 1.370 146.090 4.280 ;
        RECT 146.930 1.370 151.610 4.280 ;
        RECT 152.450 1.370 157.130 4.280 ;
        RECT 157.970 1.370 162.650 4.280 ;
        RECT 163.490 1.370 168.170 4.280 ;
        RECT 169.010 1.370 173.690 4.280 ;
        RECT 174.530 1.370 179.210 4.280 ;
        RECT 180.050 1.370 183.900 4.280 ;
      LAYER met3 ;
        RECT 0.065 165.600 182.555 180.705 ;
        RECT 4.400 164.200 180.600 165.600 ;
        RECT 0.065 160.160 182.555 164.200 ;
        RECT 4.400 158.760 180.600 160.160 ;
        RECT 0.065 154.720 182.555 158.760 ;
        RECT 4.400 153.320 180.600 154.720 ;
        RECT 0.065 149.280 182.555 153.320 ;
        RECT 4.400 147.880 180.600 149.280 ;
        RECT 0.065 143.840 182.555 147.880 ;
        RECT 4.400 142.440 180.600 143.840 ;
        RECT 0.065 138.400 182.555 142.440 ;
        RECT 4.400 137.000 180.600 138.400 ;
        RECT 0.065 132.960 182.555 137.000 ;
        RECT 4.400 131.560 180.600 132.960 ;
        RECT 0.065 127.520 182.555 131.560 ;
        RECT 4.400 126.120 180.600 127.520 ;
        RECT 0.065 122.080 182.555 126.120 ;
        RECT 4.400 120.680 180.600 122.080 ;
        RECT 0.065 116.640 182.555 120.680 ;
        RECT 4.400 115.240 180.600 116.640 ;
        RECT 0.065 111.200 182.555 115.240 ;
        RECT 4.400 109.800 180.600 111.200 ;
        RECT 0.065 105.760 182.555 109.800 ;
        RECT 4.400 104.360 180.600 105.760 ;
        RECT 0.065 100.320 182.555 104.360 ;
        RECT 4.400 98.920 180.600 100.320 ;
        RECT 0.065 94.880 182.555 98.920 ;
        RECT 4.400 93.480 180.600 94.880 ;
        RECT 0.065 89.440 182.555 93.480 ;
        RECT 4.400 88.040 180.600 89.440 ;
        RECT 0.065 84.000 182.555 88.040 ;
        RECT 4.400 82.600 180.600 84.000 ;
        RECT 0.065 78.560 182.555 82.600 ;
        RECT 4.400 77.160 180.600 78.560 ;
        RECT 0.065 73.120 182.555 77.160 ;
        RECT 4.400 71.720 180.600 73.120 ;
        RECT 0.065 67.680 182.555 71.720 ;
        RECT 4.400 66.280 180.600 67.680 ;
        RECT 0.065 62.240 182.555 66.280 ;
        RECT 4.400 60.840 180.600 62.240 ;
        RECT 0.065 56.800 182.555 60.840 ;
        RECT 4.400 55.400 180.600 56.800 ;
        RECT 0.065 51.360 182.555 55.400 ;
        RECT 4.400 49.960 180.600 51.360 ;
        RECT 0.065 45.920 182.555 49.960 ;
        RECT 4.400 44.520 180.600 45.920 ;
        RECT 0.065 40.480 182.555 44.520 ;
        RECT 4.400 39.080 180.600 40.480 ;
        RECT 0.065 35.040 182.555 39.080 ;
        RECT 4.400 33.640 180.600 35.040 ;
        RECT 0.065 29.600 182.555 33.640 ;
        RECT 4.400 28.200 180.600 29.600 ;
        RECT 0.065 24.160 182.555 28.200 ;
        RECT 4.400 22.760 180.600 24.160 ;
        RECT 0.065 18.720 182.555 22.760 ;
        RECT 4.400 17.320 180.600 18.720 ;
        RECT 0.065 5.275 182.555 17.320 ;
      LAYER met4 ;
        RECT 4.895 180.160 171.745 180.705 ;
        RECT 4.895 6.295 5.320 180.160 ;
        RECT 7.720 6.295 171.745 180.160 ;
  END
END fpgacell
END LIBRARY

