`default_nettype none
module fa (
  //put your ports here
  inout logic test,
  output logic f
);
  assign test = 1'b1;
  assign f = test;
//your code starts here ...
endmodule
