VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fpga
  CLASS BLOCK ;
  FOREIGN fpga ;
  ORIGIN 0.000 0.000 ;
  SIZE 450.000 BY 490.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 248.030 486.000 248.310 490.000 ;
    END
  END clk
  PIN config_data_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END config_data_in
  PIN config_data_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 251.640 450.000 252.240 ;
    END
  END config_data_out
  PIN config_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.424700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 260.910 486.000 261.190 490.000 ;
    END
  END config_en
  PIN io_east_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 139.440 450.000 140.040 ;
    END
  END io_east_in[0]
  PIN io_east_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 207.440 450.000 208.040 ;
    END
  END io_east_in[10]
  PIN io_east_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 214.240 450.000 214.840 ;
    END
  END io_east_in[11]
  PIN io_east_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 221.040 450.000 221.640 ;
    END
  END io_east_in[12]
  PIN io_east_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 227.840 450.000 228.440 ;
    END
  END io_east_in[13]
  PIN io_east_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END io_east_in[14]
  PIN io_east_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END io_east_in[15]
  PIN io_east_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 350.240 450.000 350.840 ;
    END
  END io_east_in[16]
  PIN io_east_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 357.040 450.000 357.640 ;
    END
  END io_east_in[17]
  PIN io_east_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 363.840 450.000 364.440 ;
    END
  END io_east_in[18]
  PIN io_east_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 370.640 450.000 371.240 ;
    END
  END io_east_in[19]
  PIN io_east_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 146.240 450.000 146.840 ;
    END
  END io_east_in[1]
  PIN io_east_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 377.440 450.000 378.040 ;
    END
  END io_east_in[20]
  PIN io_east_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 384.240 450.000 384.840 ;
    END
  END io_east_in[21]
  PIN io_east_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 391.040 450.000 391.640 ;
    END
  END io_east_in[22]
  PIN io_east_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 397.840 450.000 398.440 ;
    END
  END io_east_in[23]
  PIN io_east_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 404.640 450.000 405.240 ;
    END
  END io_east_in[24]
  PIN io_east_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 411.440 450.000 412.040 ;
    END
  END io_east_in[25]
  PIN io_east_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 418.240 450.000 418.840 ;
    END
  END io_east_in[26]
  PIN io_east_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 425.040 450.000 425.640 ;
    END
  END io_east_in[27]
  PIN io_east_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 431.840 450.000 432.440 ;
    END
  END io_east_in[28]
  PIN io_east_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 438.640 450.000 439.240 ;
    END
  END io_east_in[29]
  PIN io_east_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 153.040 450.000 153.640 ;
    END
  END io_east_in[2]
  PIN io_east_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END io_east_in[30]
  PIN io_east_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END io_east_in[31]
  PIN io_east_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 159.840 450.000 160.440 ;
    END
  END io_east_in[3]
  PIN io_east_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 166.640 450.000 167.240 ;
    END
  END io_east_in[4]
  PIN io_east_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 173.440 450.000 174.040 ;
    END
  END io_east_in[5]
  PIN io_east_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 180.240 450.000 180.840 ;
    END
  END io_east_in[6]
  PIN io_east_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 187.040 450.000 187.640 ;
    END
  END io_east_in[7]
  PIN io_east_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 193.840 450.000 194.440 ;
    END
  END io_east_in[8]
  PIN io_east_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 200.640 450.000 201.240 ;
    END
  END io_east_in[9]
  PIN io_east_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 47.640 450.000 48.240 ;
    END
  END io_east_out[0]
  PIN io_east_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 112.240 450.000 112.840 ;
    END
  END io_east_out[10]
  PIN io_east_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 119.040 450.000 119.640 ;
    END
  END io_east_out[11]
  PIN io_east_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 125.840 450.000 126.440 ;
    END
  END io_east_out[12]
  PIN io_east_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 132.640 450.000 133.240 ;
    END
  END io_east_out[13]
  PIN io_east_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.840 4.000 262.440 ;
    END
  END io_east_out[14]
  PIN io_east_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 302.640 4.000 303.240 ;
    END
  END io_east_out[15]
  PIN io_east_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 255.040 450.000 255.640 ;
    END
  END io_east_out[16]
  PIN io_east_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 261.840 450.000 262.440 ;
    END
  END io_east_out[17]
  PIN io_east_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 268.640 450.000 269.240 ;
    END
  END io_east_out[18]
  PIN io_east_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 275.440 450.000 276.040 ;
    END
  END io_east_out[19]
  PIN io_east_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 51.040 450.000 51.640 ;
    END
  END io_east_out[1]
  PIN io_east_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 282.240 450.000 282.840 ;
    END
  END io_east_out[20]
  PIN io_east_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 289.040 450.000 289.640 ;
    END
  END io_east_out[21]
  PIN io_east_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 295.840 450.000 296.440 ;
    END
  END io_east_out[22]
  PIN io_east_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 302.640 450.000 303.240 ;
    END
  END io_east_out[23]
  PIN io_east_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 309.440 450.000 310.040 ;
    END
  END io_east_out[24]
  PIN io_east_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 316.240 450.000 316.840 ;
    END
  END io_east_out[25]
  PIN io_east_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 323.040 450.000 323.640 ;
    END
  END io_east_out[26]
  PIN io_east_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 329.840 450.000 330.440 ;
    END
  END io_east_out[27]
  PIN io_east_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 336.640 450.000 337.240 ;
    END
  END io_east_out[28]
  PIN io_east_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 343.440 450.000 344.040 ;
    END
  END io_east_out[29]
  PIN io_east_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 57.840 450.000 58.440 ;
    END
  END io_east_out[2]
  PIN io_east_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END io_east_out[30]
  PIN io_east_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END io_east_out[31]
  PIN io_east_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 64.640 450.000 65.240 ;
    END
  END io_east_out[3]
  PIN io_east_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 71.440 450.000 72.040 ;
    END
  END io_east_out[4]
  PIN io_east_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 78.240 450.000 78.840 ;
    END
  END io_east_out[5]
  PIN io_east_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 85.040 450.000 85.640 ;
    END
  END io_east_out[6]
  PIN io_east_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 91.840 450.000 92.440 ;
    END
  END io_east_out[7]
  PIN io_east_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 98.640 450.000 99.240 ;
    END
  END io_east_out[8]
  PIN io_east_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 105.440 450.000 106.040 ;
    END
  END io_east_out[9]
  PIN io_north_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 74.150 486.000 74.430 490.000 ;
    END
  END io_north_in[0]
  PIN io_north_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 128.890 486.000 129.170 490.000 ;
    END
  END io_north_in[10]
  PIN io_north_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 135.330 486.000 135.610 490.000 ;
    END
  END io_north_in[11]
  PIN io_north_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 138.550 486.000 138.830 490.000 ;
    END
  END io_north_in[12]
  PIN io_north_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 144.990 486.000 145.270 490.000 ;
    END
  END io_north_in[13]
  PIN io_north_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END io_north_in[14]
  PIN io_north_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END io_north_in[15]
  PIN io_north_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 273.790 486.000 274.070 490.000 ;
    END
  END io_north_in[16]
  PIN io_north_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 280.230 486.000 280.510 490.000 ;
    END
  END io_north_in[17]
  PIN io_north_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 283.450 486.000 283.730 490.000 ;
    END
  END io_north_in[18]
  PIN io_north_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 289.890 486.000 290.170 490.000 ;
    END
  END io_north_in[19]
  PIN io_north_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 77.370 486.000 77.650 490.000 ;
    END
  END io_north_in[1]
  PIN io_north_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 296.330 486.000 296.610 490.000 ;
    END
  END io_north_in[20]
  PIN io_north_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 299.550 486.000 299.830 490.000 ;
    END
  END io_north_in[21]
  PIN io_north_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 305.990 486.000 306.270 490.000 ;
    END
  END io_north_in[22]
  PIN io_north_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 312.430 486.000 312.710 490.000 ;
    END
  END io_north_in[23]
  PIN io_north_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 318.870 486.000 319.150 490.000 ;
    END
  END io_north_in[24]
  PIN io_north_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 322.090 486.000 322.370 490.000 ;
    END
  END io_north_in[25]
  PIN io_north_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 328.530 486.000 328.810 490.000 ;
    END
  END io_north_in[26]
  PIN io_north_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 334.970 486.000 335.250 490.000 ;
    END
  END io_north_in[27]
  PIN io_north_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 338.190 486.000 338.470 490.000 ;
    END
  END io_north_in[28]
  PIN io_north_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 344.630 486.000 344.910 490.000 ;
    END
  END io_north_in[29]
  PIN io_north_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 83.810 486.000 84.090 490.000 ;
    END
  END io_north_in[2]
  PIN io_north_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END io_north_in[30]
  PIN io_north_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END io_north_in[31]
  PIN io_north_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 90.250 486.000 90.530 490.000 ;
    END
  END io_north_in[3]
  PIN io_north_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 96.690 486.000 96.970 490.000 ;
    END
  END io_north_in[4]
  PIN io_north_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 99.910 486.000 100.190 490.000 ;
    END
  END io_north_in[5]
  PIN io_north_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 106.350 486.000 106.630 490.000 ;
    END
  END io_north_in[6]
  PIN io_north_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 112.790 486.000 113.070 490.000 ;
    END
  END io_north_in[7]
  PIN io_north_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 116.010 486.000 116.290 490.000 ;
    END
  END io_north_in[8]
  PIN io_north_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 122.450 486.000 122.730 490.000 ;
    END
  END io_north_in[9]
  PIN io_north_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 151.430 486.000 151.710 490.000 ;
    END
  END io_north_out[0]
  PIN io_north_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 206.170 486.000 206.450 490.000 ;
    END
  END io_north_out[10]
  PIN io_north_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 212.610 486.000 212.890 490.000 ;
    END
  END io_north_out[11]
  PIN io_north_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 215.830 486.000 216.110 490.000 ;
    END
  END io_north_out[12]
  PIN io_north_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 222.270 486.000 222.550 490.000 ;
    END
  END io_north_out[13]
  PIN io_north_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.040 4.000 289.640 ;
    END
  END io_north_out[14]
  PIN io_north_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END io_north_out[15]
  PIN io_north_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 351.070 486.000 351.350 490.000 ;
    END
  END io_north_out[16]
  PIN io_north_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 357.510 486.000 357.790 490.000 ;
    END
  END io_north_out[17]
  PIN io_north_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 360.730 486.000 361.010 490.000 ;
    END
  END io_north_out[18]
  PIN io_north_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 367.170 486.000 367.450 490.000 ;
    END
  END io_north_out[19]
  PIN io_north_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 154.650 486.000 154.930 490.000 ;
    END
  END io_north_out[1]
  PIN io_north_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 373.610 486.000 373.890 490.000 ;
    END
  END io_north_out[20]
  PIN io_north_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 376.830 486.000 377.110 490.000 ;
    END
  END io_north_out[21]
  PIN io_north_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 383.270 486.000 383.550 490.000 ;
    END
  END io_north_out[22]
  PIN io_north_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 389.710 486.000 389.990 490.000 ;
    END
  END io_north_out[23]
  PIN io_north_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 396.150 486.000 396.430 490.000 ;
    END
  END io_north_out[24]
  PIN io_north_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 399.370 486.000 399.650 490.000 ;
    END
  END io_north_out[25]
  PIN io_north_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 405.810 486.000 406.090 490.000 ;
    END
  END io_north_out[26]
  PIN io_north_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 412.250 486.000 412.530 490.000 ;
    END
  END io_north_out[27]
  PIN io_north_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 445.440 450.000 446.040 ;
    END
  END io_north_out[28]
  PIN io_north_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 442.040 450.000 442.640 ;
    END
  END io_north_out[29]
  PIN io_north_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 161.090 486.000 161.370 490.000 ;
    END
  END io_north_out[2]
  PIN io_north_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 234.640 4.000 235.240 ;
    END
  END io_north_out[30]
  PIN io_north_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 275.440 4.000 276.040 ;
    END
  END io_north_out[31]
  PIN io_north_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 167.530 486.000 167.810 490.000 ;
    END
  END io_north_out[3]
  PIN io_north_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 173.970 486.000 174.250 490.000 ;
    END
  END io_north_out[4]
  PIN io_north_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 177.190 486.000 177.470 490.000 ;
    END
  END io_north_out[5]
  PIN io_north_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 183.630 486.000 183.910 490.000 ;
    END
  END io_north_out[6]
  PIN io_north_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 190.070 486.000 190.350 490.000 ;
    END
  END io_north_out[7]
  PIN io_north_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 193.290 486.000 193.570 490.000 ;
    END
  END io_north_out[8]
  PIN io_north_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 199.730 486.000 200.010 490.000 ;
    END
  END io_north_out[9]
  PIN io_south_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 4.000 ;
    END
  END io_south_in[0]
  PIN io_south_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 4.000 ;
    END
  END io_south_in[10]
  PIN io_south_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END io_south_in[11]
  PIN io_south_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END io_south_in[12]
  PIN io_south_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END io_south_in[13]
  PIN io_south_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END io_south_in[14]
  PIN io_south_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END io_south_in[15]
  PIN io_south_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 354.290 0.000 354.570 4.000 ;
    END
  END io_south_in[16]
  PIN io_south_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 357.510 0.000 357.790 4.000 ;
    END
  END io_south_in[17]
  PIN io_south_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 363.950 0.000 364.230 4.000 ;
    END
  END io_south_in[18]
  PIN io_south_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 370.390 0.000 370.670 4.000 ;
    END
  END io_south_in[19]
  PIN io_south_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END io_south_in[1]
  PIN io_south_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 376.830 0.000 377.110 4.000 ;
    END
  END io_south_in[20]
  PIN io_south_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 380.050 0.000 380.330 4.000 ;
    END
  END io_south_in[21]
  PIN io_south_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 386.490 0.000 386.770 4.000 ;
    END
  END io_south_in[22]
  PIN io_south_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 392.930 0.000 393.210 4.000 ;
    END
  END io_south_in[23]
  PIN io_south_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 396.150 0.000 396.430 4.000 ;
    END
  END io_south_in[24]
  PIN io_south_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 402.590 0.000 402.870 4.000 ;
    END
  END io_south_in[25]
  PIN io_south_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 409.030 0.000 409.310 4.000 ;
    END
  END io_south_in[26]
  PIN io_south_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 415.470 0.000 415.750 4.000 ;
    END
  END io_south_in[27]
  PIN io_south_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 44.240 450.000 44.840 ;
    END
  END io_south_in[28]
  PIN io_south_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 40.840 450.000 41.440 ;
    END
  END io_south_in[29]
  PIN io_south_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END io_south_in[2]
  PIN io_south_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END io_south_in[30]
  PIN io_south_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END io_south_in[31]
  PIN io_south_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END io_south_in[3]
  PIN io_south_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END io_south_in[4]
  PIN io_south_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END io_south_in[5]
  PIN io_south_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END io_south_in[6]
  PIN io_south_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END io_south_in[7]
  PIN io_south_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 196.510 0.000 196.790 4.000 ;
    END
  END io_south_in[8]
  PIN io_south_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END io_south_in[9]
  PIN io_south_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END io_south_out[0]
  PIN io_south_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END io_south_out[10]
  PIN io_south_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END io_south_out[11]
  PIN io_south_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END io_south_out[12]
  PIN io_south_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END io_south_out[13]
  PIN io_south_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.640 4.000 269.240 ;
    END
  END io_south_out[14]
  PIN io_south_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.840 4.000 296.440 ;
    END
  END io_south_out[15]
  PIN io_south_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 277.010 0.000 277.290 4.000 ;
    END
  END io_south_out[16]
  PIN io_south_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 280.230 0.000 280.510 4.000 ;
    END
  END io_south_out[17]
  PIN io_south_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 4.000 ;
    END
  END io_south_out[18]
  PIN io_south_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 293.110 0.000 293.390 4.000 ;
    END
  END io_south_out[19]
  PIN io_south_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END io_south_out[1]
  PIN io_south_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 299.550 0.000 299.830 4.000 ;
    END
  END io_south_out[20]
  PIN io_south_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 302.770 0.000 303.050 4.000 ;
    END
  END io_south_out[21]
  PIN io_south_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END io_south_out[22]
  PIN io_south_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 315.650 0.000 315.930 4.000 ;
    END
  END io_south_out[23]
  PIN io_south_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 318.870 0.000 319.150 4.000 ;
    END
  END io_south_out[24]
  PIN io_south_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 325.310 0.000 325.590 4.000 ;
    END
  END io_south_out[25]
  PIN io_south_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 331.750 0.000 332.030 4.000 ;
    END
  END io_south_out[26]
  PIN io_south_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 338.190 0.000 338.470 4.000 ;
    END
  END io_south_out[27]
  PIN io_south_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 341.410 0.000 341.690 4.000 ;
    END
  END io_south_out[28]
  PIN io_south_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 347.850 0.000 348.130 4.000 ;
    END
  END io_south_out[29]
  PIN io_south_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END io_south_out[2]
  PIN io_south_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END io_south_out[30]
  PIN io_south_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.040 4.000 255.640 ;
    END
  END io_south_out[31]
  PIN io_south_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END io_south_out[3]
  PIN io_south_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END io_south_out[4]
  PIN io_south_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END io_south_out[5]
  PIN io_south_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END io_south_out[6]
  PIN io_south_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END io_south_out[7]
  PIN io_south_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.510 4.000 ;
    END
  END io_south_out[8]
  PIN io_south_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 4.000 ;
    END
  END io_south_out[9]
  PIN io_west_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END io_west_in[0]
  PIN io_west_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END io_west_in[10]
  PIN io_west_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END io_west_in[11]
  PIN io_west_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END io_west_in[12]
  PIN io_west_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END io_west_in[13]
  PIN io_west_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END io_west_in[14]
  PIN io_west_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END io_west_in[15]
  PIN io_west_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 241.440 4.000 242.040 ;
    END
  END io_west_in[16]
  PIN io_west_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END io_west_in[17]
  PIN io_west_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END io_west_in[18]
  PIN io_west_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END io_west_in[19]
  PIN io_west_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END io_west_in[1]
  PIN io_west_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END io_west_in[20]
  PIN io_west_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END io_west_in[21]
  PIN io_west_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END io_west_in[22]
  PIN io_west_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 4.000 306.640 ;
    END
  END io_west_in[23]
  PIN io_west_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 309.440 4.000 310.040 ;
    END
  END io_west_in[24]
  PIN io_west_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.240 4.000 316.840 ;
    END
  END io_west_in[25]
  PIN io_west_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.040 4.000 323.640 ;
    END
  END io_west_in[26]
  PIN io_west_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.840 4.000 330.440 ;
    END
  END io_west_in[27]
  PIN io_west_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 336.640 4.000 337.240 ;
    END
  END io_west_in[28]
  PIN io_west_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 343.440 4.000 344.040 ;
    END
  END io_west_in[29]
  PIN io_west_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END io_west_in[2]
  PIN io_west_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END io_west_in[30]
  PIN io_west_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END io_west_in[31]
  PIN io_west_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END io_west_in[3]
  PIN io_west_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END io_west_in[4]
  PIN io_west_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END io_west_in[5]
  PIN io_west_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END io_west_in[6]
  PIN io_west_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END io_west_in[7]
  PIN io_west_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END io_west_in[8]
  PIN io_west_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END io_west_in[9]
  PIN io_west_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END io_west_out[0]
  PIN io_west_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.440 4.000 208.040 ;
    END
  END io_west_out[10]
  PIN io_west_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.240 4.000 214.840 ;
    END
  END io_west_out[11]
  PIN io_west_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.040 4.000 221.640 ;
    END
  END io_west_out[12]
  PIN io_west_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END io_west_out[13]
  PIN io_west_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.240 4.000 282.840 ;
    END
  END io_west_out[14]
  PIN io_west_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END io_west_out[15]
  PIN io_west_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.240 4.000 350.840 ;
    END
  END io_west_out[16]
  PIN io_west_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.040 4.000 357.640 ;
    END
  END io_west_out[17]
  PIN io_west_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.840 4.000 364.440 ;
    END
  END io_west_out[18]
  PIN io_west_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 4.000 371.240 ;
    END
  END io_west_out[19]
  PIN io_west_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END io_west_out[1]
  PIN io_west_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 377.440 4.000 378.040 ;
    END
  END io_west_out[20]
  PIN io_west_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.240 4.000 384.840 ;
    END
  END io_west_out[21]
  PIN io_west_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.040 4.000 391.640 ;
    END
  END io_west_out[22]
  PIN io_west_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.840 4.000 398.440 ;
    END
  END io_west_out[23]
  PIN io_west_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 404.640 4.000 405.240 ;
    END
  END io_west_out[24]
  PIN io_west_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 411.440 4.000 412.040 ;
    END
  END io_west_out[25]
  PIN io_west_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.240 4.000 418.840 ;
    END
  END io_west_out[26]
  PIN io_west_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.040 4.000 425.640 ;
    END
  END io_west_out[27]
  PIN io_west_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.840 4.000 432.440 ;
    END
  END io_west_out[28]
  PIN io_west_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 41.950 486.000 42.230 490.000 ;
    END
  END io_west_out[29]
  PIN io_west_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END io_west_out[2]
  PIN io_west_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.240 4.000 248.840 ;
    END
  END io_west_out[30]
  PIN io_west_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END io_west_out[31]
  PIN io_west_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END io_west_out[3]
  PIN io_west_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 4.000 167.240 ;
    END
  END io_west_out[4]
  PIN io_west_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.440 4.000 174.040 ;
    END
  END io_west_out[5]
  PIN io_west_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END io_west_out[6]
  PIN io_west_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END io_west_out[7]
  PIN io_west_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END io_west_out[8]
  PIN io_west_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.640 4.000 201.240 ;
    END
  END io_west_out[9]
  PIN le_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.860700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END le_clk
  PIN le_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.860700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END le_en
  PIN le_nrst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.860700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END le_nrst
  PIN nrst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.424700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 254.470 486.000 254.750 490.000 ;
    END
  END nrst
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -2.080 3.280 -0.480 486.320 ;
    END
    PORT
      LAYER met5 ;
        RECT -2.080 3.280 451.960 4.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -2.080 484.720 451.960 486.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 450.360 3.280 451.960 486.320 ;
    END
    PORT
      LAYER met4 ;
        RECT 184.720 -0.020 186.320 42.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 184.720 451.885 186.320 489.620 ;
    END
    PORT
      LAYER met4 ;
        RECT 364.720 -0.020 366.320 42.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 364.720 451.885 366.320 489.620 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 177.080 455.260 178.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 344.080 455.260 345.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 15.300 26.960 16.900 459.920 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -5.380 -0.020 -3.780 489.620 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 -0.020 455.260 1.580 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 488.020 455.260 489.620 ;
    END
    PORT
      LAYER met4 ;
        RECT 453.660 -0.020 455.260 489.620 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.020 -0.020 189.620 42.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.020 451.885 189.620 489.620 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.020 -0.020 369.620 42.795 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.020 451.885 369.620 489.620 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 180.380 455.260 181.980 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 347.380 455.260 348.980 ;
    END
    PORT
      LAYER met4 ;
        RECT 18.980 26.960 20.580 459.920 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 444.550 478.805 ;
      LAYER li1 ;
        RECT 5.520 10.795 444.360 478.805 ;
      LAYER met1 ;
        RECT 4.210 10.640 447.970 478.960 ;
      LAYER met2 ;
        RECT 4.230 485.720 41.670 486.725 ;
        RECT 42.510 485.720 73.870 486.725 ;
        RECT 74.710 485.720 77.090 486.725 ;
        RECT 77.930 485.720 83.530 486.725 ;
        RECT 84.370 485.720 89.970 486.725 ;
        RECT 90.810 485.720 96.410 486.725 ;
        RECT 97.250 485.720 99.630 486.725 ;
        RECT 100.470 485.720 106.070 486.725 ;
        RECT 106.910 485.720 112.510 486.725 ;
        RECT 113.350 485.720 115.730 486.725 ;
        RECT 116.570 485.720 122.170 486.725 ;
        RECT 123.010 485.720 128.610 486.725 ;
        RECT 129.450 485.720 135.050 486.725 ;
        RECT 135.890 485.720 138.270 486.725 ;
        RECT 139.110 485.720 144.710 486.725 ;
        RECT 145.550 485.720 151.150 486.725 ;
        RECT 151.990 485.720 154.370 486.725 ;
        RECT 155.210 485.720 160.810 486.725 ;
        RECT 161.650 485.720 167.250 486.725 ;
        RECT 168.090 485.720 173.690 486.725 ;
        RECT 174.530 485.720 176.910 486.725 ;
        RECT 177.750 485.720 183.350 486.725 ;
        RECT 184.190 485.720 189.790 486.725 ;
        RECT 190.630 485.720 193.010 486.725 ;
        RECT 193.850 485.720 199.450 486.725 ;
        RECT 200.290 485.720 205.890 486.725 ;
        RECT 206.730 485.720 212.330 486.725 ;
        RECT 213.170 485.720 215.550 486.725 ;
        RECT 216.390 485.720 221.990 486.725 ;
        RECT 222.830 485.720 247.750 486.725 ;
        RECT 248.590 485.720 254.190 486.725 ;
        RECT 255.030 485.720 260.630 486.725 ;
        RECT 261.470 485.720 273.510 486.725 ;
        RECT 274.350 485.720 279.950 486.725 ;
        RECT 280.790 485.720 283.170 486.725 ;
        RECT 284.010 485.720 289.610 486.725 ;
        RECT 290.450 485.720 296.050 486.725 ;
        RECT 296.890 485.720 299.270 486.725 ;
        RECT 300.110 485.720 305.710 486.725 ;
        RECT 306.550 485.720 312.150 486.725 ;
        RECT 312.990 485.720 318.590 486.725 ;
        RECT 319.430 485.720 321.810 486.725 ;
        RECT 322.650 485.720 328.250 486.725 ;
        RECT 329.090 485.720 334.690 486.725 ;
        RECT 335.530 485.720 337.910 486.725 ;
        RECT 338.750 485.720 344.350 486.725 ;
        RECT 345.190 485.720 350.790 486.725 ;
        RECT 351.630 485.720 357.230 486.725 ;
        RECT 358.070 485.720 360.450 486.725 ;
        RECT 361.290 485.720 366.890 486.725 ;
        RECT 367.730 485.720 373.330 486.725 ;
        RECT 374.170 485.720 376.550 486.725 ;
        RECT 377.390 485.720 382.990 486.725 ;
        RECT 383.830 485.720 389.430 486.725 ;
        RECT 390.270 485.720 395.870 486.725 ;
        RECT 396.710 485.720 399.090 486.725 ;
        RECT 399.930 485.720 405.530 486.725 ;
        RECT 406.370 485.720 411.970 486.725 ;
        RECT 412.810 485.720 447.950 486.725 ;
        RECT 4.230 4.280 447.950 485.720 ;
        RECT 4.230 4.000 6.250 4.280 ;
        RECT 7.090 4.000 9.470 4.280 ;
        RECT 10.310 4.000 12.690 4.280 ;
        RECT 13.530 4.000 15.910 4.280 ;
        RECT 16.750 4.000 19.130 4.280 ;
        RECT 19.970 4.000 22.350 4.280 ;
        RECT 23.190 4.000 25.570 4.280 ;
        RECT 26.410 4.000 28.790 4.280 ;
        RECT 29.630 4.000 32.010 4.280 ;
        RECT 32.850 4.000 35.230 4.280 ;
        RECT 36.070 4.000 38.450 4.280 ;
        RECT 39.290 4.000 41.670 4.280 ;
        RECT 42.510 4.000 44.890 4.280 ;
        RECT 45.730 4.000 48.110 4.280 ;
        RECT 48.950 4.000 51.330 4.280 ;
        RECT 52.170 4.000 54.550 4.280 ;
        RECT 55.390 4.000 57.770 4.280 ;
        RECT 58.610 4.000 60.990 4.280 ;
        RECT 61.830 4.000 67.430 4.280 ;
        RECT 68.270 4.000 77.090 4.280 ;
        RECT 77.930 4.000 80.310 4.280 ;
        RECT 81.150 4.000 86.750 4.280 ;
        RECT 87.590 4.000 93.190 4.280 ;
        RECT 94.030 4.000 96.410 4.280 ;
        RECT 97.250 4.000 102.850 4.280 ;
        RECT 103.690 4.000 109.290 4.280 ;
        RECT 110.130 4.000 115.730 4.280 ;
        RECT 116.570 4.000 118.950 4.280 ;
        RECT 119.790 4.000 125.390 4.280 ;
        RECT 126.230 4.000 131.830 4.280 ;
        RECT 132.670 4.000 135.050 4.280 ;
        RECT 135.890 4.000 141.490 4.280 ;
        RECT 142.330 4.000 147.930 4.280 ;
        RECT 148.770 4.000 154.370 4.280 ;
        RECT 155.210 4.000 157.590 4.280 ;
        RECT 158.430 4.000 164.030 4.280 ;
        RECT 164.870 4.000 170.470 4.280 ;
        RECT 171.310 4.000 173.690 4.280 ;
        RECT 174.530 4.000 180.130 4.280 ;
        RECT 180.970 4.000 186.570 4.280 ;
        RECT 187.410 4.000 193.010 4.280 ;
        RECT 193.850 4.000 196.230 4.280 ;
        RECT 197.070 4.000 202.670 4.280 ;
        RECT 203.510 4.000 209.110 4.280 ;
        RECT 209.950 4.000 212.330 4.280 ;
        RECT 213.170 4.000 218.770 4.280 ;
        RECT 219.610 4.000 225.210 4.280 ;
        RECT 226.050 4.000 276.730 4.280 ;
        RECT 277.570 4.000 279.950 4.280 ;
        RECT 280.790 4.000 286.390 4.280 ;
        RECT 287.230 4.000 292.830 4.280 ;
        RECT 293.670 4.000 299.270 4.280 ;
        RECT 300.110 4.000 302.490 4.280 ;
        RECT 303.330 4.000 308.930 4.280 ;
        RECT 309.770 4.000 315.370 4.280 ;
        RECT 316.210 4.000 318.590 4.280 ;
        RECT 319.430 4.000 325.030 4.280 ;
        RECT 325.870 4.000 331.470 4.280 ;
        RECT 332.310 4.000 337.910 4.280 ;
        RECT 338.750 4.000 341.130 4.280 ;
        RECT 341.970 4.000 347.570 4.280 ;
        RECT 348.410 4.000 354.010 4.280 ;
        RECT 354.850 4.000 357.230 4.280 ;
        RECT 358.070 4.000 363.670 4.280 ;
        RECT 364.510 4.000 370.110 4.280 ;
        RECT 370.950 4.000 376.550 4.280 ;
        RECT 377.390 4.000 379.770 4.280 ;
        RECT 380.610 4.000 386.210 4.280 ;
        RECT 387.050 4.000 392.650 4.280 ;
        RECT 393.490 4.000 395.870 4.280 ;
        RECT 396.710 4.000 402.310 4.280 ;
        RECT 403.150 4.000 408.750 4.280 ;
        RECT 409.590 4.000 415.190 4.280 ;
        RECT 416.030 4.000 447.950 4.280 ;
      LAYER met3 ;
        RECT 3.950 446.440 447.975 486.705 ;
        RECT 3.950 445.040 445.600 446.440 ;
        RECT 3.950 443.040 447.975 445.040 ;
        RECT 3.950 441.640 445.600 443.040 ;
        RECT 3.950 439.640 447.975 441.640 ;
        RECT 3.950 438.240 445.600 439.640 ;
        RECT 3.950 432.840 447.975 438.240 ;
        RECT 4.400 431.440 445.600 432.840 ;
        RECT 3.950 426.040 447.975 431.440 ;
        RECT 4.400 424.640 445.600 426.040 ;
        RECT 3.950 419.240 447.975 424.640 ;
        RECT 4.400 417.840 445.600 419.240 ;
        RECT 3.950 412.440 447.975 417.840 ;
        RECT 4.400 411.040 445.600 412.440 ;
        RECT 3.950 405.640 447.975 411.040 ;
        RECT 4.400 404.240 445.600 405.640 ;
        RECT 3.950 398.840 447.975 404.240 ;
        RECT 4.400 397.440 445.600 398.840 ;
        RECT 3.950 392.040 447.975 397.440 ;
        RECT 4.400 390.640 445.600 392.040 ;
        RECT 3.950 385.240 447.975 390.640 ;
        RECT 4.400 383.840 445.600 385.240 ;
        RECT 3.950 378.440 447.975 383.840 ;
        RECT 4.400 377.040 445.600 378.440 ;
        RECT 3.950 371.640 447.975 377.040 ;
        RECT 4.400 370.240 445.600 371.640 ;
        RECT 3.950 364.840 447.975 370.240 ;
        RECT 4.400 363.440 445.600 364.840 ;
        RECT 3.950 358.040 447.975 363.440 ;
        RECT 4.400 356.640 445.600 358.040 ;
        RECT 3.950 351.240 447.975 356.640 ;
        RECT 4.400 349.840 445.600 351.240 ;
        RECT 3.950 344.440 447.975 349.840 ;
        RECT 4.400 343.040 445.600 344.440 ;
        RECT 3.950 337.640 447.975 343.040 ;
        RECT 4.400 336.240 445.600 337.640 ;
        RECT 3.950 330.840 447.975 336.240 ;
        RECT 4.400 329.440 445.600 330.840 ;
        RECT 3.950 324.040 447.975 329.440 ;
        RECT 4.400 322.640 445.600 324.040 ;
        RECT 3.950 317.240 447.975 322.640 ;
        RECT 4.400 315.840 445.600 317.240 ;
        RECT 3.950 310.440 447.975 315.840 ;
        RECT 4.400 309.040 445.600 310.440 ;
        RECT 3.950 307.040 447.975 309.040 ;
        RECT 4.400 305.640 447.975 307.040 ;
        RECT 3.950 303.640 447.975 305.640 ;
        RECT 4.400 302.240 445.600 303.640 ;
        RECT 3.950 300.240 447.975 302.240 ;
        RECT 4.400 298.840 447.975 300.240 ;
        RECT 3.950 296.840 447.975 298.840 ;
        RECT 4.400 295.440 445.600 296.840 ;
        RECT 3.950 293.440 447.975 295.440 ;
        RECT 4.400 292.040 447.975 293.440 ;
        RECT 3.950 290.040 447.975 292.040 ;
        RECT 4.400 288.640 445.600 290.040 ;
        RECT 3.950 286.640 447.975 288.640 ;
        RECT 4.400 285.240 447.975 286.640 ;
        RECT 3.950 283.240 447.975 285.240 ;
        RECT 4.400 281.840 445.600 283.240 ;
        RECT 3.950 279.840 447.975 281.840 ;
        RECT 4.400 278.440 447.975 279.840 ;
        RECT 3.950 276.440 447.975 278.440 ;
        RECT 4.400 275.040 445.600 276.440 ;
        RECT 3.950 273.040 447.975 275.040 ;
        RECT 4.400 271.640 447.975 273.040 ;
        RECT 3.950 269.640 447.975 271.640 ;
        RECT 4.400 268.240 445.600 269.640 ;
        RECT 3.950 266.240 447.975 268.240 ;
        RECT 4.400 264.840 447.975 266.240 ;
        RECT 3.950 262.840 447.975 264.840 ;
        RECT 4.400 261.440 445.600 262.840 ;
        RECT 3.950 259.440 447.975 261.440 ;
        RECT 4.400 258.040 447.975 259.440 ;
        RECT 3.950 256.040 447.975 258.040 ;
        RECT 4.400 254.640 445.600 256.040 ;
        RECT 3.950 252.640 447.975 254.640 ;
        RECT 4.400 251.240 445.600 252.640 ;
        RECT 3.950 249.240 447.975 251.240 ;
        RECT 4.400 247.840 447.975 249.240 ;
        RECT 3.950 245.840 447.975 247.840 ;
        RECT 4.400 244.440 447.975 245.840 ;
        RECT 3.950 242.440 447.975 244.440 ;
        RECT 4.400 241.040 447.975 242.440 ;
        RECT 3.950 239.040 447.975 241.040 ;
        RECT 4.400 237.640 447.975 239.040 ;
        RECT 3.950 235.640 447.975 237.640 ;
        RECT 4.400 234.240 447.975 235.640 ;
        RECT 3.950 232.240 447.975 234.240 ;
        RECT 4.400 230.840 447.975 232.240 ;
        RECT 3.950 228.840 447.975 230.840 ;
        RECT 4.400 227.440 445.600 228.840 ;
        RECT 3.950 225.440 447.975 227.440 ;
        RECT 4.400 224.040 447.975 225.440 ;
        RECT 3.950 222.040 447.975 224.040 ;
        RECT 4.400 220.640 445.600 222.040 ;
        RECT 3.950 218.640 447.975 220.640 ;
        RECT 4.400 217.240 447.975 218.640 ;
        RECT 3.950 215.240 447.975 217.240 ;
        RECT 4.400 213.840 445.600 215.240 ;
        RECT 3.950 208.440 447.975 213.840 ;
        RECT 4.400 207.040 445.600 208.440 ;
        RECT 3.950 201.640 447.975 207.040 ;
        RECT 4.400 200.240 445.600 201.640 ;
        RECT 3.950 194.840 447.975 200.240 ;
        RECT 4.400 193.440 445.600 194.840 ;
        RECT 3.950 188.040 447.975 193.440 ;
        RECT 4.400 186.640 445.600 188.040 ;
        RECT 3.950 181.240 447.975 186.640 ;
        RECT 4.400 179.840 445.600 181.240 ;
        RECT 3.950 174.440 447.975 179.840 ;
        RECT 4.400 173.040 445.600 174.440 ;
        RECT 3.950 167.640 447.975 173.040 ;
        RECT 4.400 166.240 445.600 167.640 ;
        RECT 3.950 160.840 447.975 166.240 ;
        RECT 4.400 159.440 445.600 160.840 ;
        RECT 3.950 154.040 447.975 159.440 ;
        RECT 4.400 152.640 445.600 154.040 ;
        RECT 3.950 147.240 447.975 152.640 ;
        RECT 4.400 145.840 445.600 147.240 ;
        RECT 3.950 140.440 447.975 145.840 ;
        RECT 4.400 139.040 445.600 140.440 ;
        RECT 3.950 133.640 447.975 139.040 ;
        RECT 4.400 132.240 445.600 133.640 ;
        RECT 3.950 126.840 447.975 132.240 ;
        RECT 4.400 125.440 445.600 126.840 ;
        RECT 3.950 120.040 447.975 125.440 ;
        RECT 4.400 118.640 445.600 120.040 ;
        RECT 3.950 113.240 447.975 118.640 ;
        RECT 4.400 111.840 445.600 113.240 ;
        RECT 3.950 106.440 447.975 111.840 ;
        RECT 4.400 105.040 445.600 106.440 ;
        RECT 3.950 99.640 447.975 105.040 ;
        RECT 4.400 98.240 445.600 99.640 ;
        RECT 3.950 92.840 447.975 98.240 ;
        RECT 4.400 91.440 445.600 92.840 ;
        RECT 3.950 86.040 447.975 91.440 ;
        RECT 4.400 84.640 445.600 86.040 ;
        RECT 3.950 79.240 447.975 84.640 ;
        RECT 4.400 77.840 445.600 79.240 ;
        RECT 3.950 72.440 447.975 77.840 ;
        RECT 4.400 71.040 445.600 72.440 ;
        RECT 3.950 65.640 447.975 71.040 ;
        RECT 4.400 64.240 445.600 65.640 ;
        RECT 3.950 58.840 447.975 64.240 ;
        RECT 4.400 57.440 445.600 58.840 ;
        RECT 3.950 52.040 447.975 57.440 ;
        RECT 3.950 50.640 445.600 52.040 ;
        RECT 3.950 48.640 447.975 50.640 ;
        RECT 3.950 47.240 445.600 48.640 ;
        RECT 3.950 45.240 447.975 47.240 ;
        RECT 3.950 43.840 445.600 45.240 ;
        RECT 3.950 41.840 447.975 43.840 ;
        RECT 3.950 40.440 445.600 41.840 ;
        RECT 3.950 10.715 447.975 40.440 ;
      LAYER met4 ;
        RECT 3.975 460.320 184.320 476.505 ;
        RECT 3.975 26.560 14.900 460.320 ;
        RECT 17.300 26.560 18.580 460.320 ;
        RECT 20.980 451.485 184.320 460.320 ;
        RECT 186.720 451.485 187.620 476.505 ;
        RECT 190.020 451.485 364.320 476.505 ;
        RECT 366.720 451.485 367.620 476.505 ;
        RECT 370.020 451.485 446.825 476.505 ;
        RECT 20.980 43.195 446.825 451.485 ;
        RECT 20.980 26.560 184.320 43.195 ;
        RECT 3.975 22.615 184.320 26.560 ;
        RECT 186.720 22.615 187.620 43.195 ;
        RECT 190.020 22.615 364.320 43.195 ;
        RECT 366.720 22.615 367.620 43.195 ;
        RECT 370.020 22.615 446.825 43.195 ;
      LAYER met5 ;
        RECT 44.720 350.580 429.620 431.980 ;
        RECT 44.720 183.580 429.620 342.480 ;
        RECT 44.720 50.080 429.620 175.480 ;
  END
END fpga
END LIBRARY

