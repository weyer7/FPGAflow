* NGSPICE file created from matrix_mult.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

.subckt matrix_mult VGND VPWR bit_period[0] bit_period[10] bit_period[11] bit_period[12]
+ bit_period[13] bit_period[1] bit_period[2] bit_period[3] bit_period[4] bit_period[5]
+ bit_period[6] bit_period[7] bit_period[8] bit_period[9] clk confirmation data_read
+ n_rst serial_in serial_out tx_busy
XFILLER_39_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0985_ clknet_3_1__leaf_clk _0035_ net29 VGND VGND VPWR VPWR parallel_out1\[6\] sky130_fd_sc_hd__dfstp_1
XFILLER_42_217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_40 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0770_ parallel_out2\[0\] parallel_out2\[6\] parallel_out2\[1\] parallel_out2\[5\]
+ VGND VGND VPWR VPWR _0333_ sky130_fd_sc_hd__a22oi_1
XTAP_TAPCELL_ROW_11_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0968_ clknet_3_6__leaf_clk uart_rcv.tim.clock_count.next_cnt_out\[13\] net38 VGND
+ VGND VPWR VPWR uart_rcv.tim.clk_cnt\[13\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_34_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0899_ _0426_ _0429_ VGND VGND VPWR VPWR _0430_ sky130_fd_sc_hd__nand2_1
XFILLER_2_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0822_ _0063_ net15 _0167_ _0375_ VGND VGND VPWR VPWR _0378_ sky130_fd_sc_hd__o31a_1
X_0684_ _0256_ _0267_ _0257_ VGND VGND VPWR VPWR _0268_ sky130_fd_sc_hd__a21oi_1
X_0753_ rx_data\[6\] uart_rcv.data_buff.packet_data\[6\] _0321_ VGND VGND VPWR VPWR
+ _0011_ sky130_fd_sc_hd__mux2_1
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1021_ clknet_3_7__leaf_clk uart_tx.count.next_cnt_out\[9\] net39 VGND VGND VPWR
+ VPWR uart_tx.clk_cnt\[9\] sky130_fd_sc_hd__dfrtp_1
X_0805_ parallel_out2\[7\] parallel_out2\[2\] parallel_out2\[6\] parallel_out2\[3\]
+ VGND VGND VPWR VPWR _0365_ sky130_fd_sc_hd__a22o_1
X_0667_ _0248_ _0249_ VGND VGND VPWR VPWR _0251_ sky130_fd_sc_hd__nor2_1
X_0736_ _0313_ _0315_ VGND VGND VPWR VPWR uart_rcv.control.next_state\[2\] sky130_fd_sc_hd__or2_1
X_0598_ _0070_ uart_tx.clk_cnt\[12\] _0186_ _0188_ _0190_ VGND VGND VPWR VPWR _0197_
+ sky130_fd_sc_hd__a2111o_1
XFILLER_29_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0452_ net45 VGND VGND VPWR VPWR _0072_ sky130_fd_sc_hd__inv_2
X_0521_ uart_rcv.tim.clk_cnt\[4\] uart_rcv.tim.clk_cnt\[5\] uart_rcv.tim.clk_cnt\[6\]
+ _0124_ VGND VGND VPWR VPWR _0130_ sky130_fd_sc_hd__and4_1
XFILLER_13_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1004_ clknet_3_2__leaf_clk _0054_ net31 VGND VGND VPWR VPWR uart_rcv.data_buff.packet_data\[1\]
+ sky130_fd_sc_hd__dfstp_1
X_0719_ _0258_ _0259_ VGND VGND VPWR VPWR _0302_ sky130_fd_sc_hd__nand2_1
XFILLER_17_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0504_ _0115_ _0117_ _0118_ uart_rcv.control.packet_done VGND VGND VPWR VPWR uart_rcv.tim.clock_count.next_cnt_out\[0\]
+ sky130_fd_sc_hd__a211oi_1
XTAP_TAPCELL_ROW_17_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_6__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_6__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_9_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0984_ clknet_3_1__leaf_clk _0034_ net29 VGND VGND VPWR VPWR parallel_out1\[5\] sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_6_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_28_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0967_ clknet_3_6__leaf_clk uart_rcv.tim.clock_count.next_cnt_out\[12\] net38 VGND
+ VGND VPWR VPWR uart_rcv.tim.clk_cnt\[12\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0898_ _0427_ _0428_ VGND VGND VPWR VPWR _0429_ sky130_fd_sc_hd__xnor2_1
XFILLER_15_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0821_ _0080_ _0323_ _0376_ _0063_ VGND VGND VPWR VPWR _0377_ sky130_fd_sc_hd__a22o_1
X_0752_ rx_data\[5\] uart_rcv.data_buff.packet_data\[5\] _0321_ VGND VGND VPWR VPWR
+ _0010_ sky130_fd_sc_hd__mux2_1
XFILLER_43_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0683_ prod_adder.gen_for_loop\[3\].adder_n.b _0265_ _0266_ VGND VGND VPWR VPWR _0267_
+ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_0_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmatrix_mult_40 VGND VGND VPWR VPWR matrix_mult_40/HI tx_busy sky130_fd_sc_hd__conb_1
X_1020_ clknet_3_7__leaf_clk uart_tx.count.next_cnt_out\[8\] net37 VGND VGND VPWR
+ VPWR uart_tx.clk_cnt\[8\] sky130_fd_sc_hd__dfrtp_1
X_0804_ _0359_ _0363_ VGND VGND VPWR VPWR _0364_ sky130_fd_sc_hd__xnor2_1
X_0735_ uart_rcv.control.state\[2\] uart_rcv.control.state\[0\] uart_rcv.control.state\[1\]
+ VGND VGND VPWR VPWR _0315_ sky130_fd_sc_hd__and3b_1
X_0666_ uart_tx.tx_ctrl.state\[0\] uart_tx.tx_ctrl.state\[1\] VGND VGND VPWR VPWR
+ _0250_ sky130_fd_sc_hd__or2_1
X_0597_ _0193_ _0194_ _0195_ VGND VGND VPWR VPWR _0196_ sky130_fd_sc_hd__or3b_1
XFILLER_43_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0451_ net5 VGND VGND VPWR VPWR _0071_ sky130_fd_sc_hd__inv_2
X_0520_ _0128_ _0129_ net21 VGND VGND VPWR VPWR uart_rcv.tim.clock_count.next_cnt_out\[5\]
+ sky130_fd_sc_hd__and3b_1
X_1003_ clknet_3_2__leaf_clk _0053_ net31 VGND VGND VPWR VPWR uart_rcv.data_buff.packet_data\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_34_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0718_ prod_adder.gen_for_loop\[0\].adder_n.b prod_adder.gen_for_loop\[0\].adder_n.a
+ _0296_ VGND VGND VPWR VPWR _0301_ sky130_fd_sc_hd__o21a_1
X_0649_ net9 uart_tx.count.next_cnt_out\[4\] VGND VGND VPWR VPWR _0234_ sky130_fd_sc_hd__xor2_1
XFILLER_40_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0503_ uart_rcv.tim.clk_cnt\[0\] _0116_ VGND VGND VPWR VPWR _0118_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_17_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0983_ clknet_3_1__leaf_clk _0033_ net29 VGND VGND VPWR VPWR parallel_out1\[4\] sky130_fd_sc_hd__dfstp_1
XFILLER_27_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_19_Left_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_34_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0966_ clknet_3_6__leaf_clk uart_rcv.tim.clock_count.next_cnt_out\[11\] net33 VGND
+ VGND VPWR VPWR uart_rcv.tim.clk_cnt\[11\] sky130_fd_sc_hd__dfrtp_1
X_0897_ _0416_ _0420_ _0417_ VGND VGND VPWR VPWR _0428_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_2_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_4_Left_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0820_ _0079_ _0080_ _0166_ VGND VGND VPWR VPWR _0376_ sky130_fd_sc_hd__and3_1
X_0751_ rx_data\[4\] uart_rcv.data_buff.packet_data\[4\] _0321_ VGND VGND VPWR VPWR
+ _0009_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0682_ _0263_ _0264_ prod_adder.gen_for_loop\[3\].adder_n.a VGND VGND VPWR VPWR _0266_
+ sky130_fd_sc_hd__a21o_1
XFILLER_36_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0949_ clknet_3_5__leaf_clk _0022_ net35 VGND VGND VPWR VPWR prod_adder.gen_for_loop\[7\].adder_n.b
+ sky130_fd_sc_hd__dfstp_1
XFILLER_7_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0803_ _0351_ _0353_ _0352_ VGND VGND VPWR VPWR _0363_ sky130_fd_sc_hd__o21bai_1
X_0665_ uart_tx.tx_ctrl.state\[0\] uart_tx.tx_ctrl.state\[1\] VGND VGND VPWR VPWR
+ _0249_ sky130_fd_sc_hd__nor2_1
X_0734_ uart_rcv.control.packet_done _0116_ _0313_ _0314_ VGND VGND VPWR VPWR uart_rcv.control.next_state\[0\]
+ sky130_fd_sc_hd__a211o_1
X_0596_ _0071_ uart_tx.clk_cnt\[13\] _0179_ _0189_ _0191_ VGND VGND VPWR VPWR _0195_
+ sky130_fd_sc_hd__o2111a_1
Xhold10 uart_rcv.shift_strobe VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_7_Left_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0450_ net4 VGND VGND VPWR VPWR _0070_ sky130_fd_sc_hd__inv_2
X_1002_ clknet_3_4__leaf_clk _0052_ net35 VGND VGND VPWR VPWR prod_adder.gen_for_loop\[7\].adder_n.a
+ sky130_fd_sc_hd__dfstp_1
XFILLER_34_111 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0717_ _0251_ _0273_ _0287_ _0297_ _0003_ VGND VGND VPWR VPWR _0300_ sky130_fd_sc_hd__a2111oi_1
X_0648_ _0064_ uart_tx.count.next_cnt_out\[3\] VGND VGND VPWR VPWR _0233_ sky130_fd_sc_hd__xnor2_1
X_0579_ uart_tx.clk_cnt\[12\] net4 VGND VGND VPWR VPWR _0178_ sky130_fd_sc_hd__and2b_1
XFILLER_15_89 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_33_Left_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0502_ uart_rcv.control.state\[0\] uart_rcv.control.state\[2\] uart_rcv.tim.clk_cnt\[0\]
+ uart_rcv.control.state\[1\] VGND VGND VPWR VPWR _0117_ sky130_fd_sc_hd__and4bb_1
XTAP_TAPCELL_ROW_17_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0982_ clknet_3_1__leaf_clk _0032_ net29 VGND VGND VPWR VPWR parallel_out1\[3\] sky130_fd_sc_hd__dfstp_1
XFILLER_27_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_36_Left_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_20_Left_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0896_ parallel_out1\[2\] parallel_out1\[5\] _0413_ _0412_ VGND VGND VPWR VPWR _0427_
+ sky130_fd_sc_hd__a31o_1
X_0965_ clknet_3_6__leaf_clk uart_rcv.tim.clock_count.next_cnt_out\[10\] net38 VGND
+ VGND VPWR VPWR uart_rcv.tim.clk_cnt\[10\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_2_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0750_ rx_data\[3\] uart_rcv.data_buff.packet_data\[3\] _0321_ VGND VGND VPWR VPWR
+ _0008_ sky130_fd_sc_hd__mux2_1
X_0681_ prod_adder.gen_for_loop\[3\].adder_n.a _0263_ _0264_ VGND VGND VPWR VPWR _0265_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_0_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0948_ clknet_3_4__leaf_clk _0021_ net35 VGND VGND VPWR VPWR prod_adder.gen_for_loop\[6\].adder_n.b
+ sky130_fd_sc_hd__dfstp_1
X_0879_ parallel_out1\[2\] parallel_out1\[5\] VGND VGND VPWR VPWR _0411_ sky130_fd_sc_hd__nand2_1
XFILLER_7_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0802_ parallel_out2\[7\] parallel_out2\[3\] parallel_out2\[2\] parallel_out2\[6\]
+ VGND VGND VPWR VPWR _0362_ sky130_fd_sc_hd__and4_1
X_0664_ uart_tx.tx_ctrl.state\[0\] uart_tx.tx_ctrl.state\[1\] VGND VGND VPWR VPWR
+ _0248_ sky130_fd_sc_hd__and2_1
X_0733_ uart_rcv.control.state\[2\] uart_rcv.sbd.new_sample uart_rcv.sbd.old_sample
+ _0312_ VGND VGND VPWR VPWR _0314_ sky130_fd_sc_hd__and4bb_1
X_0595_ _0065_ uart_tx.clk_cnt\[6\] _0177_ _0184_ _0185_ VGND VGND VPWR VPWR _0194_
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_1_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold11 uart_rcv.tim.bit_count.next_cnt_out\[0\] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1001_ clknet_3_4__leaf_clk _0051_ net35 VGND VGND VPWR VPWR prod_adder.gen_for_loop\[6\].adder_n.a
+ sky130_fd_sc_hd__dfstp_1
XFILLER_34_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0578_ uart_tx.clk_cnt\[9\] net14 VGND VGND VPWR VPWR _0177_ sky130_fd_sc_hd__nand2b_1
X_0716_ _0281_ _0298_ _0299_ VGND VGND VPWR VPWR _0003_ sky130_fd_sc_hd__or3_1
X_0647_ net6 uart_tx.count.next_cnt_out\[1\] VGND VGND VPWR VPWR _0232_ sky130_fd_sc_hd__xor2_1
XFILLER_40_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0501_ uart_rcv.control.state\[0\] uart_rcv.control.state\[2\] uart_rcv.control.state\[1\]
+ VGND VGND VPWR VPWR _0116_ sky130_fd_sc_hd__nor3b_2
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_159 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_55 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0981_ clknet_3_1__leaf_clk _0031_ net28 VGND VGND VPWR VPWR parallel_out1\[2\] sky130_fd_sc_hd__dfstp_1
XFILLER_8_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0964_ clknet_3_3__leaf_clk uart_rcv.tim.clock_count.next_cnt_out\[9\] net33 VGND
+ VGND VPWR VPWR uart_rcv.tim.clk_cnt\[9\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_34_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0895_ _0422_ _0425_ VGND VGND VPWR VPWR _0426_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_2_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0680_ prod_adder.gen_for_loop\[2\].adder_n.a _0258_ _0261_ prod_adder.gen_for_loop\[2\].adder_n.b
+ VGND VGND VPWR VPWR _0264_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_0_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0947_ clknet_3_5__leaf_clk _0020_ net36 VGND VGND VPWR VPWR prod_adder.gen_for_loop\[5\].adder_n.b
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_30_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0878_ _0409_ _0410_ prod_adder.gen_for_loop\[2\].adder_n.a _0384_ VGND VGND VPWR
+ VPWR _0047_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_11_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload0 clknet_3_0__leaf_clk VGND VGND VPWR VPWR clkload0/Y sky130_fd_sc_hd__inv_4
X_0801_ _0361_ prod_adder.gen_for_loop\[4\].adder_n.b net22 VGND VGND VPWR VPWR _0019_
+ sky130_fd_sc_hd__mux2_1
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0663_ _0070_ uart_tx.count.next_cnt_out\[12\] _0243_ _0244_ _0247_ VGND VGND VPWR
+ VPWR uart_tx.count.next_roflag sky130_fd_sc_hd__o2111a_1
XFILLER_6_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0732_ cntrl.framing_error _0312_ uart_rcv.control.state\[2\] VGND VGND VPWR VPWR
+ _0313_ sky130_fd_sc_hd__and3b_1
X_0594_ _0065_ uart_tx.clk_cnt\[6\] _0180_ _0181_ _0187_ VGND VGND VPWR VPWR _0193_
+ sky130_fd_sc_hd__a2111o_1
XFILLER_37_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold12 uart_rcv.tim.bit_cnt\[2\] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1000_ clknet_3_4__leaf_clk _0050_ net35 VGND VGND VPWR VPWR prod_adder.gen_for_loop\[5\].adder_n.a
+ sky130_fd_sc_hd__dfstp_1
X_0715_ _0248_ _0277_ VGND VGND VPWR VPWR _0299_ sky130_fd_sc_hd__and2b_1
X_0577_ net1 uart_tx.clk_cnt\[0\] VGND VGND VPWR VPWR _0176_ sky130_fd_sc_hd__and2b_1
X_0646_ net12 uart_tx.count.next_cnt_out\[7\] VGND VGND VPWR VPWR _0231_ sky130_fd_sc_hd__xor2_1
XFILLER_25_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0500_ _0109_ _0114_ VGND VGND VPWR VPWR _0115_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0629_ uart_tx.clk_cnt\[9\] _0218_ VGND VGND VPWR VPWR _0219_ sky130_fd_sc_hd__and2_1
XFILLER_26_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0980_ clknet_3_3__leaf_clk _0030_ net33 VGND VGND VPWR VPWR parallel_out1\[1\] sky130_fd_sc_hd__dfstp_1
XFILLER_8_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0894_ _0423_ _0424_ VGND VGND VPWR VPWR _0425_ sky130_fd_sc_hd__nor2_1
X_0963_ clknet_3_3__leaf_clk uart_rcv.tim.clock_count.next_cnt_out\[8\] net33 VGND
+ VGND VPWR VPWR uart_rcv.tim.clk_cnt\[8\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_2_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0946_ clknet_3_5__leaf_clk _0019_ net36 VGND VGND VPWR VPWR prod_adder.gen_for_loop\[4\].adder_n.b
+ sky130_fd_sc_hd__dfstp_1
X_0877_ _0401_ _0407_ _0408_ _0384_ VGND VGND VPWR VPWR _0410_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_30_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload1 clknet_3_2__leaf_clk VGND VGND VPWR VPWR clkload1/X sky130_fd_sc_hd__clkbuf_8
XFILLER_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0800_ _0359_ _0360_ VGND VGND VPWR VPWR _0361_ sky130_fd_sc_hd__and2_1
X_0731_ uart_rcv.control.state\[1\] uart_rcv.control.state\[0\] VGND VGND VPWR VPWR
+ _0312_ sky130_fd_sc_hd__nor2_1
X_0662_ net3 _0225_ _0229_ net5 _0246_ VGND VGND VPWR VPWR _0247_ sky130_fd_sc_hd__o221a_1
X_0593_ uart_tx.clk_cnt\[2\] net7 VGND VGND VPWR VPWR _0192_ sky130_fd_sc_hd__and2b_1
XFILLER_37_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0929_ clknet_3_3__leaf_clk _0005_ net32 VGND VGND VPWR VPWR rx_data\[0\] sky130_fd_sc_hd__dfstp_1
XFILLER_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold13 uart_tx.clk_cnt\[0\] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0645_ net14 uart_tx.count.next_cnt_out\[9\] VGND VGND VPWR VPWR _0230_ sky130_fd_sc_hd__xor2_1
X_0714_ uart_tx.tx_ctrl.state\[2\] _0248_ _0294_ VGND VGND VPWR VPWR _0298_ sky130_fd_sc_hd__and3_1
X_0576_ uart_tx.clk_cnt\[4\] net9 VGND VGND VPWR VPWR _0175_ sky130_fd_sc_hd__and2b_1
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0628_ _0218_ net20 _0217_ VGND VGND VPWR VPWR uart_tx.count.next_cnt_out\[8\] sky130_fd_sc_hd__and3b_1
XFILLER_7_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0559_ _0149_ _0151_ _0152_ _0156_ VGND VGND VPWR VPWR _0160_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_8_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0893_ parallel_out1\[2\] parallel_out1\[6\] parallel_out1\[1\] parallel_out1\[7\]
+ VGND VGND VPWR VPWR _0424_ sky130_fd_sc_hd__a22oi_1
X_0962_ clknet_3_6__leaf_clk uart_rcv.tim.clock_count.next_cnt_out\[7\] net38 VGND
+ VGND VPWR VPWR uart_rcv.tim.clk_cnt\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_24_Left_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0945_ clknet_3_5__leaf_clk _0018_ net36 VGND VGND VPWR VPWR prod_adder.gen_for_loop\[3\].adder_n.b
+ sky130_fd_sc_hd__dfstp_1
X_0876_ _0407_ _0408_ _0401_ VGND VGND VPWR VPWR _0409_ sky130_fd_sc_hd__a21oi_1
XFILLER_18_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload2 clknet_3_3__leaf_clk VGND VGND VPWR VPWR clkload2/Y sky130_fd_sc_hd__clkinv_2
X_0661_ net3 _0225_ _0245_ VGND VGND VPWR VPWR _0246_ sky130_fd_sc_hd__a21oi_1
XFILLER_6_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0730_ _0116_ _0311_ VGND VGND VPWR VPWR uart_rcv.control.next_state\[1\] sky130_fd_sc_hd__nand2b_1
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0592_ uart_tx.clk_cnt\[0\] net1 VGND VGND VPWR VPWR _0191_ sky130_fd_sc_hd__nand2b_1
XFILLER_37_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0859_ parallel_out2\[2\] rx_data\[2\] net23 VGND VGND VPWR VPWR _0039_ sky130_fd_sc_hd__mux2_1
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0928_ clknet_3_7__leaf_clk _0004_ net37 VGND VGND VPWR VPWR uart_tx.tx_ctrl.state\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold14 prod_adder.gen_for_loop\[1\].adder_n.a VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_134 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0644_ _0229_ VGND VGND VPWR VPWR uart_tx.count.next_cnt_out\[13\] sky130_fd_sc_hd__inv_2
X_0713_ uart_tx.tx_ctrl.state\[2\] _0251_ _0294_ _0296_ VGND VGND VPWR VPWR _0297_
+ sky130_fd_sc_hd__a31o_1
XPHY_EDGE_ROW_27_Left_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0575_ net5 uart_tx.clk_cnt\[13\] VGND VGND VPWR VPWR _0174_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_11_Left_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0627_ uart_tx.clk_cnt\[7\] uart_tx.clk_cnt\[8\] _0214_ VGND VGND VPWR VPWR _0218_
+ sky130_fd_sc_hd__and3_1
X_0558_ net14 uart_rcv.tim.clock_count.next_cnt_out\[9\] VGND VGND VPWR VPWR _0159_
+ sky130_fd_sc_hd__xor2_1
XFILLER_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0489_ net8 uart_rcv.tim.clk_cnt\[3\] VGND VGND VPWR VPWR _0104_ sky130_fd_sc_hd__and2b_1
XFILLER_21_151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_235 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0961_ clknet_3_3__leaf_clk uart_rcv.tim.clock_count.next_cnt_out\[6\] net32 VGND
+ VGND VPWR VPWR uart_rcv.tim.clk_cnt\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_32_224 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0892_ parallel_out1\[7\] parallel_out1\[2\] parallel_out1\[6\] parallel_out1\[1\]
+ VGND VGND VPWR VPWR _0423_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_25_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_7__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_7__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_0944_ clknet_3_4__leaf_clk _0017_ net35 VGND VGND VPWR VPWR prod_adder.gen_for_loop\[2\].adder_n.b
+ sky130_fd_sc_hd__dfstp_1
X_0875_ _0405_ _0406_ _0404_ VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_41_Left_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload3 clknet_3_4__leaf_clk VGND VGND VPWR VPWR clkload3/Y sky130_fd_sc_hd__clkinv_4
X_0660_ _0068_ uart_tx.count.next_cnt_out\[10\] VGND VGND VPWR VPWR _0245_ sky130_fd_sc_hd__xnor2_1
XFILLER_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0591_ uart_tx.clk_cnt\[5\] net10 VGND VGND VPWR VPWR _0190_ sky130_fd_sc_hd__and2b_1
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0927_ clknet_3_5__leaf_clk _0003_ net36 VGND VGND VPWR VPWR uart_tx.tx_ctrl.state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_0789_ prod_adder.gen_for_loop\[3\].adder_n.b net22 _0349_ _0350_ VGND VGND VPWR
+ VPWR _0018_ sky130_fd_sc_hd__a22o_1
X_0858_ parallel_out2\[1\] rx_data\[1\] net23 VGND VGND VPWR VPWR _0038_ sky130_fd_sc_hd__mux2_1
XFILLER_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold15 uart_rcv.tim.bit_cnt\[1\] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0643_ uart_tx.clk_cnt\[13\] _0226_ _0228_ VGND VGND VPWR VPWR _0229_ sky130_fd_sc_hd__a21o_1
X_0712_ uart_tx.tx_ctrl.state\[2\] _0250_ _0295_ VGND VGND VPWR VPWR _0296_ sky130_fd_sc_hd__a21oi_1
X_0574_ uart_tx.clk_cnt\[8\] net13 VGND VGND VPWR VPWR _0173_ sky130_fd_sc_hd__and2b_1
XFILLER_0_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0557_ _0148_ _0150_ _0157_ _0155_ VGND VGND VPWR VPWR _0158_ sky130_fd_sc_hd__or4b_1
X_0626_ uart_tx.clk_cnt\[7\] _0214_ uart_tx.clk_cnt\[8\] VGND VGND VPWR VPWR _0217_
+ sky130_fd_sc_hd__a21o_1
X_0488_ uart_rcv.tim.clk_cnt\[9\] net14 VGND VGND VPWR VPWR _0103_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0609_ uart_tx.clk_cnt\[0\] uart_tx.clk_cnt\[1\] uart_tx.clk_cnt\[2\] VGND VGND VPWR
+ VPWR _0206_ sky130_fd_sc_hd__a21o_1
XFILLER_41_247 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_244 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0960_ clknet_3_3__leaf_clk uart_rcv.tim.clock_count.next_cnt_out\[5\] net30 VGND
+ VGND VPWR VPWR uart_rcv.tim.clk_cnt\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_32_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0891_ parallel_out1\[3\] parallel_out1\[5\] VGND VGND VPWR VPWR _0422_ sky130_fd_sc_hd__nand2_1
XFILLER_4_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0943_ clknet_3_4__leaf_clk _0016_ net35 VGND VGND VPWR VPWR prod_adder.gen_for_loop\[1\].adder_n.b
+ sky130_fd_sc_hd__dfstp_1
X_0874_ _0404_ _0405_ _0406_ VGND VGND VPWR VPWR _0407_ sky130_fd_sc_hd__or3_1
XFILLER_11_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload4 clknet_3_5__leaf_clk VGND VGND VPWR VPWR clkload4/Y sky130_fd_sc_hd__inv_8
X_0590_ net9 uart_tx.clk_cnt\[4\] VGND VGND VPWR VPWR _0189_ sky130_fd_sc_hd__nand2b_1
XFILLER_37_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0857_ parallel_out2\[0\] rx_data\[0\] net23 VGND VGND VPWR VPWR _0037_ sky130_fd_sc_hd__mux2_1
XFILLER_20_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0926_ clknet_3_5__leaf_clk _0002_ net36 VGND VGND VPWR VPWR uart_tx.tx_ctrl.state\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_0788_ _0346_ _0348_ net22 VGND VGND VPWR VPWR _0350_ sky130_fd_sc_hd__a21oi_1
Xhold16 cntrl.state\[0\] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_3_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0711_ uart_tx.tx_ctrl.state\[2\] _0248_ _0294_ VGND VGND VPWR VPWR _0295_ sky130_fd_sc_hd__o21ai_1
X_0642_ uart_tx.clk_cnt\[13\] _0226_ net20 VGND VGND VPWR VPWR _0228_ sky130_fd_sc_hd__o21ai_1
X_0573_ uart_tx.clk_cnt\[10\] net2 VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__and2b_1
XFILLER_25_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0909_ prod_adder.gen_for_loop\[5\].adder_n.a _0438_ _0383_ VGND VGND VPWR VPWR _0050_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0625_ uart_tx.clk_cnt\[7\] _0214_ _0216_ net20 VGND VGND VPWR VPWR uart_tx.count.next_cnt_out\[7\]
+ sky130_fd_sc_hd__o211a_1
X_0556_ net6 uart_rcv.tim.clock_count.next_cnt_out\[1\] VGND VGND VPWR VPWR _0157_
+ sky130_fd_sc_hd__xor2_1
X_0487_ uart_rcv.tim.clk_cnt\[2\] net7 VGND VGND VPWR VPWR _0102_ sky130_fd_sc_hd__and2b_1
XFILLER_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0608_ net20 _0204_ _0205_ VGND VGND VPWR VPWR uart_tx.count.next_cnt_out\[1\] sky130_fd_sc_hd__and3_1
X_0539_ uart_rcv.tim.clk_cnt\[11\] _0140_ net21 VGND VGND VPWR VPWR _0143_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_5_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0890_ prod_adder.gen_for_loop\[3\].adder_n.a _0421_ _0383_ VGND VGND VPWR VPWR _0048_
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout30 net31 VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_4
XFILLER_13_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0942_ clknet_3_4__leaf_clk _0015_ net35 VGND VGND VPWR VPWR prod_adder.gen_for_loop\[0\].adder_n.b
+ sky130_fd_sc_hd__dfstp_1
X_0873_ parallel_out1\[0\] parallel_out1\[6\] parallel_out1\[1\] parallel_out1\[5\]
+ VGND VGND VPWR VPWR _0406_ sky130_fd_sc_hd__a22oi_1
XFILLER_34_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload5 clknet_3_6__leaf_clk VGND VGND VPWR VPWR clkload5/Y sky130_fd_sc_hd__inv_6
XFILLER_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0787_ _0346_ _0348_ VGND VGND VPWR VPWR _0349_ sky130_fd_sc_hd__or2_1
X_0856_ parallel_out1\[7\] rx_data\[7\] _0083_ VGND VGND VPWR VPWR _0036_ sky130_fd_sc_hd__mux2_1
X_0925_ clknet_3_5__leaf_clk _0001_ net37 VGND VGND VPWR VPWR uart_tx.tx_ctrl.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_43_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0641_ _0226_ _0227_ VGND VGND VPWR VPWR uart_tx.count.next_cnt_out\[12\] sky130_fd_sc_hd__nor2_1
X_0710_ uart_tx.tx_ctrl.state\[4\] uart_tx.tx_ctrl.state\[3\] VGND VGND VPWR VPWR
+ _0294_ sky130_fd_sc_hd__nor2_1
X_0572_ _0167_ _0170_ VGND VGND VPWR VPWR _0171_ sky130_fd_sc_hd__and2b_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_140 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0839_ cntrl.overrun_error cntrl.framing_error _0373_ VGND VGND VPWR VPWR _0394_
+ sky130_fd_sc_hd__o21ai_1
X_0908_ _0435_ _0437_ VGND VGND VPWR VPWR _0438_ sky130_fd_sc_hd__xnor2_1
Xoutput18 net18 VGND VGND VPWR VPWR data_read sky130_fd_sc_hd__buf_2
XFILLER_16_107 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_195 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_15_Left_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0624_ uart_tx.clk_cnt\[7\] _0214_ VGND VGND VPWR VPWR _0216_ sky130_fd_sc_hd__nand2_1
XFILLER_38_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0555_ _0065_ uart_rcv.tim.clock_count.next_cnt_out\[6\] VGND VGND VPWR VPWR _0156_
+ sky130_fd_sc_hd__xnor2_1
X_0486_ net1 uart_rcv.tim.clk_cnt\[0\] VGND VGND VPWR VPWR _0101_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_5_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0607_ uart_tx.clk_cnt\[0\] uart_tx.clk_cnt\[1\] VGND VGND VPWR VPWR _0205_ sky130_fd_sc_hd__or2_1
X_0538_ uart_rcv.tim.clk_cnt\[10\] uart_rcv.tim.clk_cnt\[11\] _0137_ VGND VGND VPWR
+ VPWR _0142_ sky130_fd_sc_hd__and3_1
XFILLER_37_28 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0469_ _0085_ _0086_ VGND VGND VPWR VPWR _0087_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_28_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_18_Left_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout31 net32 VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__clkbuf_4
Xfanout20 _0203_ VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_0_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0941_ clknet_3_0__leaf_clk _0014_ net27 VGND VGND VPWR VPWR cntrl.overrun_error
+ sky130_fd_sc_hd__dfrtp_1
X_0872_ parallel_out1\[0\] parallel_out1\[6\] parallel_out1\[1\] parallel_out1\[5\]
+ VGND VGND VPWR VPWR _0405_ sky130_fd_sc_hd__and4_1
Xclkload6 clknet_3_7__leaf_clk VGND VGND VPWR VPWR clkload6/Y sky130_fd_sc_hd__inv_6
XPHY_EDGE_ROW_3_Left_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0924_ clknet_3_5__leaf_clk _0000_ net37 VGND VGND VPWR VPWR uart_tx.tx_ctrl.state\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_0786_ _0343_ _0347_ VGND VGND VPWR VPWR _0348_ sky130_fd_sc_hd__or2_1
X_0855_ parallel_out1\[6\] rx_data\[6\] _0083_ VGND VGND VPWR VPWR _0035_ sky130_fd_sc_hd__mux2_1
XFILLER_3_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0640_ uart_tx.clk_cnt\[12\] _0223_ _0203_ VGND VGND VPWR VPWR _0227_ sky130_fd_sc_hd__o21ai_1
X_0571_ uart_tx.tx_ctrl.state\[0\] _0169_ VGND VGND VPWR VPWR _0170_ sky130_fd_sc_hd__nor2_1
XFILLER_33_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0907_ _0430_ _0436_ VGND VGND VPWR VPWR _0437_ sky130_fd_sc_hd__xnor2_1
X_0769_ parallel_out2\[0\] parallel_out2\[6\] parallel_out2\[1\] parallel_out2\[5\]
+ VGND VGND VPWR VPWR _0332_ sky130_fd_sc_hd__and4_1
X_0838_ _0388_ _0389_ _0392_ VGND VGND VPWR VPWR _0393_ sky130_fd_sc_hd__or3_1
Xoutput19 net19 VGND VGND VPWR VPWR serial_out sky130_fd_sc_hd__buf_2
XFILLER_16_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_6_Left_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_32 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0623_ _0214_ _0215_ _0203_ VGND VGND VPWR VPWR uart_tx.count.next_cnt_out\[6\] sky130_fd_sc_hd__and3b_1
X_0554_ net13 uart_rcv.tim.clock_count.next_cnt_out\[8\] VGND VGND VPWR VPWR _0155_
+ sky130_fd_sc_hd__xnor2_1
X_0485_ net6 uart_rcv.tim.clk_cnt\[1\] VGND VGND VPWR VPWR _0100_ sky130_fd_sc_hd__nand2b_1
XFILLER_38_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_188 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_244 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_22_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_32_Left_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0606_ uart_tx.clk_cnt\[0\] uart_tx.clk_cnt\[1\] VGND VGND VPWR VPWR _0204_ sky130_fd_sc_hd__nand2_1
X_0537_ _0141_ VGND VGND VPWR VPWR uart_rcv.tim.clock_count.next_cnt_out\[10\] sky130_fd_sc_hd__inv_2
X_0468_ cntrl.state\[3\] cntrl.state\[2\] VGND VGND VPWR VPWR _0086_ sky130_fd_sc_hd__nand2b_1
XFILLER_5_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_3_2__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_24_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout21 _0119_ VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_2
XFILLER_13_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout32 net34 VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_0_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0940_ clknet_3_0__leaf_clk _0013_ net26 VGND VGND VPWR VPWR cntrl.data_ready sky130_fd_sc_hd__dfrtp_1
XFILLER_20_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0871_ parallel_out1\[4\] parallel_out1\[2\] VGND VGND VPWR VPWR _0404_ sky130_fd_sc_hd__and2_1
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0854_ parallel_out1\[5\] rx_data\[5\] _0083_ VGND VGND VPWR VPWR _0034_ sky130_fd_sc_hd__mux2_1
X_0923_ uart_rcv.sbc.stop_bit net17 net25 VGND VGND VPWR VPWR _0061_ sky130_fd_sc_hd__mux2_1
X_0785_ parallel_out2\[4\] parallel_out2\[3\] _0342_ VGND VGND VPWR VPWR _0347_ sky130_fd_sc_hd__a21oi_1
XFILLER_3_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_96 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_194 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_84 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0570_ uart_tx.tx_ctrl.state\[4\] uart_tx.tx_ctrl.state\[1\] uart_tx.tx_ctrl.state\[2\]
+ uart_tx.tx_ctrl.state\[3\] VGND VGND VPWR VPWR _0169_ sky130_fd_sc_hd__or4_1
X_0837_ cntrl.state\[0\] _0168_ _0390_ _0391_ VGND VGND VPWR VPWR _0392_ sky130_fd_sc_hd__a211o_1
X_0906_ _0422_ _0424_ _0423_ VGND VGND VPWR VPWR _0436_ sky130_fd_sc_hd__o21bai_1
X_0768_ parallel_out2\[4\] parallel_out2\[2\] VGND VGND VPWR VPWR _0331_ sky130_fd_sc_hd__and2_1
X_0699_ prod_adder.gen_for_loop\[3\].adder_n.b _0266_ _0267_ _0282_ net24 VGND VGND
+ VPWR VPWR _0283_ sky130_fd_sc_hd__o221a_1
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0484_ uart_rcv.tim.clk_cnt\[7\] net12 VGND VGND VPWR VPWR _0099_ sky130_fd_sc_hd__and2b_1
XFILLER_7_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0622_ uart_tx.clk_cnt\[6\] _0212_ VGND VGND VPWR VPWR _0215_ sky130_fd_sc_hd__or2_1
X_0553_ net12 uart_rcv.tim.clock_count.next_cnt_out\[7\] VGND VGND VPWR VPWR _0154_
+ sky130_fd_sc_hd__xor2_1
XFILLER_38_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0467_ cntrl.state\[0\] _0084_ VGND VGND VPWR VPWR _0085_ sky130_fd_sc_hd__nand2_1
X_0536_ _0139_ _0140_ VGND VGND VPWR VPWR _0141_ sky130_fd_sc_hd__or2_1
X_0605_ _0196_ _0201_ _0171_ VGND VGND VPWR VPWR _0203_ sky130_fd_sc_hd__o21ba_1
X_1019_ clknet_3_7__leaf_clk uart_tx.count.next_cnt_out\[7\] net37 VGND VGND VPWR
+ VPWR uart_tx.clk_cnt\[7\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_36_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0519_ uart_rcv.tim.clk_cnt\[5\] _0126_ VGND VGND VPWR VPWR _0129_ sky130_fd_sc_hd__or2_1
Xfanout22 _0326_ VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__buf_2
XFILLER_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout33 net34 VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_24_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_40 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0870_ net54 _0384_ _0403_ VGND VGND VPWR VPWR _0046_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_30_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0999_ clknet_3_4__leaf_clk _0049_ net35 VGND VGND VPWR VPWR prod_adder.gen_for_loop\[4\].adder_n.a
+ sky130_fd_sc_hd__dfstp_1
XFILLER_39_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0853_ parallel_out1\[4\] rx_data\[4\] _0083_ VGND VGND VPWR VPWR _0033_ sky130_fd_sc_hd__mux2_1
X_0922_ uart_rcv.data_buff.packet_data\[7\] uart_rcv.sbc.stop_bit net25 VGND VGND
+ VPWR VPWR _0060_ sky130_fd_sc_hd__mux2_1
X_0784_ _0336_ _0345_ VGND VGND VPWR VPWR _0346_ sky130_fd_sc_hd__xnor2_1
Xinput1 bit_period[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_2
XFILLER_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_96 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0836_ _0079_ _0086_ VGND VGND VPWR VPWR _0391_ sky130_fd_sc_hd__nor2_1
X_0905_ _0433_ _0434_ VGND VGND VPWR VPWR _0435_ sky130_fd_sc_hd__nand2b_1
X_0767_ _0330_ prod_adder.gen_for_loop\[1\].adder_n.b net22 VGND VGND VPWR VPWR _0016_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0698_ prod_adder.gen_for_loop\[3\].adder_n.b _0265_ VGND VGND VPWR VPWR _0282_ sky130_fd_sc_hd__and2_1
XFILLER_15_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0621_ uart_tx.clk_cnt\[4\] uart_tx.clk_cnt\[5\] uart_tx.clk_cnt\[6\] _0208_ VGND
+ VGND VPWR VPWR _0214_ sky130_fd_sc_hd__and4_1
X_0552_ _0070_ uart_rcv.tim.clock_count.next_cnt_out\[12\] VGND VGND VPWR VPWR _0153_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0483_ uart_rcv.tim.clk_cnt\[10\] _0068_ _0066_ net13 VGND VGND VPWR VPWR _0098_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0819_ cntrl.data_ready cntrl.overrun_error cntrl.framing_error _0374_ VGND VGND
+ VPWR VPWR _0375_ sky130_fd_sc_hd__or4_1
XFILLER_29_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0604_ net53 _0202_ _0171_ VGND VGND VPWR VPWR uart_tx.count.next_cnt_out\[0\] sky130_fd_sc_hd__a21oi_1
X_0466_ cntrl.state\[1\] cntrl.state\[4\] VGND VGND VPWR VPWR _0084_ sky130_fd_sc_hd__nor2_1
X_0535_ uart_rcv.tim.clk_cnt\[10\] _0130_ _0138_ VGND VGND VPWR VPWR _0140_ sky130_fd_sc_hd__and3_1
X_1018_ clknet_3_7__leaf_clk uart_tx.count.next_cnt_out\[6\] net37 VGND VGND VPWR
+ VPWR uart_tx.clk_cnt\[6\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_36_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0518_ uart_rcv.tim.clk_cnt\[4\] uart_rcv.tim.clk_cnt\[5\] _0124_ VGND VGND VPWR
+ VPWR _0128_ sky130_fd_sc_hd__and3_1
X_0449_ net3 VGND VGND VPWR VPWR _0069_ sky130_fd_sc_hd__inv_2
Xfanout34 net16 VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_2
Xfanout23 _0087_ VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_24_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_52 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0998_ clknet_3_4__leaf_clk _0048_ net36 VGND VGND VPWR VPWR prod_adder.gen_for_loop\[3\].adder_n.a
+ sky130_fd_sc_hd__dfstp_1
XFILLER_10_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0921_ uart_rcv.data_buff.packet_data\[6\] uart_rcv.data_buff.packet_data\[7\] net25
+ VGND VGND VPWR VPWR _0059_ sky130_fd_sc_hd__mux2_1
X_0783_ _0331_ _0332_ _0333_ VGND VGND VPWR VPWR _0345_ sky130_fd_sc_hd__o21ba_1
X_0852_ parallel_out1\[3\] rx_data\[3\] _0083_ VGND VGND VPWR VPWR _0032_ sky130_fd_sc_hd__mux2_1
Xinput2 bit_period[10] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__buf_1
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0904_ parallel_out1\[7\] parallel_out1\[2\] parallel_out1\[6\] parallel_out1\[3\]
+ VGND VGND VPWR VPWR _0434_ sky130_fd_sc_hd__a22o_1
X_0835_ cntrl.state\[4\] _0325_ _0385_ VGND VGND VPWR VPWR _0390_ sky130_fd_sc_hd__o21ai_1
X_0766_ _0328_ _0329_ VGND VGND VPWR VPWR _0330_ sky130_fd_sc_hd__and2_1
X_0697_ uart_tx.tx_ctrl.state\[4\] uart_tx.tx_ctrl.state\[2\] uart_tx.tx_ctrl.state\[3\]
+ VGND VGND VPWR VPWR _0281_ sky130_fd_sc_hd__nor3b_1
XTAP_TAPCELL_ROW_19_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0620_ _0212_ _0213_ net20 VGND VGND VPWR VPWR uart_tx.count.next_cnt_out\[5\] sky130_fd_sc_hd__and3b_1
X_0551_ net1 uart_rcv.tim.clock_count.next_cnt_out\[0\] VGND VGND VPWR VPWR _0152_
+ sky130_fd_sc_hd__xor2_1
X_0482_ net5 uart_rcv.tim.clk_cnt\[13\] VGND VGND VPWR VPWR _0097_ sky130_fd_sc_hd__nand2b_1
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_8_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0818_ _0081_ _0085_ _0373_ VGND VGND VPWR VPWR _0374_ sky130_fd_sc_hd__o21ba_1
X_0749_ rx_data\[2\] uart_rcv.data_buff.packet_data\[2\] _0321_ VGND VGND VPWR VPWR
+ _0007_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_13_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0534_ uart_rcv.tim.clk_cnt\[10\] _0137_ net21 VGND VGND VPWR VPWR _0139_ sky130_fd_sc_hd__o21ai_1
X_0603_ _0196_ _0201_ VGND VGND VPWR VPWR _0202_ sky130_fd_sc_hd__or2_1
X_0465_ _0079_ _0082_ VGND VGND VPWR VPWR _0083_ sky130_fd_sc_hd__nor2_4
X_1017_ clknet_3_7__leaf_clk uart_tx.count.next_cnt_out\[5\] net37 VGND VGND VPWR
+ VPWR uart_tx.clk_cnt\[5\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_36_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0517_ _0126_ _0127_ VGND VGND VPWR VPWR uart_rcv.tim.clock_count.next_cnt_out\[4\]
+ sky130_fd_sc_hd__nor2_1
X_0448_ net2 VGND VGND VPWR VPWR _0068_ sky130_fd_sc_hd__inv_2
Xfanout35 net36 VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_4
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_242 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_30_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0997_ clknet_3_4__leaf_clk _0047_ net38 VGND VGND VPWR VPWR prod_adder.gen_for_loop\[2\].adder_n.a
+ sky130_fd_sc_hd__dfstp_1
XFILLER_10_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_39_Left_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0920_ uart_rcv.data_buff.packet_data\[5\] uart_rcv.data_buff.packet_data\[6\] net25
+ VGND VGND VPWR VPWR _0058_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_23_Left_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0782_ parallel_out2\[4\] parallel_out2\[3\] _0342_ VGND VGND VPWR VPWR _0344_ sky130_fd_sc_hd__nand3_1
X_0851_ parallel_out1\[2\] rx_data\[2\] _0083_ VGND VGND VPWR VPWR _0031_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput3 bit_period[11] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0834_ _0083_ _0377_ net23 _0374_ VGND VGND VPWR VPWR _0389_ sky130_fd_sc_hd__or4b_1
X_0903_ parallel_out1\[7\] parallel_out1\[3\] parallel_out1\[2\] parallel_out1\[6\]
+ VGND VGND VPWR VPWR _0433_ sky130_fd_sc_hd__and4_1
XFILLER_33_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0765_ parallel_out2\[4\] parallel_out2\[1\] parallel_out2\[5\] parallel_out2\[0\]
+ VGND VGND VPWR VPWR _0329_ sky130_fd_sc_hd__a22o_1
X_0696_ _0277_ _0279_ VGND VGND VPWR VPWR _0280_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_19_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0550_ net7 uart_rcv.tim.clock_count.next_cnt_out\[2\] VGND VGND VPWR VPWR _0151_
+ sky130_fd_sc_hd__xor2_1
X_0481_ uart_rcv.tim.clk_cnt\[0\] net1 VGND VGND VPWR VPWR _0096_ sky130_fd_sc_hd__nand2b_1
X_0817_ _0086_ _0372_ VGND VGND VPWR VPWR _0373_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_26_Left_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_10_Left_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0679_ _0258_ _0261_ prod_adder.gen_for_loop\[2\].adder_n.a VGND VGND VPWR VPWR _0263_
+ sky130_fd_sc_hd__a21o_1
X_0748_ rx_data\[1\] uart_rcv.data_buff.packet_data\[1\] _0321_ VGND VGND VPWR VPWR
+ _0006_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0464_ _0063_ _0080_ VGND VGND VPWR VPWR _0082_ sky130_fd_sc_hd__nand2_1
X_0533_ _0137_ net21 _0136_ VGND VGND VPWR VPWR uart_rcv.tim.clock_count.next_cnt_out\[9\]
+ sky130_fd_sc_hd__and3b_1
X_0602_ _0197_ _0198_ _0199_ _0200_ VGND VGND VPWR VPWR _0201_ sky130_fd_sc_hd__or4_1
X_1016_ clknet_3_7__leaf_clk uart_tx.count.next_cnt_out\[4\] net37 VGND VGND VPWR
+ VPWR uart_tx.clk_cnt\[4\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_36_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0447_ uart_rcv.tim.clk_cnt\[9\] VGND VGND VPWR VPWR _0067_ sky130_fd_sc_hd__inv_2
X_0516_ uart_rcv.tim.clk_cnt\[4\] _0124_ net21 VGND VGND VPWR VPWR _0127_ sky130_fd_sc_hd__o21ai_1
Xfanout25 uart_rcv.shift_strobe VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_4
Xfanout36 net39 VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__buf_2
XFILLER_22_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0996_ clknet_3_4__leaf_clk _0046_ net36 VGND VGND VPWR VPWR prod_adder.gen_for_loop\[1\].adder_n.a
+ sky130_fd_sc_hd__dfstp_1
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0850_ parallel_out1\[1\] rx_data\[1\] _0083_ VGND VGND VPWR VPWR _0030_ sky130_fd_sc_hd__mux2_1
X_0781_ parallel_out2\[4\] parallel_out2\[3\] _0342_ VGND VGND VPWR VPWR _0343_ sky130_fd_sc_hd__and3_1
Xinput4 bit_period[12] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_1
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0979_ clknet_3_3__leaf_clk _0029_ net33 VGND VGND VPWR VPWR parallel_out1\[0\] sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_40_Left_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0833_ _0063_ _0168_ _0323_ _0381_ VGND VGND VPWR VPWR _0388_ sky130_fd_sc_hd__a22o_1
X_0902_ prod_adder.gen_for_loop\[4\].adder_n.a _0432_ _0383_ VGND VGND VPWR VPWR _0049_
+ sky130_fd_sc_hd__mux2_1
X_0764_ parallel_out2\[1\] parallel_out2\[5\] _0327_ VGND VGND VPWR VPWR _0328_ sky130_fd_sc_hd__nand3_1
X_0695_ _0268_ _0278_ VGND VGND VPWR VPWR _0279_ sky130_fd_sc_hd__xnor2_1
XFILLER_15_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0480_ net10 uart_rcv.tim.clk_cnt\[5\] VGND VGND VPWR VPWR _0095_ sky130_fd_sc_hd__xnor2_1
X_0816_ _0063_ _0084_ VGND VGND VPWR VPWR _0372_ sky130_fd_sc_hd__nand2_1
X_0747_ rx_data\[0\] uart_rcv.data_buff.packet_data\[0\] _0321_ VGND VGND VPWR VPWR
+ _0005_ sky130_fd_sc_hd__mux2_1
X_0678_ prod_adder.gen_for_loop\[2\].adder_n.a _0258_ _0261_ VGND VGND VPWR VPWR _0262_
+ sky130_fd_sc_hd__and3_1
XFILLER_8_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0601_ _0068_ uart_tx.clk_cnt\[10\] _0176_ _0183_ _0192_ VGND VGND VPWR VPWR _0200_
+ sky130_fd_sc_hd__a2111o_1
X_0463_ cntrl.state\[3\] cntrl.state\[2\] VGND VGND VPWR VPWR _0081_ sky130_fd_sc_hd__or2_1
X_0532_ uart_rcv.tim.clk_cnt\[7\] uart_rcv.tim.clk_cnt\[8\] uart_rcv.tim.clk_cnt\[9\]
+ VGND VGND VPWR VPWR _0138_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_36_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1015_ clknet_3_6__leaf_clk uart_tx.count.next_cnt_out\[3\] net38 VGND VGND VPWR
+ VPWR uart_tx.clk_cnt\[3\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_4_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_244 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0446_ uart_rcv.tim.clk_cnt\[8\] VGND VGND VPWR VPWR _0066_ sky130_fd_sc_hd__inv_2
X_0515_ uart_rcv.tim.clk_cnt\[4\] _0124_ VGND VGND VPWR VPWR _0126_ sky130_fd_sc_hd__and2_1
Xfanout26 net34 VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_4
Xfanout37 net39 VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_4
XFILLER_13_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0995_ clknet_3_4__leaf_clk _0045_ net35 VGND VGND VPWR VPWR prod_adder.gen_for_loop\[0\].adder_n.a
+ sky130_fd_sc_hd__dfstp_1
XFILLER_6_218 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0780_ _0338_ _0341_ VGND VGND VPWR VPWR _0342_ sky130_fd_sc_hd__xnor2_1
Xinput5 bit_period[13] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_2
XFILLER_36_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0978_ clknet_3_0__leaf_clk _0028_ net26 VGND VGND VPWR VPWR cntrl.state\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_2_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0832_ _0379_ _0387_ VGND VGND VPWR VPWR _0024_ sky130_fd_sc_hd__xnor2_1
X_0763_ _0327_ prod_adder.gen_for_loop\[0\].adder_n.b _0326_ VGND VGND VPWR VPWR _0015_
+ sky130_fd_sc_hd__mux2_1
X_0901_ _0430_ _0431_ VGND VGND VPWR VPWR _0432_ sky130_fd_sc_hd__and2_1
X_0694_ _0253_ _0254_ VGND VGND VPWR VPWR _0278_ sky130_fd_sc_hd__nand2b_1
XFILLER_32_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_16_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_139 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0815_ cntrl.framing_error _0315_ _0371_ _0311_ VGND VGND VPWR VPWR _0023_ sky130_fd_sc_hd__o211a_1
X_0746_ uart_rcv.control.state\[1\] uart_rcv.control.state\[0\] uart_rcv.control.state\[2\]
+ VGND VGND VPWR VPWR _0321_ sky130_fd_sc_hd__and3b_4
X_0677_ prod_adder.gen_for_loop\[1\].adder_n.b prod_adder.gen_for_loop\[1\].adder_n.a
+ prod_adder.gen_for_loop\[0\].adder_n.b prod_adder.gen_for_loop\[0\].adder_n.a VGND
+ VGND VPWR VPWR _0261_ sky130_fd_sc_hd__a22o_1
XFILLER_43_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_194 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0531_ uart_rcv.tim.clk_cnt\[7\] uart_rcv.tim.clk_cnt\[8\] uart_rcv.tim.clk_cnt\[9\]
+ _0130_ VGND VGND VPWR VPWR _0137_ sky130_fd_sc_hd__and4_1
X_0600_ _0064_ uart_tx.clk_cnt\[3\] _0173_ _0175_ _0178_ VGND VGND VPWR VPWR _0199_
+ sky130_fd_sc_hd__a2111o_1
X_0462_ cntrl.state\[3\] cntrl.state\[2\] VGND VGND VPWR VPWR _0080_ sky130_fd_sc_hd__nor2_1
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1014_ clknet_3_6__leaf_clk uart_tx.count.next_cnt_out\[2\] net38 VGND VGND VPWR
+ VPWR uart_tx.clk_cnt\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_34_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0729_ uart_rcv.control.state\[1\] uart_rcv.control.state\[2\] uart_rcv.control.state\[0\]
+ VGND VGND VPWR VPWR _0311_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_4_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0514_ _0124_ _0125_ _0119_ VGND VGND VPWR VPWR uart_rcv.tim.clock_count.next_cnt_out\[3\]
+ sky130_fd_sc_hd__and3b_1
X_0445_ net11 VGND VGND VPWR VPWR _0065_ sky130_fd_sc_hd__inv_2
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout27 net34 VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_2
XFILLER_22_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout38 net39 VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_32_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0994_ clknet_3_1__leaf_clk _0044_ net28 VGND VGND VPWR VPWR parallel_out2\[7\] sky130_fd_sc_hd__dfstp_2
XFILLER_5_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_131 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput6 bit_period[1] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_2
XFILLER_36_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0977_ clknet_3_0__leaf_clk _0027_ net26 VGND VGND VPWR VPWR cntrl.state\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_42_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_3__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_2_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0900_ _0426_ _0429_ VGND VGND VPWR VPWR _0431_ sky130_fd_sc_hd__or2_1
XFILLER_25_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0762_ parallel_out2\[0\] parallel_out2\[4\] VGND VGND VPWR VPWR _0327_ sky130_fd_sc_hd__and2_1
X_0831_ _0380_ _0384_ _0386_ VGND VGND VPWR VPWR _0387_ sky130_fd_sc_hd__and3_1
X_0693_ uart_tx.tx_ctrl.state\[4\] uart_tx.tx_ctrl.state\[2\] uart_tx.tx_ctrl.state\[3\]
+ VGND VGND VPWR VPWR _0277_ sky130_fd_sc_hd__and3b_1
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap24 _0281_ VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__buf_1
XFILLER_30_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_16_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0814_ uart_rcv.sbc.stop_bit _0315_ VGND VGND VPWR VPWR _0371_ sky130_fd_sc_hd__nand2_1
X_0676_ prod_adder.gen_for_loop\[0\].adder_n.b prod_adder.gen_for_loop\[0\].adder_n.a
+ VGND VGND VPWR VPWR _0260_ sky130_fd_sc_hd__nand2_1
X_0745_ _0286_ uart_tx.tx_ctrl.state\[4\] _0319_ VGND VGND VPWR VPWR _0004_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_39_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0530_ uart_rcv.tim.clk_cnt\[9\] _0135_ VGND VGND VPWR VPWR _0136_ sky130_fd_sc_hd__or2_1
X_0461_ cntrl.state\[4\] cntrl.state\[1\] VGND VGND VPWR VPWR _0079_ sky130_fd_sc_hd__nand2b_2
XPHY_EDGE_ROW_14_Left_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1013_ clknet_3_6__leaf_clk uart_tx.count.next_cnt_out\[1\] net38 VGND VGND VPWR
+ VPWR uart_tx.clk_cnt\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_34_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0659_ net5 _0229_ VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_4_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0728_ _0251_ _0284_ _0310_ VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__a21o_1
XFILLER_27_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0513_ uart_rcv.tim.clk_cnt\[3\] _0122_ VGND VGND VPWR VPWR _0125_ sky130_fd_sc_hd__or2_1
X_0444_ net8 VGND VGND VPWR VPWR _0064_ sky130_fd_sc_hd__inv_2
Xfanout39 net16 VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__buf_2
Xfanout28 net34 VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_4
X_0993_ clknet_3_1__leaf_clk _0043_ net28 VGND VGND VPWR VPWR parallel_out2\[6\] sky130_fd_sc_hd__dfstp_1
XFILLER_8_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_143 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_17_Left_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput7 bit_period[2] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_2
X_0976_ clknet_3_1__leaf_clk _0026_ net26 VGND VGND VPWR VPWR cntrl.state\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_42_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_2_Left_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0830_ _0080_ _0382_ _0385_ _0082_ VGND VGND VPWR VPWR _0386_ sky130_fd_sc_hd__o211a_1
X_0761_ _0324_ _0325_ VGND VGND VPWR VPWR _0326_ sky130_fd_sc_hd__or2_1
X_0692_ _0271_ _0272_ VGND VGND VPWR VPWR _0276_ sky130_fd_sc_hd__xnor2_1
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0959_ clknet_3_3__leaf_clk uart_rcv.tim.clock_count.next_cnt_out\[4\] net30 VGND
+ VGND VPWR VPWR uart_rcv.tim.clk_cnt\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_23_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput10 bit_period[5] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_2
X_0813_ _0072_ net22 _0369_ _0370_ VGND VGND VPWR VPWR _0022_ sky130_fd_sc_hd__a22oi_1
XFILLER_14_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0675_ prod_adder.gen_for_loop\[1\].adder_n.b prod_adder.gen_for_loop\[1\].adder_n.a
+ VGND VGND VPWR VPWR _0259_ sky130_fd_sc_hd__nand2_1
X_0744_ _0320_ uart_tx.tx_ctrl.state\[2\] _0319_ VGND VGND VPWR VPWR _0002_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_39_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0460_ uart_rcv.tim.bit_cnt\[0\] net50 _0078_ VGND VGND VPWR VPWR uart_rcv.tim.bit_count.next_cnt_out\[0\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_21_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1012_ clknet_3_6__leaf_clk uart_tx.count.next_cnt_out\[0\] net37 VGND VGND VPWR
+ VPWR uart_tx.clk_cnt\[0\] sky130_fd_sc_hd__dfrtp_2
X_0727_ _0287_ _0288_ _0289_ _0309_ VGND VGND VPWR VPWR _0310_ sky130_fd_sc_hd__a31o_1
X_0658_ _0070_ uart_tx.count.next_cnt_out\[12\] _0230_ _0242_ VGND VGND VPWR VPWR
+ _0243_ sky130_fd_sc_hd__a211oi_1
X_0589_ uart_tx.clk_cnt\[11\] net3 VGND VGND VPWR VPWR _0188_ sky130_fd_sc_hd__and2b_1
XFILLER_25_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_31_Left_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0512_ uart_rcv.tim.clk_cnt\[1\] uart_rcv.tim.clk_cnt\[2\] uart_rcv.tim.clk_cnt\[3\]
+ _0117_ VGND VGND VPWR VPWR _0124_ sky130_fd_sc_hd__and4_1
XFILLER_3_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0443_ cntrl.state\[0\] VGND VGND VPWR VPWR _0063_ sky130_fd_sc_hd__inv_2
Xfanout29 net34 VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_2
XFILLER_13_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0992_ clknet_3_1__leaf_clk _0042_ net28 VGND VGND VPWR VPWR parallel_out2\[5\] sky130_fd_sc_hd__dfstp_2
XFILLER_39_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_95 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput8 bit_period[3] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_1
X_0975_ clknet_3_0__leaf_clk _0025_ net26 VGND VGND VPWR VPWR cntrl.state\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_19_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0760_ cntrl.state\[2\] cntrl.state\[3\] VGND VGND VPWR VPWR _0325_ sky130_fd_sc_hd__nand2b_1
X_0691_ _0274_ VGND VGND VPWR VPWR _0275_ sky130_fd_sc_hd__inv_2
XFILLER_2_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0958_ clknet_3_3__leaf_clk uart_rcv.tim.clock_count.next_cnt_out\[3\] net31 VGND
+ VGND VPWR VPWR uart_rcv.tim.clk_cnt\[3\] sky130_fd_sc_hd__dfrtp_1
X_0889_ _0418_ _0420_ VGND VGND VPWR VPWR _0421_ sky130_fd_sc_hd__xnor2_1
XFILLER_38_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput11 bit_period[6] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_1
X_0812_ _0368_ _0369_ _0370_ net22 net49 VGND VGND VPWR VPWR _0021_ sky130_fd_sc_hd__a32o_1
X_0743_ _0248_ _0275_ _0291_ _0297_ _0299_ VGND VGND VPWR VPWR _0320_ sky130_fd_sc_hd__a2111o_1
X_0674_ prod_adder.gen_for_loop\[1\].adder_n.b prod_adder.gen_for_loop\[1\].adder_n.a
+ VGND VGND VPWR VPWR _0258_ sky130_fd_sc_hd__or2_1
XFILLER_16_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_120 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1011_ clknet_3_2__leaf_clk _0061_ net30 VGND VGND VPWR VPWR uart_rcv.sbc.stop_bit
+ sky130_fd_sc_hd__dfstp_1
XFILLER_8_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0726_ _0290_ _0293_ _0304_ _0308_ VGND VGND VPWR VPWR _0309_ sky130_fd_sc_hd__a211o_1
X_0657_ _0231_ _0236_ _0241_ VGND VGND VPWR VPWR _0242_ sky130_fd_sc_hd__or3_1
X_0588_ uart_tx.clk_cnt\[7\] net12 VGND VGND VPWR VPWR _0187_ sky130_fd_sc_hd__and2b_1
XFILLER_43_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_38 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0511_ _0122_ _0123_ VGND VGND VPWR VPWR uart_rcv.tim.clock_count.next_cnt_out\[2\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_33_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0442_ uart_rcv.tim.bit_cnt\[3\] VGND VGND VPWR VPWR _0062_ sky130_fd_sc_hd__inv_2
XFILLER_3_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0709_ _0255_ _0257_ _0267_ _0292_ VGND VGND VPWR VPWR _0293_ sky130_fd_sc_hd__o31a_1
XFILLER_38_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0991_ clknet_3_1__leaf_clk _0041_ net28 VGND VGND VPWR VPWR parallel_out2\[4\] sky130_fd_sc_hd__dfstp_1
XFILLER_5_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput9 bit_period[4] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_1_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0974_ clknet_3_1__leaf_clk _0024_ net26 VGND VGND VPWR VPWR cntrl.state\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_27_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0690_ uart_tx.tx_ctrl.state\[4\] _0273_ VGND VGND VPWR VPWR _0274_ sky130_fd_sc_hd__nand2_1
XFILLER_2_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0957_ clknet_3_3__leaf_clk uart_rcv.tim.clock_count.next_cnt_out\[2\] net32 VGND
+ VGND VPWR VPWR uart_rcv.tim.clk_cnt\[2\] sky130_fd_sc_hd__dfrtp_1
X_0888_ _0409_ _0419_ VGND VGND VPWR VPWR _0420_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_16_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput12 bit_period[7] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_2
X_0811_ net22 _0362_ VGND VGND VPWR VPWR _0370_ sky130_fd_sc_hd__nor2_1
X_0673_ prod_adder.gen_for_loop\[4\].adder_n.b prod_adder.gen_for_loop\[4\].adder_n.a
+ VGND VGND VPWR VPWR _0257_ sky130_fd_sc_hd__nor2_1
X_0742_ _0316_ _0251_ VGND VGND VPWR VPWR _0001_ sky130_fd_sc_hd__and2b_1
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1010_ clknet_3_2__leaf_clk _0060_ net30 VGND VGND VPWR VPWR uart_rcv.data_buff.packet_data\[7\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_34_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0725_ _0260_ _0301_ _0306_ _0307_ VGND VGND VPWR VPWR _0308_ sky130_fd_sc_hd__a22o_1
X_0656_ _0237_ _0238_ _0239_ _0240_ VGND VGND VPWR VPWR _0241_ sky130_fd_sc_hd__or4_1
X_0587_ net6 uart_tx.clk_cnt\[1\] VGND VGND VPWR VPWR _0186_ sky130_fd_sc_hd__and2b_1
XFILLER_43_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0510_ uart_rcv.tim.clk_cnt\[2\] _0120_ _0119_ VGND VGND VPWR VPWR _0123_ sky130_fd_sc_hd__o21ai_1
Xhold1 uart_rcv.sbd.sync_phase VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0639_ uart_tx.clk_cnt\[11\] uart_tx.clk_cnt\[12\] _0221_ VGND VGND VPWR VPWR _0226_
+ sky130_fd_sc_hd__and3_1
X_0708_ _0249_ _0277_ _0291_ VGND VGND VPWR VPWR _0292_ sky130_fd_sc_hd__a21o_1
XFILLER_0_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0990_ clknet_3_1__leaf_clk _0040_ net28 VGND VGND VPWR VPWR parallel_out2\[3\] sky130_fd_sc_hd__dfstp_2
XFILLER_5_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0973_ clknet_3_2__leaf_clk uart_rcv.tim.bit_count.next_cnt_out\[3\] net32 VGND VGND
+ VPWR VPWR uart_rcv.tim.bit_cnt\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_27_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0956_ clknet_3_3__leaf_clk uart_rcv.tim.clock_count.next_cnt_out\[1\] net32 VGND
+ VGND VPWR VPWR uart_rcv.tim.clk_cnt\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_32_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0887_ _0404_ _0405_ _0406_ VGND VGND VPWR VPWR _0419_ sky130_fd_sc_hd__o21ba_1
XFILLER_11_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput13 bit_period[8] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_2
X_0810_ parallel_out2\[7\] parallel_out2\[3\] _0364_ _0365_ VGND VGND VPWR VPWR _0369_
+ sky130_fd_sc_hd__nand4_1
X_0672_ prod_adder.gen_for_loop\[4\].adder_n.b prod_adder.gen_for_loop\[4\].adder_n.a
+ VGND VGND VPWR VPWR _0256_ sky130_fd_sc_hd__nand2_1
X_0741_ net46 _0316_ _0319_ VGND VGND VPWR VPWR _0000_ sky130_fd_sc_hd__nor3_1
XFILLER_37_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0939_ clknet_3_2__leaf_clk net41 net30 VGND VGND VPWR VPWR uart_rcv.sbd.new_sample
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_7_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0724_ _0249_ net24 _0298_ VGND VGND VPWR VPWR _0307_ sky130_fd_sc_hd__a21o_1
X_0655_ net1 uart_tx.count.next_cnt_out\[0\] VGND VGND VPWR VPWR _0240_ sky130_fd_sc_hd__xor2_1
X_0586_ net10 uart_tx.clk_cnt\[5\] VGND VGND VPWR VPWR _0185_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_35_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Left_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2 uart_rcv.sbd.new_sample VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__dlygate4sd3_1
X_0707_ _0248_ net24 VGND VGND VPWR VPWR _0291_ sky130_fd_sc_hd__and2_1
X_0638_ _0225_ VGND VGND VPWR VPWR uart_tx.count.next_cnt_out\[11\] sky130_fd_sc_hd__inv_2
X_0569_ _0167_ VGND VGND VPWR VPWR _0168_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_35_Left_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_61 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_95 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0972_ clknet_3_2__leaf_clk uart_rcv.tim.bit_count.next_cnt_out\[2\] net32 VGND VGND
+ VPWR VPWR uart_rcv.tim.bit_cnt\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_42_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_38_Left_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_22_Left_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0886_ _0416_ _0417_ VGND VGND VPWR VPWR _0418_ sky130_fd_sc_hd__nor2_1
XFILLER_32_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0955_ clknet_3_3__leaf_clk uart_rcv.tim.clock_count.next_cnt_out\[0\] net31 VGND
+ VGND VPWR VPWR uart_rcv.tim.clk_cnt\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_15_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_94 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput14 bit_period[9] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_2
X_0740_ _0169_ _0317_ _0318_ _0170_ _0167_ VGND VGND VPWR VPWR _0319_ sky130_fd_sc_hd__a32o_1
X_0671_ prod_adder.gen_for_loop\[4\].adder_n.b prod_adder.gen_for_loop\[4\].adder_n.a
+ VGND VGND VPWR VPWR _0255_ sky130_fd_sc_hd__and2_1
XFILLER_20_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0869_ _0383_ _0401_ _0402_ VGND VGND VPWR VPWR _0403_ sky130_fd_sc_hd__and3_1
X_0938_ clknet_3_3__leaf_clk net42 net30 VGND VGND VPWR VPWR uart_rcv.sbd.old_sample
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_7_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0723_ prod_adder.gen_for_loop\[2\].adder_n.b _0305_ VGND VGND VPWR VPWR _0306_ sky130_fd_sc_hd__xor2_1
X_0585_ net12 uart_tx.clk_cnt\[7\] VGND VGND VPWR VPWR _0184_ sky130_fd_sc_hd__nand2b_1
X_0654_ net7 uart_tx.count.next_cnt_out\[2\] VGND VGND VPWR VPWR _0239_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_26_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold3 cntrl.data_ready VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0706_ _0255_ _0257_ _0267_ VGND VGND VPWR VPWR _0290_ sky130_fd_sc_hd__o21ai_1
X_0637_ _0223_ _0224_ VGND VGND VPWR VPWR _0225_ sky130_fd_sc_hd__or2_1
X_0499_ _0110_ _0111_ _0112_ _0113_ VGND VGND VPWR VPWR _0114_ sky130_fd_sc_hd__and4_1
X_0568_ _0081_ _0166_ VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__or2_2
XFILLER_13_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0971_ clknet_3_2__leaf_clk uart_rcv.tim.bit_count.next_cnt_out\[1\] net32 VGND VGND
+ VPWR VPWR uart_rcv.tim.bit_cnt\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_41_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0954_ clknet_3_3__leaf_clk uart_rcv.tim.clock_count.next_roflag net31 VGND VGND
+ VPWR VPWR uart_rcv.shift_strobe sky130_fd_sc_hd__dfrtp_1
X_0885_ parallel_out1\[4\] parallel_out1\[3\] _0415_ VGND VGND VPWR VPWR _0417_ sky130_fd_sc_hd__and3_1
XFILLER_14_110 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0670_ prod_adder.gen_for_loop\[5\].adder_n.b prod_adder.gen_for_loop\[5\].adder_n.a
+ VGND VGND VPWR VPWR _0254_ sky130_fd_sc_hd__or2_1
Xinput15 confirmation VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_1
XFILLER_37_235 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0799_ _0355_ _0358_ VGND VGND VPWR VPWR _0360_ sky130_fd_sc_hd__or2_1
X_0868_ parallel_out1\[4\] parallel_out1\[1\] parallel_out1\[5\] parallel_out1\[0\]
+ VGND VGND VPWR VPWR _0402_ sky130_fd_sc_hd__a22o_1
X_0937_ clknet_3_2__leaf_clk net17 net30 VGND VGND VPWR VPWR uart_rcv.sbd.sync_phase
+ sky130_fd_sc_hd__dfstp_1
XFILLER_43_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_4__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_4__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_0722_ _0262_ _0263_ VGND VGND VPWR VPWR _0305_ sky130_fd_sc_hd__and2b_1
X_0653_ net10 uart_tx.count.next_cnt_out\[5\] VGND VGND VPWR VPWR _0238_ sky130_fd_sc_hd__xor2_1
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0584_ uart_tx.clk_cnt\[3\] net8 VGND VGND VPWR VPWR _0183_ sky130_fd_sc_hd__and2b_1
XFILLER_4_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4 uart_rcv.tim.bit_cnt\[3\] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_22_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_32_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0636_ uart_tx.clk_cnt\[11\] _0221_ _0203_ VGND VGND VPWR VPWR _0224_ sky130_fd_sc_hd__o21ai_1
X_0705_ _0252_ _0269_ _0270_ VGND VGND VPWR VPWR _0289_ sky130_fd_sc_hd__or3_1
X_0498_ _0064_ uart_rcv.tim.clk_cnt\[3\] net14 _0067_ _0095_ VGND VGND VPWR VPWR _0113_
+ sky130_fd_sc_hd__o221a_1
X_0567_ cntrl.state\[1\] cntrl.state\[4\] VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__nand2b_1
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0619_ uart_tx.clk_cnt\[4\] _0208_ uart_tx.clk_cnt\[5\] VGND VGND VPWR VPWR _0213_
+ sky130_fd_sc_hd__a21o_1
XFILLER_5_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0970_ clknet_3_2__leaf_clk net51 net32 VGND VGND VPWR VPWR uart_rcv.tim.bit_cnt\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_35_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0884_ parallel_out1\[4\] parallel_out1\[3\] _0415_ VGND VGND VPWR VPWR _0416_ sky130_fd_sc_hd__a21oi_1
X_0953_ clknet_3_2__leaf_clk _0023_ net30 VGND VGND VPWR VPWR cntrl.framing_error
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput16 n_rst VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__buf_1
XFILLER_37_247 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0936_ clknet_3_2__leaf_clk _0012_ net30 VGND VGND VPWR VPWR rx_data\[7\] sky130_fd_sc_hd__dfstp_1
X_0798_ _0355_ _0358_ VGND VGND VPWR VPWR _0359_ sky130_fd_sc_hd__nand2_1
X_0867_ parallel_out1\[0\] parallel_out1\[4\] parallel_out1\[1\] parallel_out1\[5\]
+ VGND VGND VPWR VPWR _0401_ sky130_fd_sc_hd__nand4_1
XTAP_TAPCELL_ROW_38_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0583_ net14 uart_tx.clk_cnt\[9\] VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__and2b_1
XFILLER_6_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0721_ uart_tx.tx_ctrl.state\[2\] _0251_ _0294_ _0303_ _0300_ VGND VGND VPWR VPWR
+ _0304_ sky130_fd_sc_hd__a41o_1
X_0652_ net13 uart_tx.count.next_cnt_out\[8\] VGND VGND VPWR VPWR _0237_ sky130_fd_sc_hd__xor2_1
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0919_ uart_rcv.data_buff.packet_data\[4\] uart_rcv.data_buff.packet_data\[5\] net25
+ VGND VGND VPWR VPWR _0057_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_26_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold5 prod_adder.gen_for_loop\[7\].adder_n.b VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_3_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0635_ uart_tx.clk_cnt\[11\] _0221_ VGND VGND VPWR VPWR _0223_ sky130_fd_sc_hd__and2_1
X_0566_ uart_rcv.tim.bit_count.next_cnt_out\[1\] uart_rcv.tim.bit_count.next_cnt_out\[2\]
+ uart_rcv.tim.bit_count.next_cnt_out\[3\] uart_rcv.tim.bit_count.next_cnt_out\[0\]
+ VGND VGND VPWR VPWR uart_rcv.tim.bit_count.next_roflag sky130_fd_sc_hd__and4bb_1
X_0704_ _0252_ _0270_ _0269_ VGND VGND VPWR VPWR _0288_ sky130_fd_sc_hd__o21ai_1
X_0497_ _0065_ uart_rcv.tim.clk_cnt\[6\] _0101_ _0102_ _0104_ VGND VGND VPWR VPWR
+ _0112_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0618_ uart_tx.clk_cnt\[4\] uart_tx.clk_cnt\[5\] _0208_ VGND VGND VPWR VPWR _0212_
+ sky130_fd_sc_hd__and3_1
X_0549_ _0064_ uart_rcv.tim.clock_count.next_cnt_out\[3\] VGND VGND VPWR VPWR _0150_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_5_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_142 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0952_ clknet_3_2__leaf_clk uart_rcv.control.next_state\[2\] net30 VGND VGND VPWR
+ VPWR uart_rcv.control.state\[2\] sky130_fd_sc_hd__dfrtp_1
X_0883_ _0411_ _0414_ VGND VGND VPWR VPWR _0415_ sky130_fd_sc_hd__xnor2_1
XFILLER_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput17 serial_in VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_15_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0935_ clknet_3_0__leaf_clk _0011_ net26 VGND VGND VPWR VPWR rx_data\[6\] sky130_fd_sc_hd__dfstp_1
X_0866_ prod_adder.gen_for_loop\[0\].adder_n.a _0384_ _0400_ VGND VGND VPWR VPWR _0045_
+ sky130_fd_sc_hd__a21o_1
X_0797_ _0356_ _0357_ VGND VGND VPWR VPWR _0358_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_38_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0720_ _0260_ _0302_ VGND VGND VPWR VPWR _0303_ sky130_fd_sc_hd__xor2_1
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0651_ _0232_ _0233_ _0234_ _0235_ VGND VGND VPWR VPWR _0236_ sky130_fd_sc_hd__or4_1
X_0582_ net7 uart_tx.clk_cnt\[2\] VGND VGND VPWR VPWR _0181_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_43_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0918_ uart_rcv.data_buff.packet_data\[3\] uart_rcv.data_buff.packet_data\[4\] net25
+ VGND VGND VPWR VPWR _0056_ sky130_fd_sc_hd__mux2_1
X_0849_ parallel_out1\[0\] rx_data\[0\] _0083_ VGND VGND VPWR VPWR _0029_ sky130_fd_sc_hd__mux2_1
XFILLER_17_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold6 uart_tx.tx_ctrl.state\[0\] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0703_ _0250_ _0274_ _0285_ VGND VGND VPWR VPWR _0287_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_29_Left_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0634_ _0221_ _0222_ VGND VGND VPWR VPWR uart_tx.count.next_cnt_out\[10\] sky130_fd_sc_hd__nor2_1
X_0496_ _0069_ uart_rcv.tim.clk_cnt\[11\] _0094_ _0099_ _0103_ VGND VGND VPWR VPWR
+ _0111_ sky130_fd_sc_hd__a2111oi_1
X_0565_ _0163_ _0165_ VGND VGND VPWR VPWR uart_rcv.tim.clock_count.next_roflag sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_13_Left_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0479_ uart_rcv.tim.clk_cnt\[1\] net6 VGND VGND VPWR VPWR _0094_ sky130_fd_sc_hd__and2b_1
X_0617_ net20 _0210_ _0211_ VGND VGND VPWR VPWR uart_tx.count.next_cnt_out\[4\] sky130_fd_sc_hd__and3_1
X_0548_ net10 uart_rcv.tim.clock_count.next_cnt_out\[5\] VGND VGND VPWR VPWR _0149_
+ sky130_fd_sc_hd__xor2_1
XFILLER_39_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_16_Left_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0882_ _0412_ _0413_ VGND VGND VPWR VPWR _0414_ sky130_fd_sc_hd__and2b_1
XFILLER_32_168 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0951_ clknet_3_2__leaf_clk uart_rcv.control.next_state\[1\] net31 VGND VGND VPWR
+ VPWR uart_rcv.control.state\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_1_Left_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0934_ clknet_3_0__leaf_clk _0010_ net26 VGND VGND VPWR VPWR rx_data\[5\] sky130_fd_sc_hd__dfstp_1
X_0865_ parallel_out1\[0\] parallel_out1\[4\] _0383_ VGND VGND VPWR VPWR _0400_ sky130_fd_sc_hd__and3_1
X_0796_ _0344_ _0346_ _0347_ VGND VGND VPWR VPWR _0357_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_43_Left_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_138 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0650_ _0065_ uart_tx.count.next_cnt_out\[6\] VGND VGND VPWR VPWR _0235_ sky130_fd_sc_hd__xnor2_1
X_0581_ net13 uart_tx.clk_cnt\[8\] VGND VGND VPWR VPWR _0180_ sky130_fd_sc_hd__and2b_1
XFILLER_19_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0848_ _0399_ cntrl.state\[4\] _0379_ VGND VGND VPWR VPWR _0028_ sky130_fd_sc_hd__mux2_1
X_0779_ _0339_ _0340_ VGND VGND VPWR VPWR _0341_ sky130_fd_sc_hd__and2b_1
X_0917_ uart_rcv.data_buff.packet_data\[2\] uart_rcv.data_buff.packet_data\[3\] net25
+ VGND VGND VPWR VPWR _0055_ sky130_fd_sc_hd__mux2_1
XFILLER_33_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold7 prod_adder.gen_for_loop\[6\].adder_n.a VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0633_ uart_tx.clk_cnt\[10\] _0219_ net20 VGND VGND VPWR VPWR _0222_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_40_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0702_ _0274_ _0285_ VGND VGND VPWR VPWR _0286_ sky130_fd_sc_hd__nand2_1
X_0564_ _0071_ uart_rcv.tim.clock_count.next_cnt_out\[13\] _0153_ _0164_ VGND VGND
+ VPWR VPWR _0165_ sky130_fd_sc_hd__a211o_1
X_0495_ _0069_ uart_rcv.tim.clk_cnt\[11\] _0093_ _0097_ _0100_ VGND VGND VPWR VPWR
+ _0110_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_200 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Left_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0616_ uart_tx.clk_cnt\[4\] _0208_ VGND VGND VPWR VPWR _0211_ sky130_fd_sc_hd__or2_1
X_0478_ net12 uart_rcv.tim.clk_cnt\[7\] VGND VGND VPWR VPWR _0093_ sky130_fd_sc_hd__nand2b_1
X_0547_ net9 uart_rcv.tim.clock_count.next_cnt_out\[4\] VGND VGND VPWR VPWR _0148_
+ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0881_ parallel_out1\[0\] parallel_out1\[7\] parallel_out1\[6\] parallel_out1\[1\]
+ VGND VGND VPWR VPWR _0413_ sky130_fd_sc_hd__a22o_1
X_0950_ clknet_3_2__leaf_clk uart_rcv.control.next_state\[0\] net31 VGND VGND VPWR
+ VPWR uart_rcv.control.state\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0864_ parallel_out2\[7\] rx_data\[7\] _0087_ VGND VGND VPWR VPWR _0044_ sky130_fd_sc_hd__mux2_1
X_0795_ parallel_out2\[2\] parallel_out2\[5\] _0340_ _0339_ VGND VGND VPWR VPWR _0356_
+ sky130_fd_sc_hd__a31o_1
XFILLER_9_151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0933_ clknet_3_0__leaf_clk _0009_ net26 VGND VGND VPWR VPWR rx_data\[4\] sky130_fd_sc_hd__dfstp_1
XFILLER_3_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_217 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0580_ uart_tx.clk_cnt\[1\] net6 VGND VGND VPWR VPWR _0179_ sky130_fd_sc_hd__nand2b_1
XFILLER_33_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0916_ uart_rcv.data_buff.packet_data\[1\] uart_rcv.data_buff.packet_data\[2\] net25
+ VGND VGND VPWR VPWR _0054_ sky130_fd_sc_hd__mux2_1
X_0778_ parallel_out2\[0\] parallel_out2\[7\] parallel_out2\[6\] parallel_out2\[1\]
+ VGND VGND VPWR VPWR _0340_ sky130_fd_sc_hd__a22o_1
X_0847_ _0398_ _0388_ _0393_ VGND VGND VPWR VPWR _0399_ sky130_fd_sc_hd__or3b_1
XFILLER_3_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold8 cntrl.overrun_error VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__dlygate4sd3_1
X_0563_ _0069_ uart_rcv.tim.clock_count.next_cnt_out\[11\] VGND VGND VPWR VPWR _0164_
+ sky130_fd_sc_hd__xnor2_1
X_0632_ uart_tx.clk_cnt\[9\] uart_tx.clk_cnt\[10\] _0218_ VGND VGND VPWR VPWR _0221_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_40_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0701_ _0248_ _0277_ VGND VGND VPWR VPWR _0285_ sky130_fd_sc_hd__nand2_1
X_0494_ _0098_ _0105_ _0107_ _0108_ VGND VGND VPWR VPWR _0109_ sky130_fd_sc_hd__and4_1
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0615_ uart_tx.clk_cnt\[4\] _0208_ VGND VGND VPWR VPWR _0210_ sky130_fd_sc_hd__nand2_1
X_0546_ _0147_ VGND VGND VPWR VPWR uart_rcv.tim.clock_count.next_cnt_out\[13\] sky130_fd_sc_hd__inv_2
XFILLER_38_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0477_ net7 uart_rcv.tim.clk_cnt\[2\] VGND VGND VPWR VPWR _0092_ sky130_fd_sc_hd__and2b_1
XFILLER_5_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0529_ _0135_ net21 _0134_ VGND VGND VPWR VPWR uart_rcv.tim.clock_count.next_cnt_out\[8\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_25_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0880_ parallel_out1\[0\] parallel_out1\[7\] parallel_out1\[6\] parallel_out1\[1\]
+ VGND VGND VPWR VPWR _0412_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_18_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0932_ clknet_3_0__leaf_clk _0008_ net26 VGND VGND VPWR VPWR rx_data\[3\] sky130_fd_sc_hd__dfstp_1
X_0863_ parallel_out2\[6\] rx_data\[6\] net23 VGND VGND VPWR VPWR _0043_ sky130_fd_sc_hd__mux2_1
X_0794_ _0351_ _0354_ VGND VGND VPWR VPWR _0355_ sky130_fd_sc_hd__xnor2_1
XFILLER_9_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0915_ uart_rcv.data_buff.packet_data\[0\] uart_rcv.data_buff.packet_data\[1\] net25
+ VGND VGND VPWR VPWR _0053_ sky130_fd_sc_hd__mux2_1
X_0777_ parallel_out2\[0\] parallel_out2\[7\] parallel_out2\[6\] parallel_out2\[1\]
+ VGND VGND VPWR VPWR _0339_ sky130_fd_sc_hd__and4_1
X_0846_ cntrl.overrun_error cntrl.framing_error _0374_ VGND VGND VPWR VPWR _0398_
+ sky130_fd_sc_hd__o21ba_1
XFILLER_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold9 prod_adder.gen_for_loop\[6\].adder_n.b VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_3_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0700_ _0275_ _0276_ _0280_ _0283_ VGND VGND VPWR VPWR _0284_ sky130_fd_sc_hd__a211o_1
X_0631_ _0219_ _0220_ VGND VGND VPWR VPWR uart_tx.count.next_cnt_out\[9\] sky130_fd_sc_hd__nor2_1
X_0562_ _0158_ _0159_ _0160_ _0162_ VGND VGND VPWR VPWR _0163_ sky130_fd_sc_hd__or4_1
X_0493_ net13 _0066_ _0070_ uart_rcv.tim.clk_cnt\[12\] _0092_ VGND VGND VPWR VPWR
+ _0108_ sky130_fd_sc_hd__a221oi_1
X_0829_ _0084_ _0381_ VGND VGND VPWR VPWR _0385_ sky130_fd_sc_hd__nand2_1
XFILLER_28_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0476_ net52 _0073_ _0091_ VGND VGND VPWR VPWR uart_rcv.tim.bit_count.next_cnt_out\[2\]
+ sky130_fd_sc_hd__o21a_1
X_0545_ _0145_ _0146_ net21 VGND VGND VPWR VPWR _0147_ sky130_fd_sc_hd__or3b_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0614_ _0208_ _0209_ net20 VGND VGND VPWR VPWR uart_tx.count.next_cnt_out\[3\] sky130_fd_sc_hd__and3b_1
XFILLER_14_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0459_ uart_rcv.control.packet_done _0077_ VGND VGND VPWR VPWR _0078_ sky130_fd_sc_hd__nor2_1
X_0528_ _0066_ _0133_ VGND VGND VPWR VPWR _0135_ sky130_fd_sc_hd__nor2_1
XFILLER_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0862_ parallel_out2\[5\] rx_data\[5\] net23 VGND VGND VPWR VPWR _0042_ sky130_fd_sc_hd__mux2_1
X_0931_ clknet_3_1__leaf_clk _0007_ net28 VGND VGND VPWR VPWR rx_data\[2\] sky130_fd_sc_hd__dfstp_1
X_0793_ _0352_ _0353_ VGND VGND VPWR VPWR _0354_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_5_Left_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0845_ net56 _0391_ _0390_ VGND VGND VPWR VPWR _0027_ sky130_fd_sc_hd__a21o_1
X_0914_ _0440_ _0441_ prod_adder.gen_for_loop\[7\].adder_n.a _0383_ VGND VGND VPWR
+ VPWR _0052_ sky130_fd_sc_hd__o2bb2a_1
X_0776_ parallel_out2\[2\] parallel_out2\[5\] VGND VGND VPWR VPWR _0338_ sky130_fd_sc_hd__nand2_1
XFILLER_30_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0630_ uart_tx.clk_cnt\[9\] _0218_ net20 VGND VGND VPWR VPWR _0220_ sky130_fd_sc_hd__o21ai_1
X_0492_ _0065_ uart_rcv.tim.clk_cnt\[6\] _0071_ uart_rcv.tim.clk_cnt\[13\] _0106_
+ VGND VGND VPWR VPWR _0107_ sky130_fd_sc_hd__o221a_1
X_0561_ net5 _0147_ _0154_ _0161_ VGND VGND VPWR VPWR _0162_ sky130_fd_sc_hd__a211o_1
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0759_ _0063_ _0079_ VGND VGND VPWR VPWR _0324_ sky130_fd_sc_hd__or2_1
X_0828_ _0325_ _0372_ VGND VGND VPWR VPWR _0384_ sky130_fd_sc_hd__or2_2
XFILLER_8_218 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Left_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0613_ uart_tx.clk_cnt\[3\] _0207_ VGND VGND VPWR VPWR _0209_ sky130_fd_sc_hd__or2_1
X_0475_ uart_rcv.control.packet_done _0074_ VGND VGND VPWR VPWR _0091_ sky130_fd_sc_hd__nor2_1
X_0544_ uart_rcv.tim.clk_cnt\[12\] uart_rcv.tim.clk_cnt\[13\] _0142_ VGND VGND VPWR
+ VPWR _0146_ sky130_fd_sc_hd__and3_1
XFILLER_38_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_5__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_5__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_30_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_34_Left_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0458_ _0062_ uart_rcv.tim.bit_cnt\[2\] uart_rcv.tim.bit_cnt\[1\] uart_rcv.tim.bit_cnt\[0\]
+ uart_rcv.shift_strobe VGND VGND VPWR VPWR _0077_ sky130_fd_sc_hd__o311a_1
XFILLER_26_103 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0527_ _0066_ _0133_ VGND VGND VPWR VPWR _0134_ sky130_fd_sc_hd__nand2_1
XFILLER_1_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_18_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_37_Left_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0792_ parallel_out2\[2\] parallel_out2\[6\] parallel_out2\[1\] parallel_out2\[7\]
+ VGND VGND VPWR VPWR _0353_ sky130_fd_sc_hd__a22oi_1
X_0861_ parallel_out2\[4\] rx_data\[4\] net23 VGND VGND VPWR VPWR _0041_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_21_Left_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0930_ clknet_3_3__leaf_clk _0006_ net32 VGND VGND VPWR VPWR rx_data\[1\] sky130_fd_sc_hd__dfstp_1
XFILLER_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_29_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_164 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0775_ _0336_ _0337_ prod_adder.gen_for_loop\[2\].adder_n.b net22 VGND VGND VPWR
+ VPWR _0017_ sky130_fd_sc_hd__a2bb2o_1
X_0844_ _0397_ cntrl.state\[2\] _0379_ VGND VGND VPWR VPWR _0026_ sky130_fd_sc_hd__mux2_1
X_0913_ _0439_ _0440_ _0441_ _0384_ net47 VGND VGND VPWR VPWR _0051_ sky130_fd_sc_hd__a32o_1
XFILLER_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0491_ net9 uart_rcv.tim.clk_cnt\[4\] VGND VGND VPWR VPWR _0106_ sky130_fd_sc_hd__xnor2_1
X_0560_ net2 _0141_ VGND VGND VPWR VPWR _0161_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0758_ _0063_ _0079_ VGND VGND VPWR VPWR _0323_ sky130_fd_sc_hd__nor2_1
X_0827_ _0325_ _0372_ VGND VGND VPWR VPWR _0383_ sky130_fd_sc_hd__nor2_2
X_0689_ uart_tx.tx_ctrl.state\[2\] uart_tx.tx_ctrl.state\[3\] VGND VGND VPWR VPWR
+ _0273_ sky130_fd_sc_hd__nor2_1
XFILLER_28_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_226 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0612_ uart_tx.clk_cnt\[0\] uart_tx.clk_cnt\[1\] uart_tx.clk_cnt\[2\] uart_tx.clk_cnt\[3\]
+ VGND VGND VPWR VPWR _0208_ sky130_fd_sc_hd__and4_1
X_0474_ net55 _0077_ _0090_ VGND VGND VPWR VPWR uart_rcv.tim.bit_count.next_cnt_out\[1\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_38_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0543_ uart_rcv.tim.clk_cnt\[12\] _0142_ uart_rcv.tim.clk_cnt\[13\] VGND VGND VPWR
+ VPWR _0145_ sky130_fd_sc_hd__a21oi_1
X_1026_ clknet_3_7__leaf_clk uart_tx.count.next_roflag net37 VGND VGND VPWR VPWR uart_tx.count.roflag_ff
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_4_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0526_ net21 _0132_ _0133_ VGND VGND VPWR VPWR uart_rcv.tim.clock_count.next_cnt_out\[7\]
+ sky130_fd_sc_hd__and3_1
X_0457_ net44 _0074_ _0076_ uart_rcv.control.packet_done VGND VGND VPWR VPWR uart_rcv.tim.bit_count.next_cnt_out\[3\]
+ sky130_fd_sc_hd__a211oi_1
XFILLER_26_115 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1009_ clknet_3_0__leaf_clk _0059_ net27 VGND VGND VPWR VPWR uart_rcv.data_buff.packet_data\[6\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_1_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_18_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0509_ uart_rcv.tim.clk_cnt\[1\] uart_rcv.tim.clk_cnt\[2\] _0117_ VGND VGND VPWR
+ VPWR _0122_ sky130_fd_sc_hd__and3_1
XFILLER_39_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0860_ parallel_out2\[3\] rx_data\[3\] net23 VGND VGND VPWR VPWR _0040_ sky130_fd_sc_hd__mux2_1
X_0791_ parallel_out2\[7\] parallel_out2\[2\] parallel_out2\[6\] parallel_out2\[1\]
+ VGND VGND VPWR VPWR _0352_ sky130_fd_sc_hd__and4_1
X_0989_ clknet_3_1__leaf_clk _0039_ net28 VGND VGND VPWR VPWR parallel_out2\[2\] sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_37_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0912_ _0384_ _0433_ VGND VGND VPWR VPWR _0441_ sky130_fd_sc_hd__nor2_1
XFILLER_33_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0843_ cntrl.state\[2\] _0324_ _0385_ _0396_ VGND VGND VPWR VPWR _0397_ sky130_fd_sc_hd__o211ai_1
X_0774_ _0328_ _0334_ _0335_ net22 VGND VGND VPWR VPWR _0337_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_3_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_235 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0490_ _0068_ uart_rcv.tim.clk_cnt\[10\] _0070_ uart_rcv.tim.clk_cnt\[12\] _0096_
+ VGND VGND VPWR VPWR _0105_ sky130_fd_sc_hd__o221a_1
XFILLER_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0826_ cntrl.state\[0\] _0079_ _0381_ VGND VGND VPWR VPWR _0382_ sky130_fd_sc_hd__or3_1
X_0688_ prod_adder.gen_for_loop\[7\].adder_n.b prod_adder.gen_for_loop\[7\].adder_n.a
+ VGND VGND VPWR VPWR _0272_ sky130_fd_sc_hd__xor2_1
X_0757_ net18 _0322_ VGND VGND VPWR VPWR _0014_ sky130_fd_sc_hd__nor2_1
XFILLER_28_49 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0542_ uart_rcv.tim.clk_cnt\[12\] _0142_ _0144_ VGND VGND VPWR VPWR uart_rcv.tim.clock_count.next_cnt_out\[12\]
+ sky130_fd_sc_hd__a21oi_1
X_0611_ _0207_ net20 _0206_ VGND VGND VPWR VPWR uart_tx.count.next_cnt_out\[2\] sky130_fd_sc_hd__and3b_1
X_0473_ uart_rcv.control.packet_done _0073_ VGND VGND VPWR VPWR _0090_ sky130_fd_sc_hd__nor2_1
XFILLER_38_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1025_ clknet_3_6__leaf_clk uart_tx.count.next_cnt_out\[13\] net38 VGND VGND VPWR
+ VPWR uart_tx.clk_cnt\[13\] sky130_fd_sc_hd__dfrtp_1
X_0809_ parallel_out2\[7\] parallel_out2\[3\] _0364_ _0365_ VGND VGND VPWR VPWR _0368_
+ sky130_fd_sc_hd__a22o_1
XFILLER_29_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_190 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_94 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_138 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0456_ uart_rcv.tim.bit_cnt\[3\] _0075_ _0074_ VGND VGND VPWR VPWR _0076_ sky130_fd_sc_hd__a21oi_1
XFILLER_6_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0525_ uart_rcv.tim.clk_cnt\[7\] _0130_ VGND VGND VPWR VPWR _0133_ sky130_fd_sc_hd__nand2_1
XFILLER_26_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1008_ clknet_3_0__leaf_clk _0058_ net27 VGND VGND VPWR VPWR uart_rcv.data_buff.packet_data\[5\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_1_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0508_ _0120_ _0121_ _0119_ VGND VGND VPWR VPWR uart_rcv.tim.clock_count.next_cnt_out\[1\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_9_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0790_ parallel_out2\[3\] parallel_out2\[5\] VGND VGND VPWR VPWR _0351_ sky130_fd_sc_hd__nand2_1
XFILLER_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0988_ clknet_3_1__leaf_clk _0038_ net28 VGND VGND VPWR VPWR parallel_out2\[1\] sky130_fd_sc_hd__dfstp_2
XFILLER_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_37_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0842_ cntrl.state\[0\] _0079_ _0086_ _0088_ _0380_ VGND VGND VPWR VPWR _0396_ sky130_fd_sc_hd__o311a_1
X_0911_ parallel_out1\[7\] parallel_out1\[3\] _0434_ _0437_ VGND VGND VPWR VPWR _0440_
+ sky130_fd_sc_hd__nand4_1
XFILLER_33_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0773_ _0334_ _0335_ _0328_ VGND VGND VPWR VPWR _0336_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_3_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_247 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0825_ cntrl.state\[3\] cntrl.state\[2\] VGND VGND VPWR VPWR _0381_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_31_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0687_ _0252_ _0269_ _0270_ VGND VGND VPWR VPWR _0271_ sky130_fd_sc_hd__o21ba_1
X_0756_ net43 _0321_ net48 VGND VGND VPWR VPWR _0322_ sky130_fd_sc_hd__a21oi_1
XFILLER_18_50 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0541_ uart_rcv.tim.clk_cnt\[12\] _0142_ net21 VGND VGND VPWR VPWR _0144_ sky130_fd_sc_hd__o21ai_1
X_0472_ net18 VGND VGND VPWR VPWR _0089_ sky130_fd_sc_hd__inv_2
X_0610_ uart_tx.clk_cnt\[0\] uart_tx.clk_cnt\[1\] uart_tx.clk_cnt\[2\] VGND VGND VPWR
+ VPWR _0207_ sky130_fd_sc_hd__and3_1
X_1024_ clknet_3_7__leaf_clk uart_tx.count.next_cnt_out\[12\] net39 VGND VGND VPWR
+ VPWR uart_tx.clk_cnt\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_15_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0808_ _0367_ prod_adder.gen_for_loop\[5\].adder_n.b net22 VGND VGND VPWR VPWR _0020_
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0739_ uart_tx.count.roflag_ff uart_tx.tx_ctrl.state\[0\] VGND VGND VPWR VPWR _0318_
+ sky130_fd_sc_hd__nor2_1
X_0455_ uart_rcv.tim.bit_cnt\[2\] uart_rcv.tim.bit_cnt\[1\] uart_rcv.tim.bit_cnt\[0\]
+ uart_rcv.shift_strobe VGND VGND VPWR VPWR _0075_ sky130_fd_sc_hd__or4bb_1
XFILLER_6_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0524_ uart_rcv.tim.clk_cnt\[7\] _0130_ VGND VGND VPWR VPWR _0132_ sky130_fd_sc_hd__or2_1
X_1007_ clknet_3_0__leaf_clk _0057_ net27 VGND VGND VPWR VPWR uart_rcv.data_buff.packet_data\[4\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0507_ uart_rcv.tim.clk_cnt\[1\] _0117_ VGND VGND VPWR VPWR _0121_ sky130_fd_sc_hd__or2_1
XFILLER_39_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0987_ clknet_3_1__leaf_clk _0037_ net28 VGND VGND VPWR VPWR parallel_out2\[0\] sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_37_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_25_Left_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0772_ _0332_ _0333_ _0331_ VGND VGND VPWR VPWR _0335_ sky130_fd_sc_hd__o21ai_1
X_0841_ _0395_ cntrl.state\[1\] _0379_ VGND VGND VPWR VPWR _0025_ sky130_fd_sc_hd__mux2_1
X_0910_ parallel_out1\[7\] parallel_out1\[3\] _0434_ _0437_ VGND VGND VPWR VPWR _0439_
+ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_3_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_163 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_64 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0824_ cntrl.overrun_error cntrl.framing_error _0086_ _0372_ VGND VGND VPWR VPWR
+ _0380_ sky130_fd_sc_hd__or4_1
X_0755_ net43 _0089_ _0321_ VGND VGND VPWR VPWR _0013_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_31_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0686_ prod_adder.gen_for_loop\[6\].adder_n.b prod_adder.gen_for_loop\[6\].adder_n.a
+ VGND VGND VPWR VPWR _0270_ sky130_fd_sc_hd__and2_1
XFILLER_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_18_62 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0540_ _0142_ _0143_ VGND VGND VPWR VPWR uart_rcv.tim.clock_count.next_cnt_out\[11\]
+ sky130_fd_sc_hd__nor2_1
X_0471_ _0083_ net23 VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__or2_1
X_1023_ clknet_3_7__leaf_clk uart_tx.count.next_cnt_out\[11\] net39 VGND VGND VPWR
+ VPWR uart_tx.clk_cnt\[11\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_28_Left_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Left_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0807_ _0364_ _0366_ VGND VGND VPWR VPWR _0367_ sky130_fd_sc_hd__xnor2_1
X_0738_ uart_tx.tx_ctrl.state\[1\] uart_tx.tx_ctrl.state\[3\] _0316_ VGND VGND VPWR
+ VPWR _0317_ sky130_fd_sc_hd__o21ai_1
XFILLER_30_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0669_ prod_adder.gen_for_loop\[5\].adder_n.b prod_adder.gen_for_loop\[5\].adder_n.a
+ VGND VGND VPWR VPWR _0253_ sky130_fd_sc_hd__and2_1
XFILLER_43_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0454_ uart_rcv.tim.bit_cnt\[2\] _0073_ VGND VGND VPWR VPWR _0074_ sky130_fd_sc_hd__and2_1
X_0523_ _0130_ _0131_ VGND VGND VPWR VPWR uart_rcv.tim.clock_count.next_cnt_out\[6\]
+ sky130_fd_sc_hd__nor2_1
X_1006_ clknet_3_0__leaf_clk _0056_ net27 VGND VGND VPWR VPWR uart_rcv.data_buff.packet_data\[3\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0506_ uart_rcv.tim.clk_cnt\[1\] _0117_ VGND VGND VPWR VPWR _0120_ sky130_fd_sc_hd__and2_1
XFILLER_36_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0986_ clknet_3_1__leaf_clk _0036_ net29 VGND VGND VPWR VPWR parallel_out1\[7\] sky130_fd_sc_hd__dfstp_2
XFILLER_27_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_0_Left_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0771_ _0331_ _0332_ _0333_ VGND VGND VPWR VPWR _0334_ sky130_fd_sc_hd__or3_1
X_0840_ _0085_ _0382_ _0393_ _0394_ VGND VGND VPWR VPWR _0395_ sky130_fd_sc_hd__nand4_1
XTAP_TAPCELL_ROW_3_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_42_Left_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0969_ clknet_3_2__leaf_clk uart_rcv.tim.bit_count.next_roflag net31 VGND VGND VPWR
+ VPWR uart_rcv.control.packet_done sky130_fd_sc_hd__dfrtp_4
XFILLER_2_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0823_ net17 _0377_ _0378_ VGND VGND VPWR VPWR _0379_ sky130_fd_sc_hd__a21bo_1
X_0685_ _0253_ _0268_ _0254_ VGND VGND VPWR VPWR _0269_ sky130_fd_sc_hd__o21ai_1
X_0754_ rx_data\[7\] uart_rcv.data_buff.packet_data\[7\] _0321_ VGND VGND VPWR VPWR
+ _0012_ sky130_fd_sc_hd__mux2_1
XFILLER_18_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_62 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_116 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_0470_ net23 VGND VGND VPWR VPWR _0088_ sky130_fd_sc_hd__inv_2
X_1022_ clknet_3_6__leaf_clk uart_tx.count.next_cnt_out\[10\] net38 VGND VGND VPWR
+ VPWR uart_tx.clk_cnt\[10\] sky130_fd_sc_hd__dfrtp_1
X_0806_ _0362_ _0365_ VGND VGND VPWR VPWR _0366_ sky130_fd_sc_hd__nand2b_1
X_0668_ prod_adder.gen_for_loop\[6\].adder_n.b prod_adder.gen_for_loop\[6\].adder_n.a
+ VGND VGND VPWR VPWR _0252_ sky130_fd_sc_hd__nor2_1
X_0737_ uart_tx.tx_ctrl.state\[4\] _0274_ _0285_ VGND VGND VPWR VPWR _0316_ sky130_fd_sc_hd__and3_1
X_0599_ _0069_ uart_tx.clk_cnt\[11\] _0172_ _0174_ _0182_ VGND VGND VPWR VPWR _0198_
+ sky130_fd_sc_hd__a2111o_1
XFILLER_43_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0522_ uart_rcv.tim.clk_cnt\[6\] _0128_ net21 VGND VGND VPWR VPWR _0131_ sky130_fd_sc_hd__o21ai_1
X_0453_ uart_rcv.tim.bit_cnt\[1\] uart_rcv.tim.bit_cnt\[0\] net25 VGND VGND VPWR VPWR
+ _0073_ sky130_fd_sc_hd__and3_1
XFILLER_20_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_1005_ clknet_3_1__leaf_clk _0055_ net31 VGND VGND VPWR VPWR uart_rcv.data_buff.packet_data\[2\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_34_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0505_ _0109_ _0114_ _0116_ uart_rcv.control.packet_done VGND VGND VPWR VPWR _0119_
+ sky130_fd_sc_hd__a31oi_2
.ends

