magic
tech sky130A
magscale 1 2
timestamp 1752674710
<< viali >>
rect 31500 89065 31534 89099
rect 32035 89065 32069 89099
rect 33524 89065 33558 89099
rect 34720 89065 34754 89099
rect 35255 89065 35289 89099
rect 36652 89065 36686 89099
rect 37940 89065 37974 89099
rect 39228 89065 39262 89099
rect 39763 89065 39797 89099
rect 41252 89065 41286 89099
rect 42448 89065 42482 89099
rect 42983 89065 43017 89099
rect 44380 89065 44414 89099
rect 45668 89065 45702 89099
rect 46801 89065 46835 89099
rect 56553 89065 56587 89099
rect 57749 89065 57783 89099
rect 68208 89065 68242 89099
rect 69588 89065 69622 89099
rect 70031 89065 70065 89099
rect 71428 89065 71462 89099
rect 72716 89065 72750 89099
rect 74004 89065 74038 89099
rect 74740 89065 74774 89099
rect 75936 89065 75970 89099
rect 77316 89065 77350 89099
rect 77759 89065 77793 89099
rect 79156 89065 79190 89099
rect 80444 89065 80478 89099
rect 81732 89065 81766 89099
rect 82468 89065 82502 89099
rect 25641 88929 25675 88963
rect 62257 88929 62291 88963
rect 15889 88895 15923 88929
rect 16533 88895 16567 88929
rect 19109 88895 19143 88929
rect 19753 88895 19787 88929
rect 22329 88895 22363 88929
rect 23617 88895 23651 88929
rect 24214 88895 24248 88929
rect 28769 88895 28803 88929
rect 30179 88895 30213 88929
rect 31297 88895 31331 88929
rect 32204 88895 32238 88929
rect 33323 88895 33357 88929
rect 34517 88895 34551 88929
rect 35424 88895 35458 88929
rect 36497 88895 36531 88929
rect 37737 88895 37771 88929
rect 39025 88895 39059 88929
rect 39932 88895 39966 88929
rect 41049 88895 41083 88929
rect 42245 88895 42279 88929
rect 43152 88895 43186 88929
rect 44225 88895 44259 88929
rect 45465 88895 45499 88929
rect 17933 88861 17967 88895
rect 21225 88861 21259 88895
rect 24537 88861 24571 88895
rect 26857 88861 26891 88895
rect 27501 88861 27535 88895
rect 49929 88890 49963 88924
rect 52597 88895 52631 88929
rect 53929 88895 53963 88929
rect 55817 88895 55851 88929
rect 57105 88895 57139 88929
rect 59081 88895 59115 88929
rect 60325 88895 60359 88929
rect 61658 88895 61692 88929
rect 66121 88895 66155 88929
rect 66811 88895 66845 88929
rect 68053 88895 68087 88929
rect 69433 88895 69467 88929
rect 70237 88895 70271 88929
rect 71273 88895 71307 88929
rect 72561 88895 72595 88929
rect 73801 88895 73835 88929
rect 74585 88895 74619 88929
rect 75733 88895 75767 88929
rect 77113 88895 77147 88929
rect 77965 88895 77999 88929
rect 79001 88895 79035 88929
rect 80289 88895 80323 88929
rect 81529 88895 81563 88929
rect 82313 88895 82347 88929
rect 50757 88861 50791 88895
rect 54549 88861 54583 88895
rect 58577 88861 58611 88895
rect 61981 88861 62015 88895
rect 63565 88861 63599 88895
rect 64853 88861 64887 88895
rect 16044 88793 16078 88827
rect 16697 88793 16731 88827
rect 18051 88793 18085 88827
rect 19264 88793 19298 88827
rect 19917 88793 19951 88827
rect 21087 88793 21121 88827
rect 22484 88793 22518 88827
rect 23772 88793 23806 88827
rect 25825 88793 25859 88827
rect 26975 88793 27009 88827
rect 27619 88793 27653 88827
rect 28924 88793 28958 88827
rect 30011 88793 30045 88827
rect 52761 88793 52795 88827
rect 54141 88793 54175 88827
rect 54851 88793 54885 88827
rect 55981 88793 56015 88827
rect 57260 88793 57294 88827
rect 58439 88793 58473 88827
rect 59293 88793 59327 88827
rect 60480 88793 60514 88827
rect 62441 88793 62475 88827
rect 63683 88793 63717 88827
rect 65155 88793 65189 88827
rect 66276 88793 66310 88827
rect 66995 88793 67029 88827
rect 48733 88419 48767 88453
rect 49653 88385 49687 88419
rect 49469 87331 49503 87365
rect 50481 87297 50515 87331
rect 30585 86685 30619 86719
rect 30774 86685 30808 86719
rect 50021 86714 50055 86748
rect 51033 86685 51067 86719
rect 29965 86617 29999 86651
rect 31713 86617 31747 86651
rect 5469 80803 5503 80837
rect 88637 80769 88671 80803
rect 5263 80633 5297 80667
rect 88385 80633 88419 80667
rect 5469 79715 5503 79749
rect 88637 79715 88671 79749
rect 5263 79545 5297 79579
rect 88431 79545 88465 79579
rect 5469 78627 5503 78661
rect 88637 78627 88671 78661
rect 5263 78457 5297 78491
rect 88431 78457 88465 78491
rect 5263 77641 5297 77675
rect 88569 77573 88603 77607
rect 5469 77539 5503 77573
rect 88201 77505 88235 77539
rect 88339 75941 88373 75975
rect 5469 75839 5503 75873
rect 88545 75839 88579 75873
rect 5263 75737 5297 75771
rect 88569 75397 88603 75431
rect 5469 75363 5503 75397
rect 88339 75261 88373 75295
rect 5263 75193 5297 75227
rect 88569 74309 88603 74343
rect 5469 74275 5503 74309
rect 88339 74173 88373 74207
rect 5263 74105 5297 74139
rect 5469 73187 5503 73221
rect 88633 73187 88667 73221
rect 5263 73017 5297 73051
rect 88431 73017 88465 73051
rect 5469 72099 5503 72133
rect 88615 72081 88649 72115
rect 5263 71997 5297 72031
rect 88431 71997 88465 72031
rect 88247 70501 88281 70535
rect 5469 70399 5503 70433
rect 88477 70365 88511 70399
rect 5263 70297 5297 70331
rect 88569 69957 88603 69991
rect 5469 69923 5503 69957
rect 88339 69821 88373 69855
rect 5263 69753 5297 69787
rect 88477 69277 88511 69311
rect 5469 68835 5503 68869
rect 88633 68835 88667 68869
rect 5263 68665 5297 68699
rect 88431 68665 88465 68699
rect 5469 67747 5503 67781
rect 88633 67747 88667 67781
rect 5263 67577 5297 67611
rect 88431 67577 88465 67611
rect 5469 66659 5503 66693
rect 88615 66641 88649 66675
rect 5263 66489 5297 66523
rect 88431 66489 88465 66523
rect 5376 65061 5410 65095
rect 5171 64959 5205 64993
rect 88245 64959 88279 64993
rect 88457 64857 88491 64891
rect 5171 64483 5205 64517
rect 88337 64483 88371 64517
rect 5376 64313 5410 64347
rect 88549 64313 88583 64347
rect 5171 63395 5205 63429
rect 88337 63395 88371 63429
rect 5376 63225 5410 63259
rect 88549 63225 88583 63259
rect 5376 62341 5410 62375
rect 88549 62341 88583 62375
rect 5217 62307 5251 62341
rect 88385 62307 88419 62341
rect 5217 61219 5251 61253
rect 88385 61219 88419 61253
rect 5376 61049 5410 61083
rect 88549 61049 88583 61083
rect 5171 59519 5205 59553
rect 88245 59519 88279 59553
rect 5376 59485 5410 59519
rect 88457 59417 88491 59451
rect 5171 59043 5205 59077
rect 88337 59043 88371 59077
rect 5376 58873 5410 58907
rect 88549 58873 88583 58907
rect 5171 57955 5205 57989
rect 88337 57955 88371 57989
rect 5376 57785 5410 57819
rect 88549 57785 88583 57819
rect 5171 56867 5205 56901
rect 88385 56867 88419 56901
rect 5376 56833 5410 56867
rect 88549 56833 88583 56867
rect 5171 55779 5205 55813
rect 88385 55779 88419 55813
rect 5376 55609 5410 55643
rect 88549 55609 88583 55643
rect 5217 55133 5251 55167
rect 7585 54725 7619 54759
rect 6965 54521 6999 54555
rect 88245 54079 88279 54113
rect 5217 54045 5251 54079
rect 88457 54045 88491 54079
rect 5376 53705 5410 53739
rect 5171 53603 5205 53637
rect 88337 53603 88371 53637
rect 88549 53433 88583 53467
rect 5377 53161 5411 53195
rect 5171 52991 5205 53025
rect 88477 52957 88511 52991
rect 5171 52515 5205 52549
rect 88337 52515 88371 52549
rect 5377 52345 5411 52379
rect 88549 52345 88583 52379
rect 5171 51427 5205 51461
rect 88385 51427 88419 51461
rect 5376 51325 5410 51359
rect 88549 51325 88583 51359
rect 5217 49693 5251 49727
rect 88477 49693 88511 49727
rect 88477 48605 88511 48639
rect 88337 48163 88371 48197
rect 88201 47993 88235 48027
rect 88549 47993 88583 48027
rect 5237 47109 5271 47143
rect 5539 46905 5573 46939
rect 88569 46905 88603 46939
rect 5217 45817 5251 45851
rect 5217 44729 5251 44763
rect 5217 44389 5251 44423
rect 88523 43233 88557 43267
rect 5469 43199 5503 43233
rect 5263 43097 5297 43131
rect 88293 43097 88327 43131
rect 5217 42553 5251 42587
rect 5469 42111 5503 42145
rect 88545 42111 88579 42145
rect 5263 42009 5297 42043
rect 88339 42009 88373 42043
rect 5263 41737 5297 41771
rect 88431 41737 88465 41771
rect 5469 41635 5503 41669
rect 88637 41635 88671 41669
rect 5469 39935 5503 39969
rect 88109 39901 88143 39935
rect 88477 39901 88511 39935
rect 5263 39833 5297 39867
rect 5263 38949 5297 38983
rect 88339 38949 88373 38983
rect 5469 38847 5503 38881
rect 88545 38847 88579 38881
rect 5469 37759 5503 37793
rect 88247 37725 88281 37759
rect 88477 37725 88511 37759
rect 5263 37657 5297 37691
rect 5469 36671 5503 36705
rect 88247 36637 88281 36671
rect 88477 36637 88511 36671
rect 5263 36569 5297 36603
rect 5469 36195 5503 36229
rect 88615 36177 88649 36211
rect 5263 36093 5297 36127
rect 88431 36093 88465 36127
rect 5469 34495 5503 34529
rect 88541 34489 88575 34523
rect 5263 34393 5297 34427
rect 88339 34393 88373 34427
rect 5217 33849 5251 33883
rect 5263 33509 5297 33543
rect 5469 33407 5503 33441
rect 88247 33373 88281 33407
rect 88477 33373 88511 33407
rect 5469 32319 5503 32353
rect 88247 32285 88281 32319
rect 88477 32285 88511 32319
rect 5263 32217 5297 32251
rect 5469 31231 5503 31265
rect 88541 31225 88575 31259
rect 5263 31129 5297 31163
rect 88339 31129 88373 31163
rect 5469 30755 5503 30789
rect 88615 30737 88649 30771
rect 5263 30585 5297 30619
rect 88431 30585 88465 30619
rect 5469 29055 5503 29089
rect 88541 29049 88575 29083
rect 5263 28953 5297 28987
rect 88339 28953 88373 28987
rect 5217 27967 5251 28001
rect 88245 27967 88279 28001
rect 5376 27865 5410 27899
rect 88457 27865 88491 27899
rect 5171 26879 5205 26913
rect 88245 26879 88279 26913
rect 5376 26777 5410 26811
rect 88457 26777 88491 26811
rect 5171 25791 5205 25825
rect 88245 25791 88279 25825
rect 5376 25689 5410 25723
rect 88457 25689 88491 25723
rect 5171 25315 5205 25349
rect 88385 25315 88419 25349
rect 5376 25145 5410 25179
rect 88549 25145 88583 25179
rect 5171 23615 5205 23649
rect 88245 23615 88279 23649
rect 5376 23513 5410 23547
rect 88457 23513 88491 23547
rect 5217 22527 5251 22561
rect 88245 22527 88279 22561
rect 5376 22425 5410 22459
rect 88457 22425 88491 22459
rect 5171 21439 5205 21473
rect 88245 21439 88279 21473
rect 5376 21337 5410 21371
rect 88457 21337 88491 21371
rect 5171 20351 5205 20385
rect 88245 20351 88279 20385
rect 5376 20249 5410 20283
rect 88457 20249 88491 20283
rect 5171 19875 5205 19909
rect 88385 19875 88419 19909
rect 5376 19705 5410 19739
rect 88549 19705 88583 19739
rect 5376 18209 5410 18243
rect 88457 18209 88491 18243
rect 5217 18175 5251 18209
rect 88293 18175 88327 18209
rect 5217 17087 5251 17121
rect 88245 17087 88279 17121
rect 5376 16985 5410 17019
rect 88457 16985 88491 17019
rect 5171 15999 5205 16033
rect 88245 15999 88279 16033
rect 5377 15897 5411 15931
rect 88457 15897 88491 15931
rect 5171 14911 5205 14945
rect 88245 14911 88279 14945
rect 5377 14809 5411 14843
rect 88457 14809 88491 14843
rect 5171 14435 5205 14469
rect 88385 14435 88419 14469
rect 5376 14265 5410 14299
rect 88549 14265 88583 14299
rect 82313 5697 82347 5731
rect 82497 5629 82531 5663
rect 13497 5289 13531 5323
rect 14693 5289 14727 5323
rect 31299 5289 31333 5323
rect 33323 5289 33357 5323
rect 34519 5289 34553 5323
rect 35368 5289 35402 5323
rect 36647 5289 36681 5323
rect 37739 5289 37773 5323
rect 39027 5289 39061 5323
rect 41051 5289 41085 5323
rect 44409 5289 44443 5323
rect 46433 5289 46467 5323
rect 68007 5289 68041 5323
rect 69387 5289 69421 5323
rect 70144 5289 70178 5323
rect 72515 5289 72549 5323
rect 73803 5289 73837 5323
rect 74744 5289 74778 5323
rect 75735 5289 75769 5323
rect 77115 5289 77149 5323
rect 77872 5289 77906 5323
rect 82497 5289 82531 5323
rect 32127 5221 32161 5255
rect 39855 5221 39889 5255
rect 42247 5221 42281 5255
rect 43167 5221 43201 5255
rect 71411 5221 71445 5255
rect 79231 5221 79265 5255
rect 80243 5221 80277 5255
rect 44225 5153 44259 5187
rect 46249 5153 46283 5187
rect 82313 5153 82347 5187
rect 15290 5119 15324 5153
rect 15841 5119 15875 5153
rect 16748 5119 16782 5153
rect 17865 5119 17899 5153
rect 19109 5119 19143 5153
rect 19968 5119 20002 5153
rect 21041 5119 21075 5153
rect 22283 5119 22317 5153
rect 23569 5119 23603 5153
rect 24476 5119 24510 5153
rect 25593 5119 25627 5153
rect 26789 5119 26823 5153
rect 27696 5119 27730 5153
rect 28769 5119 28803 5153
rect 30009 5119 30043 5153
rect 12713 5085 12747 5119
rect 13909 5085 13943 5119
rect 15613 5085 15647 5119
rect 31467 5113 31501 5147
rect 31989 5119 32023 5153
rect 33507 5093 33541 5127
rect 34703 5093 34737 5127
rect 35209 5119 35243 5153
rect 36497 5119 36531 5153
rect 37907 5113 37941 5147
rect 39195 5113 39229 5147
rect 39717 5119 39751 5153
rect 41235 5093 41269 5127
rect 52597 5119 52631 5153
rect 53929 5119 53963 5153
rect 54781 5119 54815 5153
rect 55817 5119 55851 5153
rect 57105 5119 57139 5153
rect 58345 5119 58379 5153
rect 59129 5119 59163 5153
rect 60325 5119 60359 5153
rect 61657 5119 61691 5153
rect 62509 5119 62543 5153
rect 63545 5119 63579 5153
rect 64833 5119 64867 5153
rect 66073 5119 66107 5153
rect 66857 5119 66891 5153
rect 42477 5085 42511 5119
rect 42957 5085 42991 5119
rect 68191 5093 68225 5127
rect 69571 5093 69605 5127
rect 69985 5119 70019 5153
rect 71273 5119 71307 5153
rect 72683 5113 72717 5147
rect 73971 5113 74005 5147
rect 74539 5119 74573 5153
rect 75919 5093 75953 5127
rect 77299 5093 77333 5127
rect 77713 5119 77747 5153
rect 79021 5085 79055 5119
rect 80473 5085 80507 5119
rect 16044 5017 16078 5051
rect 16579 5017 16613 5051
rect 18068 5017 18102 5051
rect 19264 5017 19298 5051
rect 19799 5017 19833 5051
rect 21196 5017 21230 5051
rect 22484 5017 22518 5051
rect 23772 5017 23806 5051
rect 24307 5017 24341 5051
rect 25796 5017 25830 5051
rect 26992 5017 27026 5051
rect 27527 5017 27561 5051
rect 28924 5017 28958 5051
rect 30212 5017 30246 5051
rect 52752 5017 52786 5051
rect 54132 5017 54166 5051
rect 54575 5017 54609 5051
rect 55972 5017 56006 5051
rect 57260 5017 57294 5051
rect 58548 5017 58582 5051
rect 59284 5017 59318 5051
rect 60480 5017 60514 5051
rect 61860 5017 61894 5051
rect 62303 5017 62337 5051
rect 63700 5017 63734 5051
rect 64988 5017 65022 5051
rect 66276 5017 66310 5051
rect 67012 5017 67046 5051
<< metal1 >>
rect 4876 89242 88964 89264
rect 4876 89190 18722 89242
rect 18774 89190 18786 89242
rect 18838 89190 18850 89242
rect 18902 89190 18914 89242
rect 18966 89190 18978 89242
rect 19030 89190 37722 89242
rect 37774 89190 37786 89242
rect 37838 89190 37850 89242
rect 37902 89190 37914 89242
rect 37966 89190 37978 89242
rect 38030 89190 56722 89242
rect 56774 89190 56786 89242
rect 56838 89190 56850 89242
rect 56902 89190 56914 89242
rect 56966 89190 56978 89242
rect 57030 89190 75722 89242
rect 75774 89190 75786 89242
rect 75838 89190 75850 89242
rect 75902 89190 75914 89242
rect 75966 89190 75978 89242
rect 76030 89190 88964 89242
rect 4876 89168 88964 89190
rect 31238 89056 31244 89108
rect 31296 89096 31302 89108
rect 31488 89099 31546 89105
rect 31488 89096 31500 89099
rect 31296 89068 31500 89096
rect 31296 89056 31302 89068
rect 31488 89065 31500 89068
rect 31534 89065 31546 89099
rect 31488 89059 31546 89065
rect 31882 89056 31888 89108
rect 31940 89096 31946 89108
rect 32023 89099 32081 89105
rect 32023 89096 32035 89099
rect 31940 89068 32035 89096
rect 31940 89056 31946 89068
rect 32023 89065 32035 89068
rect 32069 89065 32081 89099
rect 32023 89059 32081 89065
rect 33170 89056 33176 89108
rect 33228 89096 33234 89108
rect 33512 89099 33570 89105
rect 33512 89096 33524 89099
rect 33228 89068 33524 89096
rect 33228 89056 33234 89068
rect 33512 89065 33524 89068
rect 33558 89065 33570 89099
rect 33512 89059 33570 89065
rect 34458 89056 34464 89108
rect 34516 89096 34522 89108
rect 34708 89099 34766 89105
rect 34708 89096 34720 89099
rect 34516 89068 34720 89096
rect 34516 89056 34522 89068
rect 34708 89065 34720 89068
rect 34754 89065 34766 89099
rect 34708 89059 34766 89065
rect 35102 89056 35108 89108
rect 35160 89096 35166 89108
rect 35243 89099 35301 89105
rect 35243 89096 35255 89099
rect 35160 89068 35255 89096
rect 35160 89056 35166 89068
rect 35243 89065 35255 89068
rect 35289 89065 35301 89099
rect 35243 89059 35301 89065
rect 36390 89056 36396 89108
rect 36448 89096 36454 89108
rect 36640 89099 36698 89105
rect 36640 89096 36652 89099
rect 36448 89068 36652 89096
rect 36448 89056 36454 89068
rect 36640 89065 36652 89068
rect 36686 89065 36698 89099
rect 36640 89059 36698 89065
rect 37586 89056 37592 89108
rect 37644 89096 37650 89108
rect 37928 89099 37986 89105
rect 37928 89096 37940 89099
rect 37644 89068 37940 89096
rect 37644 89056 37650 89068
rect 37928 89065 37940 89068
rect 37974 89065 37986 89099
rect 37928 89059 37986 89065
rect 38966 89056 38972 89108
rect 39024 89096 39030 89108
rect 39216 89099 39274 89105
rect 39216 89096 39228 89099
rect 39024 89068 39228 89096
rect 39024 89056 39030 89068
rect 39216 89065 39228 89068
rect 39262 89065 39274 89099
rect 39216 89059 39274 89065
rect 39610 89056 39616 89108
rect 39668 89096 39674 89108
rect 39751 89099 39809 89105
rect 39751 89096 39763 89099
rect 39668 89068 39763 89096
rect 39668 89056 39674 89068
rect 39751 89065 39763 89068
rect 39797 89065 39809 89099
rect 39751 89059 39809 89065
rect 40898 89056 40904 89108
rect 40956 89096 40962 89108
rect 41240 89099 41298 89105
rect 41240 89096 41252 89099
rect 40956 89068 41252 89096
rect 40956 89056 40962 89068
rect 41240 89065 41252 89068
rect 41286 89065 41298 89099
rect 41240 89059 41298 89065
rect 42186 89056 42192 89108
rect 42244 89096 42250 89108
rect 42436 89099 42494 89105
rect 42436 89096 42448 89099
rect 42244 89068 42448 89096
rect 42244 89056 42250 89068
rect 42436 89065 42448 89068
rect 42482 89065 42494 89099
rect 42436 89059 42494 89065
rect 42830 89056 42836 89108
rect 42888 89096 42894 89108
rect 42971 89099 43029 89105
rect 42971 89096 42983 89099
rect 42888 89068 42983 89096
rect 42888 89056 42894 89068
rect 42971 89065 42983 89068
rect 43017 89065 43029 89099
rect 42971 89059 43029 89065
rect 44118 89056 44124 89108
rect 44176 89096 44182 89108
rect 44368 89099 44426 89105
rect 44368 89096 44380 89099
rect 44176 89068 44380 89096
rect 44176 89056 44182 89068
rect 44368 89065 44380 89068
rect 44414 89065 44426 89099
rect 44368 89059 44426 89065
rect 45406 89056 45412 89108
rect 45464 89096 45470 89108
rect 45656 89099 45714 89105
rect 45656 89096 45668 89099
rect 45464 89068 45668 89096
rect 45464 89056 45470 89068
rect 45656 89065 45668 89068
rect 45702 89065 45714 89099
rect 45656 89059 45714 89065
rect 46694 89056 46700 89108
rect 46752 89096 46758 89108
rect 46789 89099 46847 89105
rect 46789 89096 46801 89099
rect 46752 89068 46801 89096
rect 46752 89056 46758 89068
rect 46789 89065 46801 89068
rect 46835 89065 46847 89099
rect 46789 89059 46847 89065
rect 56354 89056 56360 89108
rect 56412 89096 56418 89108
rect 56541 89099 56599 89105
rect 56541 89096 56553 89099
rect 56412 89068 56553 89096
rect 56412 89056 56418 89068
rect 56541 89065 56553 89068
rect 56587 89065 56599 89099
rect 56541 89059 56599 89065
rect 57642 89056 57648 89108
rect 57700 89096 57706 89108
rect 57737 89099 57795 89105
rect 57737 89096 57749 89099
rect 57700 89068 57749 89096
rect 57700 89056 57706 89068
rect 57737 89065 57749 89068
rect 57783 89065 57795 89099
rect 57737 89059 57795 89065
rect 67946 89056 67952 89108
rect 68004 89096 68010 89108
rect 68196 89099 68254 89105
rect 68196 89096 68208 89099
rect 68004 89068 68208 89096
rect 68004 89056 68010 89068
rect 68196 89065 68208 89068
rect 68242 89065 68254 89099
rect 68196 89059 68254 89065
rect 69234 89056 69240 89108
rect 69292 89096 69298 89108
rect 69576 89099 69634 89105
rect 69576 89096 69588 89099
rect 69292 89068 69588 89096
rect 69292 89056 69298 89068
rect 69576 89065 69588 89068
rect 69622 89065 69634 89099
rect 69576 89059 69634 89065
rect 69878 89056 69884 89108
rect 69936 89096 69942 89108
rect 70019 89099 70077 89105
rect 70019 89096 70031 89099
rect 69936 89068 70031 89096
rect 69936 89056 69942 89068
rect 70019 89065 70031 89068
rect 70065 89065 70077 89099
rect 70019 89059 70077 89065
rect 71166 89056 71172 89108
rect 71224 89096 71230 89108
rect 71416 89099 71474 89105
rect 71416 89096 71428 89099
rect 71224 89068 71428 89096
rect 71224 89056 71230 89068
rect 71416 89065 71428 89068
rect 71462 89065 71474 89099
rect 71416 89059 71474 89065
rect 72454 89056 72460 89108
rect 72512 89096 72518 89108
rect 72704 89099 72762 89105
rect 72704 89096 72716 89099
rect 72512 89068 72716 89096
rect 72512 89056 72518 89068
rect 72704 89065 72716 89068
rect 72750 89065 72762 89099
rect 72704 89059 72762 89065
rect 73742 89056 73748 89108
rect 73800 89096 73806 89108
rect 73992 89099 74050 89105
rect 73992 89096 74004 89099
rect 73800 89068 74004 89096
rect 73800 89056 73806 89068
rect 73992 89065 74004 89068
rect 74038 89065 74050 89099
rect 73992 89059 74050 89065
rect 74386 89056 74392 89108
rect 74444 89096 74450 89108
rect 74728 89099 74786 89105
rect 74728 89096 74740 89099
rect 74444 89068 74740 89096
rect 74444 89056 74450 89068
rect 74728 89065 74740 89068
rect 74774 89065 74786 89099
rect 74728 89059 74786 89065
rect 75582 89056 75588 89108
rect 75640 89096 75646 89108
rect 75924 89099 75982 89105
rect 75924 89096 75936 89099
rect 75640 89068 75936 89096
rect 75640 89056 75646 89068
rect 75924 89065 75936 89068
rect 75970 89065 75982 89099
rect 75924 89059 75982 89065
rect 76962 89056 76968 89108
rect 77020 89096 77026 89108
rect 77304 89099 77362 89105
rect 77304 89096 77316 89099
rect 77020 89068 77316 89096
rect 77020 89056 77026 89068
rect 77304 89065 77316 89068
rect 77350 89065 77362 89099
rect 77304 89059 77362 89065
rect 77606 89056 77612 89108
rect 77664 89096 77670 89108
rect 77747 89099 77805 89105
rect 77747 89096 77759 89099
rect 77664 89068 77759 89096
rect 77664 89056 77670 89068
rect 77747 89065 77759 89068
rect 77793 89065 77805 89099
rect 77747 89059 77805 89065
rect 78894 89056 78900 89108
rect 78952 89096 78958 89108
rect 79144 89099 79202 89105
rect 79144 89096 79156 89099
rect 78952 89068 79156 89096
rect 78952 89056 78958 89068
rect 79144 89065 79156 89068
rect 79190 89065 79202 89099
rect 79144 89059 79202 89065
rect 80182 89056 80188 89108
rect 80240 89096 80246 89108
rect 80432 89099 80490 89105
rect 80432 89096 80444 89099
rect 80240 89068 80444 89096
rect 80240 89056 80246 89068
rect 80432 89065 80444 89068
rect 80478 89065 80490 89099
rect 80432 89059 80490 89065
rect 81470 89056 81476 89108
rect 81528 89096 81534 89108
rect 81720 89099 81778 89105
rect 81720 89096 81732 89099
rect 81528 89068 81732 89096
rect 81528 89056 81534 89068
rect 81720 89065 81732 89068
rect 81766 89065 81778 89099
rect 81720 89059 81778 89065
rect 82114 89056 82120 89108
rect 82172 89096 82178 89108
rect 82456 89099 82514 89105
rect 82456 89096 82468 89099
rect 82172 89068 82468 89096
rect 82172 89056 82178 89068
rect 82456 89065 82468 89068
rect 82502 89065 82514 89099
rect 82456 89059 82514 89065
rect 15782 88886 15788 88938
rect 15840 88926 15846 88938
rect 15877 88929 15935 88935
rect 15877 88926 15889 88929
rect 15840 88898 15889 88926
rect 15840 88886 15846 88898
rect 15877 88895 15889 88898
rect 15923 88895 15935 88929
rect 15877 88889 15935 88895
rect 16426 88886 16432 88938
rect 16484 88926 16490 88938
rect 16521 88929 16579 88935
rect 16521 88926 16533 88929
rect 16484 88898 16533 88926
rect 16484 88886 16490 88898
rect 16521 88895 16533 88898
rect 16567 88895 16579 88929
rect 16521 88889 16579 88895
rect 17714 88852 17720 88904
rect 17772 88892 17778 88904
rect 17921 88895 17979 88901
rect 17921 88892 17933 88895
rect 17772 88864 17933 88892
rect 17772 88852 17778 88864
rect 17921 88861 17933 88864
rect 17967 88861 17979 88895
rect 19094 88886 19100 88938
rect 19152 88886 19158 88938
rect 19646 88886 19652 88938
rect 19704 88926 19710 88938
rect 19741 88929 19799 88935
rect 19741 88926 19753 88929
rect 19704 88898 19753 88926
rect 19704 88886 19710 88898
rect 19741 88895 19753 88898
rect 19787 88895 19799 88929
rect 19741 88889 19799 88895
rect 17921 88855 17979 88861
rect 20934 88852 20940 88904
rect 20992 88892 20998 88904
rect 21213 88895 21271 88901
rect 21213 88892 21225 88895
rect 20992 88864 21225 88892
rect 20992 88852 20998 88864
rect 21213 88861 21225 88864
rect 21259 88861 21271 88895
rect 22222 88886 22228 88938
rect 22280 88926 22286 88938
rect 22317 88929 22375 88935
rect 22317 88926 22329 88929
rect 22280 88898 22329 88926
rect 22280 88886 22286 88898
rect 22317 88895 22329 88898
rect 22363 88895 22375 88929
rect 22317 88889 22375 88895
rect 23510 88886 23516 88938
rect 23568 88926 23574 88938
rect 23605 88929 23663 88935
rect 23605 88926 23617 88929
rect 23568 88898 23617 88926
rect 23568 88886 23574 88898
rect 23605 88895 23617 88898
rect 23651 88895 23663 88929
rect 23605 88889 23663 88895
rect 24154 88886 24160 88938
rect 24212 88935 24218 88938
rect 24212 88929 24260 88935
rect 24212 88895 24214 88929
rect 24248 88895 24260 88929
rect 25442 88920 25448 88972
rect 25500 88960 25506 88972
rect 25629 88963 25687 88969
rect 25629 88960 25641 88963
rect 25500 88932 25641 88960
rect 25500 88920 25506 88932
rect 25629 88929 25641 88932
rect 25675 88929 25687 88963
rect 25629 88923 25687 88929
rect 24212 88889 24260 88895
rect 24212 88886 24218 88889
rect 21213 88855 21271 88861
rect 24338 88852 24344 88904
rect 24396 88892 24402 88904
rect 24525 88895 24583 88901
rect 24525 88892 24537 88895
rect 24396 88864 24537 88892
rect 24396 88852 24402 88864
rect 24525 88861 24537 88864
rect 24571 88861 24583 88895
rect 24525 88855 24583 88861
rect 26730 88852 26736 88904
rect 26788 88892 26794 88904
rect 26845 88895 26903 88901
rect 26845 88892 26857 88895
rect 26788 88864 26857 88892
rect 26788 88852 26794 88864
rect 26845 88861 26857 88864
rect 26891 88861 26903 88895
rect 26845 88855 26903 88861
rect 27374 88852 27380 88904
rect 27432 88892 27438 88904
rect 27489 88895 27547 88901
rect 27489 88892 27501 88895
rect 27432 88864 27501 88892
rect 27432 88852 27438 88864
rect 27489 88861 27501 88864
rect 27535 88861 27547 88895
rect 28662 88886 28668 88938
rect 28720 88926 28726 88938
rect 28757 88929 28815 88935
rect 28757 88926 28769 88929
rect 28720 88898 28769 88926
rect 28720 88886 28726 88898
rect 28757 88895 28769 88898
rect 28803 88895 28815 88929
rect 28757 88889 28815 88895
rect 29950 88886 29956 88938
rect 30008 88926 30014 88938
rect 30167 88929 30225 88935
rect 30167 88926 30179 88929
rect 30008 88898 30179 88926
rect 30008 88886 30014 88898
rect 30167 88895 30179 88898
rect 30213 88895 30225 88929
rect 31285 88929 31343 88935
rect 31285 88926 31297 88929
rect 30980 88904 31297 88926
rect 30167 88889 30225 88895
rect 27489 88855 27547 88861
rect 30962 88852 30968 88904
rect 31020 88898 31297 88904
rect 31020 88852 31026 88898
rect 31285 88895 31297 88898
rect 31331 88895 31343 88929
rect 31285 88889 31343 88895
rect 32066 88886 32072 88938
rect 32124 88926 32130 88938
rect 32192 88929 32250 88935
rect 32192 88926 32204 88929
rect 32124 88898 32204 88926
rect 32124 88886 32130 88898
rect 32192 88895 32204 88898
rect 32238 88895 32250 88929
rect 32192 88889 32250 88895
rect 33170 88886 33176 88938
rect 33228 88926 33234 88938
rect 33311 88929 33369 88935
rect 33311 88926 33323 88929
rect 33228 88898 33323 88926
rect 33228 88886 33234 88898
rect 33311 88895 33323 88898
rect 33357 88895 33369 88929
rect 33311 88889 33369 88895
rect 34274 88886 34280 88938
rect 34332 88926 34338 88938
rect 34505 88929 34563 88935
rect 34505 88926 34517 88929
rect 34332 88898 34517 88926
rect 34332 88886 34338 88898
rect 34505 88895 34517 88898
rect 34551 88895 34563 88929
rect 34505 88889 34563 88895
rect 35378 88886 35384 88938
rect 35436 88935 35442 88938
rect 35436 88929 35470 88935
rect 35458 88895 35470 88929
rect 35436 88889 35470 88895
rect 35436 88886 35442 88889
rect 36482 88886 36488 88938
rect 36540 88886 36546 88938
rect 37586 88886 37592 88938
rect 37644 88926 37650 88938
rect 37725 88929 37783 88935
rect 37725 88926 37737 88929
rect 37644 88898 37737 88926
rect 37644 88886 37650 88898
rect 37725 88895 37737 88898
rect 37771 88895 37783 88929
rect 37725 88889 37783 88895
rect 38782 88886 38788 88938
rect 38840 88926 38846 88938
rect 39013 88929 39071 88935
rect 39013 88926 39025 88929
rect 38840 88898 39025 88926
rect 38840 88886 38846 88898
rect 39013 88895 39025 88898
rect 39059 88895 39071 88929
rect 39013 88889 39071 88895
rect 39794 88886 39800 88938
rect 39852 88926 39858 88938
rect 39920 88929 39978 88935
rect 39920 88926 39932 88929
rect 39852 88898 39932 88926
rect 39852 88886 39858 88898
rect 39920 88895 39932 88898
rect 39966 88895 39978 88929
rect 39920 88889 39978 88895
rect 40898 88886 40904 88938
rect 40956 88926 40962 88938
rect 41037 88929 41095 88935
rect 41037 88926 41049 88929
rect 40956 88898 41049 88926
rect 40956 88886 40962 88898
rect 41037 88895 41049 88898
rect 41083 88895 41095 88929
rect 41037 88889 41095 88895
rect 42002 88886 42008 88938
rect 42060 88926 42066 88938
rect 42233 88929 42291 88935
rect 42233 88926 42245 88929
rect 42060 88898 42245 88926
rect 42060 88886 42066 88898
rect 42233 88895 42245 88898
rect 42279 88895 42291 88929
rect 42233 88889 42291 88895
rect 43106 88886 43112 88938
rect 43164 88935 43170 88938
rect 43164 88929 43198 88935
rect 43186 88895 43198 88929
rect 43164 88889 43198 88895
rect 43164 88886 43170 88889
rect 44210 88886 44216 88938
rect 44268 88886 44274 88938
rect 45314 88886 45320 88938
rect 45372 88926 45378 88938
rect 45453 88929 45511 88935
rect 45453 88926 45465 88929
rect 45372 88898 45465 88926
rect 45372 88886 45378 88898
rect 45453 88895 45465 88898
rect 45499 88895 45511 88929
rect 45453 88889 45511 88895
rect 49914 88881 49920 88933
rect 49972 88881 49978 88933
rect 50006 88852 50012 88904
rect 50064 88892 50070 88904
rect 50745 88895 50803 88901
rect 50745 88892 50757 88895
rect 50064 88864 50757 88892
rect 50064 88852 50070 88864
rect 50745 88861 50757 88864
rect 50791 88861 50803 88895
rect 52490 88886 52496 88938
rect 52548 88926 52554 88938
rect 52585 88929 52643 88935
rect 52585 88926 52597 88929
rect 52548 88898 52597 88926
rect 52548 88886 52554 88898
rect 52585 88895 52597 88898
rect 52631 88895 52643 88929
rect 52585 88889 52643 88895
rect 53778 88886 53784 88938
rect 53836 88926 53842 88938
rect 53917 88929 53975 88935
rect 53917 88926 53929 88929
rect 53836 88898 53929 88926
rect 53836 88886 53842 88898
rect 53917 88895 53929 88898
rect 53963 88895 53975 88929
rect 53917 88889 53975 88895
rect 50745 88855 50803 88861
rect 54422 88852 54428 88904
rect 54480 88892 54486 88904
rect 54537 88895 54595 88901
rect 54537 88892 54549 88895
rect 54480 88864 54549 88892
rect 54480 88852 54486 88864
rect 54537 88861 54549 88864
rect 54583 88861 54595 88895
rect 55710 88886 55716 88938
rect 55768 88926 55774 88938
rect 55805 88929 55863 88935
rect 55805 88926 55817 88929
rect 55768 88898 55817 88926
rect 55768 88886 55774 88898
rect 55805 88895 55817 88898
rect 55851 88895 55863 88929
rect 55805 88889 55863 88895
rect 57090 88886 57096 88938
rect 57148 88886 57154 88938
rect 54537 88855 54595 88861
rect 58286 88852 58292 88904
rect 58344 88892 58350 88904
rect 58565 88895 58623 88901
rect 58565 88892 58577 88895
rect 58344 88864 58577 88892
rect 58344 88852 58350 88864
rect 58565 88861 58577 88864
rect 58611 88861 58623 88895
rect 58930 88886 58936 88938
rect 58988 88926 58994 88938
rect 59069 88929 59127 88935
rect 59069 88926 59081 88929
rect 58988 88898 59081 88926
rect 58988 88886 58994 88898
rect 59069 88895 59081 88898
rect 59115 88895 59127 88929
rect 59069 88889 59127 88895
rect 60218 88886 60224 88938
rect 60276 88926 60282 88938
rect 60313 88929 60371 88935
rect 60313 88926 60325 88929
rect 60276 88898 60325 88926
rect 60276 88886 60282 88898
rect 60313 88895 60325 88898
rect 60359 88895 60371 88929
rect 60313 88889 60371 88895
rect 61506 88886 61512 88938
rect 61564 88926 61570 88938
rect 61646 88929 61704 88935
rect 61646 88926 61658 88929
rect 61564 88898 61658 88926
rect 61564 88886 61570 88898
rect 61646 88895 61658 88898
rect 61692 88895 61704 88929
rect 62150 88920 62156 88972
rect 62208 88960 62214 88972
rect 62245 88963 62303 88969
rect 62245 88960 62257 88963
rect 62208 88932 62257 88960
rect 62208 88920 62214 88932
rect 62245 88929 62257 88932
rect 62291 88929 62303 88963
rect 62245 88923 62303 88929
rect 61646 88889 61704 88895
rect 61969 88895 62027 88901
rect 58565 88855 58623 88861
rect 61969 88861 61981 88895
rect 62015 88861 62027 88895
rect 61969 88855 62027 88861
rect 15506 88784 15512 88836
rect 15564 88824 15570 88836
rect 16702 88833 16708 88836
rect 16032 88827 16090 88833
rect 16032 88824 16044 88827
rect 15564 88796 16044 88824
rect 15564 88784 15570 88796
rect 16032 88793 16044 88796
rect 16078 88793 16090 88827
rect 16032 88787 16090 88793
rect 16685 88827 16708 88833
rect 16685 88793 16697 88827
rect 16685 88787 16708 88793
rect 16702 88784 16708 88787
rect 16760 88784 16766 88836
rect 17806 88784 17812 88836
rect 17864 88824 17870 88836
rect 18039 88827 18097 88833
rect 18039 88824 18051 88827
rect 17864 88796 18051 88824
rect 17864 88784 17870 88796
rect 18039 88793 18051 88796
rect 18085 88793 18097 88827
rect 18039 88787 18097 88793
rect 18634 88784 18640 88836
rect 18692 88824 18698 88836
rect 19922 88833 19928 88836
rect 19252 88827 19310 88833
rect 19252 88824 19264 88827
rect 18692 88796 19264 88824
rect 18692 88784 18698 88796
rect 19252 88793 19264 88796
rect 19298 88793 19310 88827
rect 19252 88787 19310 88793
rect 19905 88827 19928 88833
rect 19905 88793 19917 88827
rect 19905 88787 19928 88793
rect 19922 88784 19928 88787
rect 19980 88784 19986 88836
rect 21026 88784 21032 88836
rect 21084 88833 21090 88836
rect 21084 88827 21133 88833
rect 21084 88793 21087 88827
rect 21121 88793 21133 88827
rect 21084 88787 21133 88793
rect 21084 88784 21090 88787
rect 22130 88784 22136 88836
rect 22188 88824 22194 88836
rect 22472 88827 22530 88833
rect 22472 88824 22484 88827
rect 22188 88796 22484 88824
rect 22188 88784 22194 88796
rect 22472 88793 22484 88796
rect 22518 88793 22530 88827
rect 22472 88787 22530 88793
rect 23234 88784 23240 88836
rect 23292 88824 23298 88836
rect 23760 88827 23818 88833
rect 23760 88824 23772 88827
rect 23292 88796 23772 88824
rect 23292 88784 23298 88796
rect 23760 88793 23772 88796
rect 23806 88793 23818 88827
rect 23760 88787 23818 88793
rect 25442 88784 25448 88836
rect 25500 88824 25506 88836
rect 25813 88827 25871 88833
rect 25813 88824 25825 88827
rect 25500 88796 25825 88824
rect 25500 88784 25506 88796
rect 25813 88793 25825 88796
rect 25859 88793 25871 88827
rect 25813 88787 25871 88793
rect 26546 88784 26552 88836
rect 26604 88824 26610 88836
rect 27650 88833 27656 88836
rect 26963 88827 27021 88833
rect 26963 88824 26975 88827
rect 26604 88796 26975 88824
rect 26604 88784 26610 88796
rect 26963 88793 26975 88796
rect 27009 88793 27021 88827
rect 26963 88787 27021 88793
rect 27607 88827 27656 88833
rect 27607 88793 27619 88827
rect 27653 88793 27656 88827
rect 27607 88787 27656 88793
rect 27650 88784 27656 88787
rect 27708 88784 27714 88836
rect 28754 88784 28760 88836
rect 28812 88824 28818 88836
rect 28912 88827 28970 88833
rect 28912 88824 28924 88827
rect 28812 88796 28924 88824
rect 28812 88784 28818 88796
rect 28912 88793 28924 88796
rect 28958 88793 28970 88827
rect 28912 88787 28970 88793
rect 29858 88784 29864 88836
rect 29916 88824 29922 88836
rect 52766 88833 52772 88836
rect 29999 88827 30057 88833
rect 29999 88824 30011 88827
rect 29916 88796 30011 88824
rect 29916 88784 29922 88796
rect 29999 88793 30011 88796
rect 30045 88793 30057 88827
rect 29999 88787 30057 88793
rect 52749 88827 52772 88833
rect 52749 88793 52761 88827
rect 52749 88787 52772 88793
rect 52766 88784 52772 88787
rect 52824 88784 52830 88836
rect 54146 88833 54152 88836
rect 54129 88827 54152 88833
rect 54129 88793 54141 88827
rect 54129 88787 54152 88793
rect 54146 88784 54152 88787
rect 54204 88784 54210 88836
rect 54790 88784 54796 88836
rect 54848 88833 54854 88836
rect 55986 88833 55992 88836
rect 54848 88827 54897 88833
rect 54848 88793 54851 88827
rect 54885 88793 54897 88827
rect 54848 88787 54897 88793
rect 55969 88827 55992 88833
rect 55969 88793 55981 88827
rect 55969 88787 55992 88793
rect 54848 88784 54854 88787
rect 55986 88784 55992 88787
rect 56044 88784 56050 88836
rect 57090 88784 57096 88836
rect 57148 88824 57154 88836
rect 57248 88827 57306 88833
rect 57248 88824 57260 88827
rect 57148 88796 57260 88824
rect 57148 88784 57154 88796
rect 57248 88793 57260 88796
rect 57294 88793 57306 88827
rect 57248 88787 57306 88793
rect 58378 88784 58384 88836
rect 58436 88833 58442 88836
rect 59298 88833 59304 88836
rect 58436 88827 58485 88833
rect 58436 88793 58439 88827
rect 58473 88793 58485 88827
rect 58436 88787 58485 88793
rect 59281 88827 59304 88833
rect 59281 88793 59293 88827
rect 59281 88787 59304 88793
rect 58436 88784 58442 88787
rect 59298 88784 59304 88787
rect 59356 88784 59362 88836
rect 60310 88784 60316 88836
rect 60368 88824 60374 88836
rect 60468 88827 60526 88833
rect 60468 88824 60480 88827
rect 60368 88796 60480 88824
rect 60368 88784 60374 88796
rect 60468 88793 60480 88796
rect 60514 88793 60526 88827
rect 60468 88787 60526 88793
rect 61414 88784 61420 88836
rect 61472 88824 61478 88836
rect 61984 88824 62012 88855
rect 63438 88852 63444 88904
rect 63496 88892 63502 88904
rect 63553 88895 63611 88901
rect 63553 88892 63565 88895
rect 63496 88864 63565 88892
rect 63496 88852 63502 88864
rect 63553 88861 63565 88864
rect 63599 88861 63611 88895
rect 63553 88855 63611 88861
rect 64726 88852 64732 88904
rect 64784 88892 64790 88904
rect 64841 88895 64899 88901
rect 64841 88892 64853 88895
rect 64784 88864 64853 88892
rect 64784 88852 64790 88864
rect 64841 88861 64853 88864
rect 64887 88861 64899 88895
rect 66014 88886 66020 88938
rect 66072 88926 66078 88938
rect 66109 88929 66167 88935
rect 66109 88926 66121 88929
rect 66072 88898 66121 88926
rect 66072 88886 66078 88898
rect 66109 88895 66121 88898
rect 66155 88895 66167 88929
rect 66109 88889 66167 88895
rect 66658 88886 66664 88938
rect 66716 88926 66722 88938
rect 66799 88929 66857 88935
rect 66799 88926 66811 88929
rect 66716 88898 66811 88926
rect 66716 88886 66722 88898
rect 66799 88895 66811 88898
rect 66845 88895 66857 88929
rect 66799 88889 66857 88895
rect 68038 88886 68044 88938
rect 68096 88886 68102 88938
rect 69418 88886 69424 88938
rect 69476 88886 69482 88938
rect 70246 88935 70252 88938
rect 70225 88929 70252 88935
rect 70225 88895 70237 88929
rect 70225 88889 70252 88895
rect 70246 88886 70252 88889
rect 70304 88886 70310 88938
rect 71261 88929 71319 88935
rect 71261 88895 71273 88929
rect 71307 88926 71319 88929
rect 71350 88926 71356 88938
rect 71307 88898 71356 88926
rect 71307 88895 71319 88898
rect 71261 88889 71319 88895
rect 71350 88886 71356 88898
rect 71408 88886 71414 88938
rect 72454 88886 72460 88938
rect 72512 88926 72518 88938
rect 72549 88929 72607 88935
rect 72549 88926 72561 88929
rect 72512 88898 72561 88926
rect 72512 88886 72518 88898
rect 72549 88895 72561 88898
rect 72595 88895 72607 88929
rect 72549 88889 72607 88895
rect 73558 88886 73564 88938
rect 73616 88926 73622 88938
rect 73789 88929 73847 88935
rect 73789 88926 73801 88929
rect 73616 88898 73801 88926
rect 73616 88886 73622 88898
rect 73789 88895 73801 88898
rect 73835 88895 73847 88929
rect 73789 88889 73847 88895
rect 74573 88929 74631 88935
rect 74573 88895 74585 88929
rect 74619 88926 74631 88929
rect 74662 88926 74668 88938
rect 74619 88898 74668 88926
rect 74619 88895 74631 88898
rect 74573 88889 74631 88895
rect 74662 88886 74668 88898
rect 74720 88886 74726 88938
rect 75490 88886 75496 88938
rect 75548 88926 75554 88938
rect 75721 88929 75779 88935
rect 75721 88926 75733 88929
rect 75548 88898 75733 88926
rect 75548 88886 75554 88898
rect 75721 88895 75733 88898
rect 75767 88895 75779 88929
rect 75721 88889 75779 88895
rect 76870 88886 76876 88938
rect 76928 88926 76934 88938
rect 77974 88935 77980 88938
rect 77101 88929 77159 88935
rect 77101 88926 77113 88929
rect 76928 88898 77113 88926
rect 76928 88886 76934 88898
rect 77101 88895 77113 88898
rect 77147 88895 77159 88929
rect 77101 88889 77159 88895
rect 77953 88929 77980 88935
rect 77953 88895 77965 88929
rect 77953 88889 77980 88895
rect 77974 88886 77980 88889
rect 78032 88886 78038 88938
rect 78989 88929 79047 88935
rect 78989 88895 79001 88929
rect 79035 88926 79047 88929
rect 79078 88926 79084 88938
rect 79035 88898 79084 88926
rect 79035 88895 79047 88898
rect 78989 88889 79047 88895
rect 79078 88886 79084 88898
rect 79136 88886 79142 88938
rect 80274 88886 80280 88938
rect 80332 88886 80338 88938
rect 81286 88886 81292 88938
rect 81344 88926 81350 88938
rect 81517 88929 81575 88935
rect 81517 88926 81529 88929
rect 81344 88898 81529 88926
rect 81344 88886 81350 88898
rect 81517 88895 81529 88898
rect 81563 88895 81575 88929
rect 81517 88889 81575 88895
rect 82301 88929 82359 88935
rect 82301 88895 82313 88929
rect 82347 88926 82359 88929
rect 82390 88926 82396 88938
rect 82347 88898 82396 88926
rect 82347 88895 82359 88898
rect 82301 88889 82359 88895
rect 82390 88886 82396 88898
rect 82448 88886 82454 88938
rect 64841 88855 64899 88861
rect 61472 88796 62012 88824
rect 62429 88827 62487 88833
rect 61472 88784 61478 88796
rect 62429 88793 62441 88827
rect 62475 88824 62487 88827
rect 62518 88824 62524 88836
rect 62475 88796 62524 88824
rect 62475 88793 62487 88796
rect 62429 88787 62487 88793
rect 62518 88784 62524 88796
rect 62576 88784 62582 88836
rect 63714 88833 63720 88836
rect 63671 88827 63720 88833
rect 63671 88793 63683 88827
rect 63717 88793 63720 88827
rect 63671 88787 63720 88793
rect 63714 88784 63720 88787
rect 63772 88784 63778 88836
rect 65094 88784 65100 88836
rect 65152 88833 65158 88836
rect 65152 88827 65201 88833
rect 65152 88793 65155 88827
rect 65189 88793 65201 88827
rect 65152 88787 65201 88793
rect 65152 88784 65158 88787
rect 65830 88784 65836 88836
rect 65888 88824 65894 88836
rect 66264 88827 66322 88833
rect 66264 88824 66276 88827
rect 65888 88796 66276 88824
rect 65888 88784 65894 88796
rect 66264 88793 66276 88796
rect 66310 88793 66322 88827
rect 66264 88787 66322 88793
rect 66934 88784 66940 88836
rect 66992 88833 66998 88836
rect 66992 88827 67041 88833
rect 66992 88793 66995 88827
rect 67029 88793 67041 88827
rect 66992 88787 67041 88793
rect 66992 88784 66998 88787
rect 4876 88698 88964 88720
rect 4876 88646 19382 88698
rect 19434 88646 19446 88698
rect 19498 88646 19510 88698
rect 19562 88646 19574 88698
rect 19626 88646 19638 88698
rect 19690 88646 38382 88698
rect 38434 88646 38446 88698
rect 38498 88646 38510 88698
rect 38562 88646 38574 88698
rect 38626 88646 38638 88698
rect 38690 88646 57382 88698
rect 57434 88646 57446 88698
rect 57498 88646 57510 88698
rect 57562 88646 57574 88698
rect 57626 88646 57638 88698
rect 57690 88646 76382 88698
rect 76434 88646 76446 88698
rect 76498 88646 76510 88698
rect 76562 88646 76574 88698
rect 76626 88646 76638 88698
rect 76690 88646 88964 88698
rect 4876 88624 88964 88646
rect 48626 88410 48632 88462
rect 48684 88450 48690 88462
rect 48721 88453 48779 88459
rect 48721 88450 48733 88453
rect 48684 88422 48733 88450
rect 48684 88410 48690 88422
rect 48721 88419 48733 88422
rect 48767 88419 48779 88453
rect 48721 88413 48779 88419
rect 49638 88376 49644 88428
rect 49696 88376 49702 88428
rect 4876 88154 88964 88176
rect 4876 88102 18722 88154
rect 18774 88102 18786 88154
rect 18838 88102 18850 88154
rect 18902 88102 18914 88154
rect 18966 88102 18978 88154
rect 19030 88102 37722 88154
rect 37774 88102 37786 88154
rect 37838 88102 37850 88154
rect 37902 88102 37914 88154
rect 37966 88102 37978 88154
rect 38030 88102 56722 88154
rect 56774 88102 56786 88154
rect 56838 88102 56850 88154
rect 56902 88102 56914 88154
rect 56966 88102 56978 88154
rect 57030 88102 75722 88154
rect 75774 88102 75786 88154
rect 75838 88102 75850 88154
rect 75902 88102 75914 88154
rect 75966 88102 75978 88154
rect 76030 88102 88964 88154
rect 4876 88080 88964 88102
rect 4876 87610 88964 87632
rect 4876 87558 19382 87610
rect 19434 87558 19446 87610
rect 19498 87558 19510 87610
rect 19562 87558 19574 87610
rect 19626 87558 19638 87610
rect 19690 87558 38382 87610
rect 38434 87558 38446 87610
rect 38498 87558 38510 87610
rect 38562 87558 38574 87610
rect 38626 87558 38638 87610
rect 38690 87558 57382 87610
rect 57434 87558 57446 87610
rect 57498 87558 57510 87610
rect 57562 87558 57574 87610
rect 57626 87558 57638 87610
rect 57690 87558 76382 87610
rect 76434 87558 76446 87610
rect 76498 87558 76510 87610
rect 76562 87558 76574 87610
rect 76626 87558 76638 87610
rect 76690 87558 88964 87610
rect 4876 87536 88964 87558
rect 49270 87322 49276 87374
rect 49328 87362 49334 87374
rect 49457 87365 49515 87371
rect 49457 87362 49469 87365
rect 49328 87334 49469 87362
rect 49328 87322 49334 87334
rect 49457 87331 49469 87334
rect 49503 87362 49515 87365
rect 49638 87362 49644 87374
rect 49503 87334 49644 87362
rect 49503 87331 49515 87334
rect 49457 87325 49515 87331
rect 49638 87322 49644 87334
rect 49696 87322 49702 87374
rect 50469 87331 50527 87337
rect 50469 87297 50481 87331
rect 50515 87328 50527 87331
rect 83678 87328 83684 87340
rect 50515 87300 83684 87328
rect 50515 87297 50527 87300
rect 50469 87291 50527 87297
rect 83678 87288 83684 87300
rect 83736 87288 83742 87340
rect 4876 87066 88964 87088
rect 4876 87014 5954 87066
rect 6006 87014 6018 87066
rect 6070 87014 6082 87066
rect 6134 87014 6146 87066
rect 6198 87014 6210 87066
rect 6262 87014 18722 87066
rect 18774 87014 18786 87066
rect 18838 87014 18850 87066
rect 18902 87014 18914 87066
rect 18966 87014 18978 87066
rect 19030 87014 37722 87066
rect 37774 87014 37786 87066
rect 37838 87014 37850 87066
rect 37902 87014 37914 87066
rect 37966 87014 37978 87066
rect 38030 87014 56722 87066
rect 56774 87014 56786 87066
rect 56838 87014 56850 87066
rect 56902 87014 56914 87066
rect 56966 87014 56978 87066
rect 57030 87014 75722 87066
rect 75774 87014 75786 87066
rect 75838 87014 75850 87066
rect 75902 87014 75914 87066
rect 75966 87014 75978 87066
rect 76030 87014 87098 87066
rect 87150 87014 87162 87066
rect 87214 87014 87226 87066
rect 87278 87014 87290 87066
rect 87342 87014 87354 87066
rect 87406 87014 88964 87066
rect 4876 86992 88964 87014
rect 30612 86756 37494 86784
rect 7594 86676 7600 86728
rect 7652 86716 7658 86728
rect 30612 86725 30640 86756
rect 30573 86719 30640 86725
rect 7652 86688 27834 86716
rect 7652 86676 7658 86688
rect 27806 86648 27834 86688
rect 30573 86685 30585 86719
rect 30619 86688 30640 86719
rect 30762 86719 30820 86725
rect 30619 86685 30631 86688
rect 30573 86679 30631 86685
rect 30762 86685 30774 86719
rect 30808 86716 30820 86719
rect 37466 86716 37494 86756
rect 47982 86716 47988 86728
rect 30808 86685 30824 86716
rect 37466 86688 47988 86716
rect 30762 86679 30824 86685
rect 29953 86651 30011 86657
rect 29953 86648 29965 86651
rect 27806 86620 29965 86648
rect 29953 86617 29965 86620
rect 29999 86648 30011 86651
rect 30796 86648 30824 86679
rect 47982 86676 47988 86688
rect 48040 86676 48046 86728
rect 50006 86705 50012 86757
rect 50064 86705 50070 86757
rect 51021 86719 51079 86725
rect 51021 86685 51033 86719
rect 51067 86716 51079 86719
rect 84046 86716 84052 86728
rect 51067 86688 84052 86716
rect 51067 86685 51079 86688
rect 51021 86679 51079 86685
rect 84046 86676 84052 86688
rect 84104 86676 84110 86728
rect 29999 86620 30824 86648
rect 29999 86617 30011 86620
rect 29953 86611 30011 86617
rect 31698 86608 31704 86660
rect 31756 86608 31762 86660
rect 4876 86522 88964 86544
rect 4876 86470 6690 86522
rect 6742 86470 6754 86522
rect 6806 86470 6818 86522
rect 6870 86470 6882 86522
rect 6934 86470 6946 86522
rect 6998 86470 19382 86522
rect 19434 86470 19446 86522
rect 19498 86470 19510 86522
rect 19562 86470 19574 86522
rect 19626 86470 19638 86522
rect 19690 86470 38382 86522
rect 38434 86470 38446 86522
rect 38498 86470 38510 86522
rect 38562 86470 38574 86522
rect 38626 86470 38638 86522
rect 38690 86470 57382 86522
rect 57434 86470 57446 86522
rect 57498 86470 57510 86522
rect 57562 86470 57574 86522
rect 57626 86470 57638 86522
rect 57690 86470 76382 86522
rect 76434 86470 76446 86522
rect 76498 86470 76510 86522
rect 76562 86470 76574 86522
rect 76626 86470 76638 86522
rect 76690 86470 87834 86522
rect 87886 86470 87898 86522
rect 87950 86470 87962 86522
rect 88014 86470 88026 86522
rect 88078 86470 88090 86522
rect 88142 86470 88964 86522
rect 4876 86448 88964 86470
rect 4876 85978 7912 86000
rect 4876 85926 5954 85978
rect 6006 85926 6018 85978
rect 6070 85926 6082 85978
rect 6134 85926 6146 85978
rect 6198 85926 6210 85978
rect 6262 85926 7912 85978
rect 4876 85904 7912 85926
rect 86020 85978 88964 86000
rect 86020 85926 87098 85978
rect 87150 85926 87162 85978
rect 87214 85926 87226 85978
rect 87278 85926 87290 85978
rect 87342 85926 87354 85978
rect 87406 85926 88964 85978
rect 86020 85904 88964 85926
rect 4876 85434 7912 85456
rect 4876 85382 6690 85434
rect 6742 85382 6754 85434
rect 6806 85382 6818 85434
rect 6870 85382 6882 85434
rect 6934 85382 6946 85434
rect 6998 85382 7912 85434
rect 4876 85360 7912 85382
rect 86020 85434 88964 85456
rect 86020 85382 87834 85434
rect 87886 85382 87898 85434
rect 87950 85382 87962 85434
rect 88014 85382 88026 85434
rect 88078 85382 88090 85434
rect 88142 85382 88964 85434
rect 86020 85360 88964 85382
rect 4876 84890 7912 84912
rect 4876 84838 5954 84890
rect 6006 84838 6018 84890
rect 6070 84838 6082 84890
rect 6134 84838 6146 84890
rect 6198 84838 6210 84890
rect 6262 84838 7912 84890
rect 4876 84816 7912 84838
rect 86020 84890 88964 84912
rect 86020 84838 87098 84890
rect 87150 84838 87162 84890
rect 87214 84838 87226 84890
rect 87278 84838 87290 84890
rect 87342 84838 87354 84890
rect 87406 84838 88964 84890
rect 86020 84816 88964 84838
rect 4876 84346 7912 84368
rect 4876 84294 6690 84346
rect 6742 84294 6754 84346
rect 6806 84294 6818 84346
rect 6870 84294 6882 84346
rect 6934 84294 6946 84346
rect 6998 84294 7912 84346
rect 4876 84272 7912 84294
rect 86020 84346 88964 84368
rect 86020 84294 87834 84346
rect 87886 84294 87898 84346
rect 87950 84294 87962 84346
rect 88014 84294 88026 84346
rect 88078 84294 88090 84346
rect 88142 84294 88964 84346
rect 13666 84228 13672 84280
rect 13724 84268 13730 84280
rect 50006 84268 50012 84280
rect 13724 84240 50012 84268
rect 13724 84228 13730 84240
rect 50006 84228 50012 84240
rect 50064 84228 50070 84280
rect 86020 84272 88964 84294
rect 12562 84160 12568 84212
rect 12620 84200 12626 84212
rect 48902 84200 48908 84212
rect 12620 84172 48908 84200
rect 12620 84160 12626 84172
rect 48902 84160 48908 84172
rect 48960 84160 48966 84212
rect 11274 84092 11280 84144
rect 11332 84132 11338 84144
rect 31698 84132 31704 84144
rect 11332 84104 31704 84132
rect 11332 84092 11338 84104
rect 31698 84092 31704 84104
rect 31756 84132 31762 84144
rect 47798 84132 47804 84144
rect 31756 84104 47804 84132
rect 31756 84092 31762 84104
rect 47798 84092 47804 84104
rect 47856 84092 47862 84144
rect 4876 83802 7912 83824
rect 4876 83750 5954 83802
rect 6006 83750 6018 83802
rect 6070 83750 6082 83802
rect 6134 83750 6146 83802
rect 6198 83750 6210 83802
rect 6262 83750 7912 83802
rect 4876 83728 7912 83750
rect 86020 83802 88964 83824
rect 86020 83750 87098 83802
rect 87150 83750 87162 83802
rect 87214 83750 87226 83802
rect 87278 83750 87290 83802
rect 87342 83750 87354 83802
rect 87406 83750 88964 83802
rect 86020 83728 88964 83750
rect 4876 83258 7912 83280
rect 4876 83206 6690 83258
rect 6742 83206 6754 83258
rect 6806 83206 6818 83258
rect 6870 83206 6882 83258
rect 6934 83206 6946 83258
rect 6998 83206 7912 83258
rect 4876 83184 7912 83206
rect 86020 83258 88964 83280
rect 86020 83206 87834 83258
rect 87886 83206 87898 83258
rect 87950 83206 87962 83258
rect 88014 83206 88026 83258
rect 88078 83206 88090 83258
rect 88142 83206 88964 83258
rect 86020 83184 88964 83206
rect 4876 82714 7912 82736
rect 4876 82662 5954 82714
rect 6006 82662 6018 82714
rect 6070 82662 6082 82714
rect 6134 82662 6146 82714
rect 6198 82662 6210 82714
rect 6262 82662 7912 82714
rect 4876 82640 7912 82662
rect 86020 82714 88964 82736
rect 86020 82662 87098 82714
rect 87150 82662 87162 82714
rect 87214 82662 87226 82714
rect 87278 82662 87290 82714
rect 87342 82662 87354 82714
rect 87406 82662 88964 82714
rect 86020 82640 88964 82662
rect 4876 82170 7912 82192
rect 4876 82118 6690 82170
rect 6742 82118 6754 82170
rect 6806 82118 6818 82170
rect 6870 82118 6882 82170
rect 6934 82118 6946 82170
rect 6998 82118 7912 82170
rect 4876 82096 7912 82118
rect 86020 82170 88964 82192
rect 86020 82118 87834 82170
rect 87886 82118 87898 82170
rect 87950 82118 87962 82170
rect 88014 82118 88026 82170
rect 88078 82118 88090 82170
rect 88142 82118 88964 82170
rect 86020 82096 88964 82118
rect 4876 81626 7912 81648
rect 4876 81574 5954 81626
rect 6006 81574 6018 81626
rect 6070 81574 6082 81626
rect 6134 81574 6146 81626
rect 6198 81574 6210 81626
rect 6262 81574 7912 81626
rect 4876 81552 7912 81574
rect 86020 81626 88964 81648
rect 86020 81574 87098 81626
rect 87150 81574 87162 81626
rect 87214 81574 87226 81626
rect 87278 81574 87290 81626
rect 87342 81574 87354 81626
rect 87406 81574 88964 81626
rect 86020 81552 88964 81574
rect 4876 81082 7912 81104
rect 4876 81030 6690 81082
rect 6742 81030 6754 81082
rect 6806 81030 6818 81082
rect 6870 81030 6882 81082
rect 6934 81030 6946 81082
rect 6998 81030 7912 81082
rect 4876 81008 7912 81030
rect 86020 81082 88964 81104
rect 86020 81030 87834 81082
rect 87886 81030 87898 81082
rect 87950 81030 87962 81082
rect 88014 81030 88026 81082
rect 88078 81030 88090 81082
rect 88142 81030 88964 81082
rect 86020 81008 88964 81030
rect 5457 80837 5515 80843
rect 5457 80803 5469 80837
rect 5503 80803 5515 80837
rect 5457 80800 5515 80803
rect 7134 80800 7140 80812
rect 5457 80797 7140 80800
rect 5472 80772 7140 80797
rect 7134 80760 7140 80772
rect 7192 80760 7198 80812
rect 88646 80809 88652 80812
rect 88625 80803 88652 80809
rect 88625 80769 88637 80803
rect 88625 80763 88652 80769
rect 88646 80760 88652 80763
rect 88704 80760 88710 80812
rect 2902 80624 2908 80676
rect 2960 80664 2966 80676
rect 5251 80667 5309 80673
rect 5251 80664 5263 80667
rect 2960 80636 5263 80664
rect 2960 80624 2966 80636
rect 5251 80633 5263 80636
rect 5297 80633 5309 80667
rect 5251 80627 5309 80633
rect 84322 80624 84328 80676
rect 84380 80664 84386 80676
rect 88373 80667 88431 80673
rect 88373 80664 88385 80667
rect 84380 80636 88385 80664
rect 84380 80624 84386 80636
rect 88373 80633 88385 80636
rect 88419 80633 88431 80667
rect 88373 80627 88431 80633
rect 4876 80538 7912 80560
rect 4876 80486 5954 80538
rect 6006 80486 6018 80538
rect 6070 80486 6082 80538
rect 6134 80486 6146 80538
rect 6198 80486 6210 80538
rect 6262 80486 7912 80538
rect 4876 80464 7912 80486
rect 86020 80538 88964 80560
rect 86020 80486 87098 80538
rect 87150 80486 87162 80538
rect 87214 80486 87226 80538
rect 87278 80486 87290 80538
rect 87342 80486 87354 80538
rect 87406 80486 88964 80538
rect 86020 80464 88964 80486
rect 4876 79994 7912 80016
rect 4876 79942 6690 79994
rect 6742 79942 6754 79994
rect 6806 79942 6818 79994
rect 6870 79942 6882 79994
rect 6934 79942 6946 79994
rect 6998 79942 7912 79994
rect 4876 79920 7912 79942
rect 86020 79994 88964 80016
rect 86020 79942 87834 79994
rect 87886 79942 87898 79994
rect 87950 79942 87962 79994
rect 88014 79942 88026 79994
rect 88078 79942 88090 79994
rect 88142 79942 88964 79994
rect 86020 79920 88964 79942
rect 88646 79755 88652 79758
rect 5457 79749 5515 79755
rect 5457 79715 5469 79749
rect 5503 79715 5515 79749
rect 88625 79749 88652 79755
rect 5457 79712 5515 79715
rect 7134 79712 7140 79724
rect 5457 79709 7140 79712
rect 5472 79684 7140 79709
rect 7134 79672 7140 79684
rect 7192 79672 7198 79724
rect 88625 79715 88637 79749
rect 88625 79709 88652 79715
rect 88646 79706 88652 79709
rect 88704 79706 88710 79758
rect 2718 79536 2724 79588
rect 2776 79576 2782 79588
rect 5251 79579 5309 79585
rect 5251 79576 5263 79579
rect 2776 79548 5263 79576
rect 2776 79536 2782 79548
rect 5251 79545 5263 79548
rect 5297 79545 5309 79579
rect 5251 79539 5309 79545
rect 84322 79536 84328 79588
rect 84380 79576 84386 79588
rect 88419 79579 88477 79585
rect 88419 79576 88431 79579
rect 84380 79548 88431 79576
rect 84380 79536 84386 79548
rect 88419 79545 88431 79548
rect 88465 79545 88477 79579
rect 88419 79539 88477 79545
rect 4876 79450 7912 79472
rect 4876 79398 5954 79450
rect 6006 79398 6018 79450
rect 6070 79398 6082 79450
rect 6134 79398 6146 79450
rect 6198 79398 6210 79450
rect 6262 79398 7912 79450
rect 4876 79376 7912 79398
rect 86020 79450 88964 79472
rect 86020 79398 87098 79450
rect 87150 79398 87162 79450
rect 87214 79398 87226 79450
rect 87278 79398 87290 79450
rect 87342 79398 87354 79450
rect 87406 79398 88964 79450
rect 86020 79376 88964 79398
rect 4876 78906 7912 78928
rect 4876 78854 6690 78906
rect 6742 78854 6754 78906
rect 6806 78854 6818 78906
rect 6870 78854 6882 78906
rect 6934 78854 6946 78906
rect 6998 78854 7912 78906
rect 4876 78832 7912 78854
rect 86020 78906 88964 78928
rect 86020 78854 87834 78906
rect 87886 78854 87898 78906
rect 87950 78854 87962 78906
rect 88014 78854 88026 78906
rect 88078 78854 88090 78906
rect 88142 78854 88964 78906
rect 86020 78832 88964 78854
rect 88646 78667 88652 78670
rect 5457 78661 5515 78667
rect 5457 78627 5469 78661
rect 5503 78627 5515 78661
rect 88625 78661 88652 78667
rect 5457 78624 5515 78627
rect 7134 78624 7140 78636
rect 5457 78621 7140 78624
rect 5472 78596 7140 78621
rect 7134 78584 7140 78596
rect 7192 78584 7198 78636
rect 88625 78627 88637 78661
rect 88625 78621 88652 78627
rect 88646 78618 88652 78621
rect 88704 78618 88710 78670
rect 2902 78448 2908 78500
rect 2960 78488 2966 78500
rect 5251 78491 5309 78497
rect 5251 78488 5263 78491
rect 2960 78460 5263 78488
rect 2960 78448 2966 78460
rect 5251 78457 5263 78460
rect 5297 78457 5309 78491
rect 5251 78451 5309 78457
rect 84322 78448 84328 78500
rect 84380 78488 84386 78500
rect 88419 78491 88477 78497
rect 88419 78488 88431 78491
rect 84380 78460 88431 78488
rect 84380 78448 84386 78460
rect 88419 78457 88431 78460
rect 88465 78457 88477 78491
rect 88419 78451 88477 78457
rect 4876 78362 7912 78384
rect 4876 78310 5954 78362
rect 6006 78310 6018 78362
rect 6070 78310 6082 78362
rect 6134 78310 6146 78362
rect 6198 78310 6210 78362
rect 6262 78310 7912 78362
rect 4876 78288 7912 78310
rect 86020 78362 88964 78384
rect 86020 78310 87098 78362
rect 87150 78310 87162 78362
rect 87214 78310 87226 78362
rect 87278 78310 87290 78362
rect 87342 78310 87354 78362
rect 87406 78310 88964 78362
rect 86020 78288 88964 78310
rect 4876 77818 7912 77840
rect 4876 77766 6690 77818
rect 6742 77766 6754 77818
rect 6806 77766 6818 77818
rect 6870 77766 6882 77818
rect 6934 77766 6946 77818
rect 6998 77766 7912 77818
rect 4876 77744 7912 77766
rect 86020 77818 88964 77840
rect 86020 77766 87834 77818
rect 87886 77766 87898 77818
rect 87950 77766 87962 77818
rect 88014 77766 88026 77818
rect 88078 77766 88090 77818
rect 88142 77766 88964 77818
rect 86020 77744 88964 77766
rect 4374 77632 4380 77684
rect 4432 77672 4438 77684
rect 5251 77675 5309 77681
rect 5251 77672 5263 77675
rect 4432 77644 5263 77672
rect 4432 77632 4438 77644
rect 5251 77641 5263 77644
rect 5297 77641 5309 77675
rect 5251 77635 5309 77641
rect 88557 77607 88615 77613
rect 5457 77573 5515 77579
rect 5457 77539 5469 77573
rect 5503 77570 5515 77573
rect 5662 77570 5668 77582
rect 5503 77542 5668 77570
rect 5503 77539 5515 77542
rect 5457 77533 5515 77539
rect 5662 77530 5668 77542
rect 5720 77530 5726 77582
rect 88557 77573 88569 77607
rect 88603 77604 88615 77607
rect 90026 77604 90032 77616
rect 88603 77576 90032 77604
rect 88603 77573 88615 77576
rect 88557 77567 88615 77573
rect 90026 77564 90032 77576
rect 90084 77564 90090 77616
rect 88189 77539 88247 77545
rect 88189 77505 88201 77539
rect 88235 77505 88247 77539
rect 88189 77499 88247 77505
rect 84322 77428 84328 77480
rect 84380 77468 84386 77480
rect 88204 77468 88232 77499
rect 84380 77440 88232 77468
rect 84380 77428 84386 77440
rect 4876 77274 7912 77296
rect 4876 77222 5954 77274
rect 6006 77222 6018 77274
rect 6070 77222 6082 77274
rect 6134 77222 6146 77274
rect 6198 77222 6210 77274
rect 6262 77222 7912 77274
rect 4876 77200 7912 77222
rect 86020 77274 88964 77296
rect 86020 77222 87098 77274
rect 87150 77222 87162 77274
rect 87214 77222 87226 77274
rect 87278 77222 87290 77274
rect 87342 77222 87354 77274
rect 87406 77222 88964 77274
rect 86020 77200 88964 77222
rect 4876 76730 7912 76752
rect 4876 76678 6690 76730
rect 6742 76678 6754 76730
rect 6806 76678 6818 76730
rect 6870 76678 6882 76730
rect 6934 76678 6946 76730
rect 6998 76678 7912 76730
rect 4876 76656 7912 76678
rect 86020 76730 88964 76752
rect 86020 76678 87834 76730
rect 87886 76678 87898 76730
rect 87950 76678 87962 76730
rect 88014 76678 88026 76730
rect 88078 76678 88090 76730
rect 88142 76678 88964 76730
rect 86020 76656 88964 76678
rect 4876 76186 7912 76208
rect 4876 76134 5954 76186
rect 6006 76134 6018 76186
rect 6070 76134 6082 76186
rect 6134 76134 6146 76186
rect 6198 76134 6210 76186
rect 6262 76134 7912 76186
rect 4876 76112 7912 76134
rect 86020 76186 88964 76208
rect 86020 76134 87098 76186
rect 87150 76134 87162 76186
rect 87214 76134 87226 76186
rect 87278 76134 87290 76186
rect 87342 76134 87354 76186
rect 87406 76134 88964 76186
rect 86020 76112 88964 76134
rect 84322 75932 84328 75984
rect 84380 75972 84386 75984
rect 88327 75975 88385 75981
rect 88327 75972 88339 75975
rect 84380 75944 88339 75972
rect 84380 75932 84386 75944
rect 88327 75941 88339 75944
rect 88373 75941 88385 75975
rect 88327 75935 88385 75941
rect 7134 75904 7140 75916
rect 5457 75873 5515 75879
rect 5457 75839 5469 75873
rect 5503 75870 5515 75873
rect 5772 75876 7140 75904
rect 5772 75870 5800 75876
rect 5503 75842 5800 75870
rect 7134 75864 7140 75876
rect 7192 75864 7198 75916
rect 88533 75873 88591 75879
rect 5503 75839 5515 75842
rect 5457 75833 5515 75839
rect 88533 75839 88545 75873
rect 88579 75870 88591 75873
rect 88579 75848 88784 75870
rect 88579 75842 88744 75848
rect 88579 75839 88591 75842
rect 88533 75833 88591 75839
rect 88738 75796 88744 75842
rect 88796 75796 88802 75848
rect 2902 75728 2908 75780
rect 2960 75768 2966 75780
rect 5251 75771 5309 75777
rect 5251 75768 5263 75771
rect 2960 75740 5263 75768
rect 2960 75728 2966 75740
rect 5251 75737 5263 75740
rect 5297 75737 5309 75771
rect 5251 75731 5309 75737
rect 4876 75642 7912 75664
rect 4876 75590 6690 75642
rect 6742 75590 6754 75642
rect 6806 75590 6818 75642
rect 6870 75590 6882 75642
rect 6934 75590 6946 75642
rect 6998 75590 7912 75642
rect 4876 75568 7912 75590
rect 86020 75642 88964 75664
rect 86020 75590 87834 75642
rect 87886 75590 87898 75642
rect 87950 75590 87962 75642
rect 88014 75590 88026 75642
rect 88078 75590 88090 75642
rect 88142 75590 88964 75642
rect 86020 75568 88964 75590
rect 5457 75397 5515 75403
rect 5457 75363 5469 75397
rect 5503 75394 5515 75397
rect 5503 75366 5800 75394
rect 88554 75388 88560 75440
rect 88612 75388 88618 75440
rect 5503 75363 5515 75366
rect 5457 75357 5515 75363
rect 5772 75360 5800 75366
rect 7134 75360 7140 75372
rect 5772 75332 7140 75360
rect 7134 75320 7140 75332
rect 7192 75320 7198 75372
rect 84322 75252 84328 75304
rect 84380 75292 84386 75304
rect 88327 75295 88385 75301
rect 88327 75292 88339 75295
rect 84380 75264 88339 75292
rect 84380 75252 84386 75264
rect 88327 75261 88339 75264
rect 88373 75261 88385 75295
rect 88327 75255 88385 75261
rect 2902 75184 2908 75236
rect 2960 75224 2966 75236
rect 5251 75227 5309 75233
rect 5251 75224 5263 75227
rect 2960 75196 5263 75224
rect 2960 75184 2966 75196
rect 5251 75193 5263 75196
rect 5297 75193 5309 75227
rect 5251 75187 5309 75193
rect 4876 75098 7912 75120
rect 4876 75046 5954 75098
rect 6006 75046 6018 75098
rect 6070 75046 6082 75098
rect 6134 75046 6146 75098
rect 6198 75046 6210 75098
rect 6262 75046 7912 75098
rect 4876 75024 7912 75046
rect 86020 75098 88964 75120
rect 86020 75046 87098 75098
rect 87150 75046 87162 75098
rect 87214 75046 87226 75098
rect 87278 75046 87290 75098
rect 87342 75046 87354 75098
rect 87406 75046 88964 75098
rect 86020 75024 88964 75046
rect 4876 74554 7912 74576
rect 4876 74502 6690 74554
rect 6742 74502 6754 74554
rect 6806 74502 6818 74554
rect 6870 74502 6882 74554
rect 6934 74502 6946 74554
rect 6998 74502 7912 74554
rect 4876 74480 7912 74502
rect 86020 74554 88964 74576
rect 86020 74502 87834 74554
rect 87886 74502 87898 74554
rect 87950 74502 87962 74554
rect 88014 74502 88026 74554
rect 88078 74502 88090 74554
rect 88142 74502 88964 74554
rect 86020 74480 88964 74502
rect 5457 74309 5515 74315
rect 5457 74275 5469 74309
rect 5503 74306 5515 74309
rect 5503 74278 5800 74306
rect 88554 74300 88560 74352
rect 88612 74300 88618 74352
rect 5503 74275 5515 74278
rect 5457 74269 5515 74275
rect 5772 74272 5800 74278
rect 7134 74272 7140 74284
rect 5772 74244 7140 74272
rect 7134 74232 7140 74244
rect 7192 74232 7198 74284
rect 84322 74164 84328 74216
rect 84380 74204 84386 74216
rect 88327 74207 88385 74213
rect 88327 74204 88339 74207
rect 84380 74176 88339 74204
rect 84380 74164 84386 74176
rect 88327 74173 88339 74176
rect 88373 74173 88385 74207
rect 88327 74167 88385 74173
rect 2902 74096 2908 74148
rect 2960 74136 2966 74148
rect 5251 74139 5309 74145
rect 5251 74136 5263 74139
rect 2960 74108 5263 74136
rect 2960 74096 2966 74108
rect 5251 74105 5263 74108
rect 5297 74105 5309 74139
rect 5251 74099 5309 74105
rect 4876 74010 7912 74032
rect 4876 73958 5954 74010
rect 6006 73958 6018 74010
rect 6070 73958 6082 74010
rect 6134 73958 6146 74010
rect 6198 73958 6210 74010
rect 6262 73958 7912 74010
rect 4876 73936 7912 73958
rect 86020 74010 88964 74032
rect 86020 73958 87098 74010
rect 87150 73958 87162 74010
rect 87214 73958 87226 74010
rect 87278 73958 87290 74010
rect 87342 73958 87354 74010
rect 87406 73958 88964 74010
rect 86020 73936 88964 73958
rect 4876 73466 7912 73488
rect 4876 73414 6690 73466
rect 6742 73414 6754 73466
rect 6806 73414 6818 73466
rect 6870 73414 6882 73466
rect 6934 73414 6946 73466
rect 6998 73414 7912 73466
rect 4876 73392 7912 73414
rect 86020 73466 88964 73488
rect 86020 73414 87834 73466
rect 87886 73414 87898 73466
rect 87950 73414 87962 73466
rect 88014 73414 88026 73466
rect 88078 73414 88090 73466
rect 88142 73414 88964 73466
rect 86020 73392 88964 73414
rect 88646 73227 88652 73230
rect 5457 73221 5515 73227
rect 5457 73187 5469 73221
rect 5503 73218 5515 73221
rect 88621 73221 88652 73227
rect 5503 73190 5800 73218
rect 5503 73187 5515 73190
rect 5457 73181 5515 73187
rect 5772 73184 5800 73190
rect 7134 73184 7140 73196
rect 5772 73156 7140 73184
rect 7134 73144 7140 73156
rect 7192 73144 7198 73196
rect 88621 73187 88633 73221
rect 88621 73181 88652 73187
rect 88646 73178 88652 73181
rect 88704 73178 88710 73230
rect 2902 73008 2908 73060
rect 2960 73048 2966 73060
rect 5251 73051 5309 73057
rect 5251 73048 5263 73051
rect 2960 73020 5263 73048
rect 2960 73008 2966 73020
rect 5251 73017 5263 73020
rect 5297 73017 5309 73051
rect 5251 73011 5309 73017
rect 84322 73008 84328 73060
rect 84380 73048 84386 73060
rect 88419 73051 88477 73057
rect 88419 73048 88431 73051
rect 84380 73020 88431 73048
rect 84380 73008 84386 73020
rect 88419 73017 88431 73020
rect 88465 73017 88477 73051
rect 88419 73011 88477 73017
rect 4876 72922 7912 72944
rect 4876 72870 5954 72922
rect 6006 72870 6018 72922
rect 6070 72870 6082 72922
rect 6134 72870 6146 72922
rect 6198 72870 6210 72922
rect 6262 72870 7912 72922
rect 4876 72848 7912 72870
rect 86020 72922 88964 72944
rect 86020 72870 87098 72922
rect 87150 72870 87162 72922
rect 87214 72870 87226 72922
rect 87278 72870 87290 72922
rect 87342 72870 87354 72922
rect 87406 72870 88964 72922
rect 86020 72848 88964 72870
rect 4876 72378 7912 72400
rect 4876 72326 6690 72378
rect 6742 72326 6754 72378
rect 6806 72326 6818 72378
rect 6870 72326 6882 72378
rect 6934 72326 6946 72378
rect 6998 72326 7912 72378
rect 4876 72304 7912 72326
rect 86020 72378 88964 72400
rect 86020 72326 87834 72378
rect 87886 72326 87898 72378
rect 87950 72326 87962 72378
rect 88014 72326 88026 72378
rect 88078 72326 88090 72378
rect 88142 72326 88964 72378
rect 86020 72304 88964 72326
rect 5457 72133 5515 72139
rect 5457 72099 5469 72133
rect 5503 72130 5515 72133
rect 5662 72130 5668 72142
rect 5503 72102 5668 72130
rect 5503 72099 5515 72102
rect 5457 72093 5515 72099
rect 5662 72090 5668 72102
rect 5720 72090 5726 72142
rect 88603 72115 88661 72121
rect 88603 72081 88615 72115
rect 88649 72112 88661 72115
rect 88649 72096 88876 72112
rect 90118 72096 90124 72108
rect 88649 72084 90124 72096
rect 88649 72081 88661 72084
rect 88603 72075 88661 72081
rect 88848 72068 90124 72084
rect 90118 72056 90124 72068
rect 90176 72056 90182 72108
rect 4374 71988 4380 72040
rect 4432 72028 4438 72040
rect 5251 72031 5309 72037
rect 5251 72028 5263 72031
rect 4432 72000 5263 72028
rect 4432 71988 4438 72000
rect 5251 71997 5263 72000
rect 5297 71997 5309 72031
rect 5251 71991 5309 71997
rect 87174 71988 87180 72040
rect 87232 72028 87238 72040
rect 88419 72031 88477 72037
rect 88419 72028 88431 72031
rect 87232 72000 88431 72028
rect 87232 71988 87238 72000
rect 88419 71997 88431 72000
rect 88465 71997 88477 72031
rect 88419 71991 88477 71997
rect 4876 71834 7912 71856
rect 4876 71782 5954 71834
rect 6006 71782 6018 71834
rect 6070 71782 6082 71834
rect 6134 71782 6146 71834
rect 6198 71782 6210 71834
rect 6262 71782 7912 71834
rect 4876 71760 7912 71782
rect 86020 71834 88964 71856
rect 86020 71782 87098 71834
rect 87150 71782 87162 71834
rect 87214 71782 87226 71834
rect 87278 71782 87290 71834
rect 87342 71782 87354 71834
rect 87406 71782 88964 71834
rect 86020 71760 88964 71782
rect 4876 71290 7912 71312
rect 4876 71238 6690 71290
rect 6742 71238 6754 71290
rect 6806 71238 6818 71290
rect 6870 71238 6882 71290
rect 6934 71238 6946 71290
rect 6998 71238 7912 71290
rect 4876 71216 7912 71238
rect 86020 71290 88964 71312
rect 86020 71238 87834 71290
rect 87886 71238 87898 71290
rect 87950 71238 87962 71290
rect 88014 71238 88026 71290
rect 88078 71238 88090 71290
rect 88142 71238 88964 71290
rect 86020 71216 88964 71238
rect 4876 70746 7912 70768
rect 4876 70694 5954 70746
rect 6006 70694 6018 70746
rect 6070 70694 6082 70746
rect 6134 70694 6146 70746
rect 6198 70694 6210 70746
rect 6262 70694 7912 70746
rect 4876 70672 7912 70694
rect 86020 70746 88964 70768
rect 86020 70694 87098 70746
rect 87150 70694 87162 70746
rect 87214 70694 87226 70746
rect 87278 70694 87290 70746
rect 87342 70694 87354 70746
rect 87406 70694 88964 70746
rect 86020 70672 88964 70694
rect 84322 70492 84328 70544
rect 84380 70532 84386 70544
rect 88235 70535 88293 70541
rect 88235 70532 88247 70535
rect 84380 70504 88247 70532
rect 84380 70492 84386 70504
rect 88235 70501 88247 70504
rect 88281 70501 88293 70535
rect 88235 70495 88293 70501
rect 5457 70433 5515 70439
rect 5457 70399 5469 70433
rect 5503 70430 5515 70433
rect 5662 70430 5668 70442
rect 5503 70402 5668 70430
rect 5503 70399 5515 70402
rect 5457 70393 5515 70399
rect 5662 70390 5668 70402
rect 5720 70390 5726 70442
rect 88465 70399 88523 70405
rect 88465 70365 88477 70399
rect 88511 70396 88523 70399
rect 89934 70396 89940 70408
rect 88511 70368 89940 70396
rect 88511 70365 88523 70368
rect 88465 70359 88523 70365
rect 89934 70356 89940 70368
rect 89992 70356 89998 70408
rect 2902 70288 2908 70340
rect 2960 70328 2966 70340
rect 5251 70331 5309 70337
rect 5251 70328 5263 70331
rect 2960 70300 5263 70328
rect 2960 70288 2966 70300
rect 5251 70297 5263 70300
rect 5297 70297 5309 70331
rect 5251 70291 5309 70297
rect 4876 70202 7912 70224
rect 4876 70150 6690 70202
rect 6742 70150 6754 70202
rect 6806 70150 6818 70202
rect 6870 70150 6882 70202
rect 6934 70150 6946 70202
rect 6998 70150 7912 70202
rect 4876 70128 7912 70150
rect 86020 70202 88964 70224
rect 86020 70150 87834 70202
rect 87886 70150 87898 70202
rect 87950 70150 87962 70202
rect 88014 70150 88026 70202
rect 88078 70150 88090 70202
rect 88142 70150 88964 70202
rect 86020 70128 88964 70150
rect 5457 69957 5515 69963
rect 5457 69923 5469 69957
rect 5503 69954 5515 69957
rect 5503 69926 5800 69954
rect 88554 69948 88560 70000
rect 88612 69948 88618 70000
rect 5503 69923 5515 69926
rect 5457 69917 5515 69923
rect 5772 69920 5800 69926
rect 7134 69920 7140 69932
rect 5772 69892 7140 69920
rect 7134 69880 7140 69892
rect 7192 69880 7198 69932
rect 84322 69812 84328 69864
rect 84380 69852 84386 69864
rect 88327 69855 88385 69861
rect 88327 69852 88339 69855
rect 84380 69824 88339 69852
rect 84380 69812 84386 69824
rect 88327 69821 88339 69824
rect 88373 69821 88385 69855
rect 88327 69815 88385 69821
rect 2902 69744 2908 69796
rect 2960 69784 2966 69796
rect 5251 69787 5309 69793
rect 5251 69784 5263 69787
rect 2960 69756 5263 69784
rect 2960 69744 2966 69756
rect 5251 69753 5263 69756
rect 5297 69753 5309 69787
rect 5251 69747 5309 69753
rect 4876 69658 7912 69680
rect 4876 69606 5954 69658
rect 6006 69606 6018 69658
rect 6070 69606 6082 69658
rect 6134 69606 6146 69658
rect 6198 69606 6210 69658
rect 6262 69606 7912 69658
rect 4876 69584 7912 69606
rect 86020 69658 88964 69680
rect 86020 69606 87098 69658
rect 87150 69606 87162 69658
rect 87214 69606 87226 69658
rect 87278 69606 87290 69658
rect 87342 69606 87354 69658
rect 87406 69606 88964 69658
rect 86020 69584 88964 69606
rect 88465 69311 88523 69317
rect 88465 69277 88477 69311
rect 88511 69308 88523 69311
rect 89934 69308 89940 69320
rect 88511 69280 89940 69308
rect 88511 69277 88523 69280
rect 88465 69271 88523 69277
rect 89934 69268 89940 69280
rect 89992 69268 89998 69320
rect 4876 69114 7912 69136
rect 4876 69062 6690 69114
rect 6742 69062 6754 69114
rect 6806 69062 6818 69114
rect 6870 69062 6882 69114
rect 6934 69062 6946 69114
rect 6998 69062 7912 69114
rect 4876 69040 7912 69062
rect 86020 69114 88964 69136
rect 86020 69062 87834 69114
rect 87886 69062 87898 69114
rect 87950 69062 87962 69114
rect 88014 69062 88026 69114
rect 88078 69062 88090 69114
rect 88142 69062 88964 69114
rect 86020 69040 88964 69062
rect 88646 68875 88652 68878
rect 5457 68869 5515 68875
rect 5457 68835 5469 68869
rect 5503 68866 5515 68869
rect 88621 68869 88652 68875
rect 5503 68838 5800 68866
rect 5503 68835 5515 68838
rect 5457 68829 5515 68835
rect 5772 68832 5800 68838
rect 7134 68832 7140 68844
rect 5772 68804 7140 68832
rect 7134 68792 7140 68804
rect 7192 68792 7198 68844
rect 88621 68835 88633 68869
rect 88621 68829 88652 68835
rect 88646 68826 88652 68829
rect 88704 68826 88710 68878
rect 2902 68656 2908 68708
rect 2960 68696 2966 68708
rect 5251 68699 5309 68705
rect 5251 68696 5263 68699
rect 2960 68668 5263 68696
rect 2960 68656 2966 68668
rect 5251 68665 5263 68668
rect 5297 68665 5309 68699
rect 5251 68659 5309 68665
rect 84322 68656 84328 68708
rect 84380 68696 84386 68708
rect 88419 68699 88477 68705
rect 88419 68696 88431 68699
rect 84380 68668 88431 68696
rect 84380 68656 84386 68668
rect 88419 68665 88431 68668
rect 88465 68665 88477 68699
rect 88419 68659 88477 68665
rect 4876 68570 7912 68592
rect 4876 68518 5954 68570
rect 6006 68518 6018 68570
rect 6070 68518 6082 68570
rect 6134 68518 6146 68570
rect 6198 68518 6210 68570
rect 6262 68518 7912 68570
rect 4876 68496 7912 68518
rect 86020 68570 88964 68592
rect 86020 68518 87098 68570
rect 87150 68518 87162 68570
rect 87214 68518 87226 68570
rect 87278 68518 87290 68570
rect 87342 68518 87354 68570
rect 87406 68518 88964 68570
rect 86020 68496 88964 68518
rect 4876 68026 7912 68048
rect 4876 67974 6690 68026
rect 6742 67974 6754 68026
rect 6806 67974 6818 68026
rect 6870 67974 6882 68026
rect 6934 67974 6946 68026
rect 6998 67974 7912 68026
rect 4876 67952 7912 67974
rect 86020 68026 88964 68048
rect 86020 67974 87834 68026
rect 87886 67974 87898 68026
rect 87950 67974 87962 68026
rect 88014 67974 88026 68026
rect 88078 67974 88090 68026
rect 88142 67974 88964 68026
rect 86020 67952 88964 67974
rect 88646 67787 88652 67790
rect 5457 67781 5515 67787
rect 5457 67747 5469 67781
rect 5503 67778 5515 67781
rect 88621 67781 88652 67787
rect 5503 67750 5800 67778
rect 5503 67747 5515 67750
rect 5457 67741 5515 67747
rect 5772 67744 5800 67750
rect 7134 67744 7140 67756
rect 5772 67716 7140 67744
rect 7134 67704 7140 67716
rect 7192 67704 7198 67756
rect 88621 67747 88633 67781
rect 88621 67741 88652 67747
rect 88646 67738 88652 67741
rect 88704 67738 88710 67790
rect 2902 67568 2908 67620
rect 2960 67608 2966 67620
rect 5251 67611 5309 67617
rect 5251 67608 5263 67611
rect 2960 67580 5263 67608
rect 2960 67568 2966 67580
rect 5251 67577 5263 67580
rect 5297 67577 5309 67611
rect 5251 67571 5309 67577
rect 84322 67568 84328 67620
rect 84380 67608 84386 67620
rect 88419 67611 88477 67617
rect 88419 67608 88431 67611
rect 84380 67580 88431 67608
rect 84380 67568 84386 67580
rect 88419 67577 88431 67580
rect 88465 67577 88477 67611
rect 88419 67571 88477 67577
rect 4876 67482 7912 67504
rect 4876 67430 5954 67482
rect 6006 67430 6018 67482
rect 6070 67430 6082 67482
rect 6134 67430 6146 67482
rect 6198 67430 6210 67482
rect 6262 67430 7912 67482
rect 4876 67408 7912 67430
rect 86020 67482 88964 67504
rect 86020 67430 87098 67482
rect 87150 67430 87162 67482
rect 87214 67430 87226 67482
rect 87278 67430 87290 67482
rect 87342 67430 87354 67482
rect 87406 67430 88964 67482
rect 86020 67408 88964 67430
rect 4876 66938 7912 66960
rect 4876 66886 6690 66938
rect 6742 66886 6754 66938
rect 6806 66886 6818 66938
rect 6870 66886 6882 66938
rect 6934 66886 6946 66938
rect 6998 66886 7912 66938
rect 4876 66864 7912 66886
rect 86020 66938 88964 66960
rect 86020 66886 87834 66938
rect 87886 66886 87898 66938
rect 87950 66886 87962 66938
rect 88014 66886 88026 66938
rect 88078 66886 88090 66938
rect 88142 66886 88964 66938
rect 86020 66864 88964 66886
rect 5478 66699 5484 66702
rect 5457 66693 5484 66699
rect 5457 66659 5469 66693
rect 5457 66653 5484 66659
rect 5478 66650 5484 66653
rect 5536 66650 5542 66702
rect 88603 66675 88661 66681
rect 88603 66641 88615 66675
rect 88649 66672 88661 66675
rect 88649 66656 88876 66672
rect 90118 66656 90124 66668
rect 88649 66644 90124 66656
rect 88649 66641 88661 66644
rect 88603 66635 88661 66641
rect 88848 66628 90124 66644
rect 90118 66616 90124 66628
rect 90176 66616 90182 66668
rect 4374 66480 4380 66532
rect 4432 66520 4438 66532
rect 5251 66523 5309 66529
rect 5251 66520 5263 66523
rect 4432 66492 5263 66520
rect 4432 66480 4438 66492
rect 5251 66489 5263 66492
rect 5297 66489 5309 66523
rect 5251 66483 5309 66489
rect 87450 66480 87456 66532
rect 87508 66520 87514 66532
rect 88419 66523 88477 66529
rect 88419 66520 88431 66523
rect 87508 66492 88431 66520
rect 87508 66480 87514 66492
rect 88419 66489 88431 66492
rect 88465 66489 88477 66523
rect 88419 66483 88477 66489
rect 4876 66394 7912 66416
rect 4876 66342 5954 66394
rect 6006 66342 6018 66394
rect 6070 66342 6082 66394
rect 6134 66342 6146 66394
rect 6198 66342 6210 66394
rect 6262 66342 7912 66394
rect 4876 66320 7912 66342
rect 86020 66394 88964 66416
rect 86020 66342 87098 66394
rect 87150 66342 87162 66394
rect 87214 66342 87226 66394
rect 87278 66342 87290 66394
rect 87342 66342 87354 66394
rect 87406 66342 88964 66394
rect 86020 66320 88964 66342
rect 4876 65850 7912 65872
rect 4876 65798 6690 65850
rect 6742 65798 6754 65850
rect 6806 65798 6818 65850
rect 6870 65798 6882 65850
rect 6934 65798 6946 65850
rect 6998 65798 7912 65850
rect 4876 65776 7912 65798
rect 86020 65850 88964 65872
rect 86020 65798 87834 65850
rect 87886 65798 87898 65850
rect 87950 65798 87962 65850
rect 88014 65798 88026 65850
rect 88078 65798 88090 65850
rect 88142 65798 88964 65850
rect 86020 65776 88964 65798
rect 4876 65306 7912 65328
rect 4876 65254 5954 65306
rect 6006 65254 6018 65306
rect 6070 65254 6082 65306
rect 6134 65254 6146 65306
rect 6198 65254 6210 65306
rect 6262 65254 7912 65306
rect 4876 65232 7912 65254
rect 86020 65306 88964 65328
rect 86020 65254 87098 65306
rect 87150 65254 87162 65306
rect 87214 65254 87226 65306
rect 87278 65254 87290 65306
rect 87342 65254 87354 65306
rect 87406 65254 88964 65306
rect 86020 65232 88964 65254
rect 5386 65101 5392 65104
rect 5364 65095 5392 65101
rect 5364 65061 5376 65095
rect 5364 65055 5392 65061
rect 5386 65052 5392 65055
rect 5444 65052 5450 65104
rect 5159 64993 5217 64999
rect 5159 64990 5171 64993
rect 2902 64916 2908 64968
rect 2960 64956 2966 64968
rect 4852 64962 5171 64990
rect 4852 64956 4880 64962
rect 2960 64928 4880 64956
rect 5159 64959 5171 64962
rect 5205 64959 5217 64993
rect 84322 64984 84328 65036
rect 84380 65024 84386 65036
rect 84380 64996 87956 65024
rect 84380 64984 84386 64996
rect 87928 64990 87956 64996
rect 88233 64993 88291 64999
rect 88233 64990 88245 64993
rect 87928 64962 88245 64990
rect 5159 64953 5217 64959
rect 88233 64959 88245 64962
rect 88279 64959 88291 64993
rect 88233 64953 88291 64959
rect 2960 64916 2966 64928
rect 88445 64891 88503 64897
rect 88445 64857 88457 64891
rect 88491 64888 88503 64891
rect 89934 64888 89940 64900
rect 88491 64860 89940 64888
rect 88491 64857 88503 64860
rect 88445 64851 88503 64857
rect 89934 64848 89940 64860
rect 89992 64848 89998 64900
rect 4876 64762 7912 64784
rect 4876 64710 6690 64762
rect 6742 64710 6754 64762
rect 6806 64710 6818 64762
rect 6870 64710 6882 64762
rect 6934 64710 6946 64762
rect 6998 64710 7912 64762
rect 4876 64688 7912 64710
rect 86020 64762 88964 64784
rect 86020 64710 87834 64762
rect 87886 64710 87898 64762
rect 87950 64710 87962 64762
rect 88014 64710 88026 64762
rect 88078 64710 88090 64762
rect 88142 64710 88964 64762
rect 86020 64688 88964 64710
rect 5159 64517 5217 64523
rect 5159 64514 5171 64517
rect 2902 64440 2908 64492
rect 2960 64480 2966 64492
rect 4852 64486 5171 64514
rect 4852 64480 4880 64486
rect 2960 64452 4880 64480
rect 5159 64483 5171 64486
rect 5205 64483 5217 64517
rect 88325 64517 88383 64523
rect 88325 64514 88337 64517
rect 5159 64477 5217 64483
rect 2960 64440 2966 64452
rect 84322 64440 84328 64492
rect 84380 64480 84386 64492
rect 88020 64486 88337 64514
rect 88020 64480 88048 64486
rect 84380 64452 88048 64480
rect 88325 64483 88337 64486
rect 88371 64483 88383 64517
rect 88325 64477 88383 64483
rect 84380 64440 84386 64452
rect 5364 64347 5422 64353
rect 5364 64313 5376 64347
rect 5410 64344 5422 64347
rect 7226 64344 7232 64356
rect 5410 64316 7232 64344
rect 5410 64313 5422 64316
rect 5364 64307 5422 64313
rect 7226 64304 7232 64316
rect 7284 64304 7290 64356
rect 88554 64353 88560 64356
rect 88537 64347 88560 64353
rect 88537 64313 88549 64347
rect 88537 64307 88560 64313
rect 88554 64304 88560 64307
rect 88612 64304 88618 64356
rect 4876 64218 7912 64240
rect 4876 64166 5954 64218
rect 6006 64166 6018 64218
rect 6070 64166 6082 64218
rect 6134 64166 6146 64218
rect 6198 64166 6210 64218
rect 6262 64166 7912 64218
rect 4876 64144 7912 64166
rect 86020 64218 88964 64240
rect 86020 64166 87098 64218
rect 87150 64166 87162 64218
rect 87214 64166 87226 64218
rect 87278 64166 87290 64218
rect 87342 64166 87354 64218
rect 87406 64166 88964 64218
rect 86020 64144 88964 64166
rect 4876 63674 7912 63696
rect 4876 63622 6690 63674
rect 6742 63622 6754 63674
rect 6806 63622 6818 63674
rect 6870 63622 6882 63674
rect 6934 63622 6946 63674
rect 6998 63622 7912 63674
rect 4876 63600 7912 63622
rect 86020 63674 88964 63696
rect 86020 63622 87834 63674
rect 87886 63622 87898 63674
rect 87950 63622 87962 63674
rect 88014 63622 88026 63674
rect 88078 63622 88090 63674
rect 88142 63622 88964 63674
rect 86020 63600 88964 63622
rect 5159 63429 5217 63435
rect 5159 63426 5171 63429
rect 2902 63352 2908 63404
rect 2960 63392 2966 63404
rect 4852 63398 5171 63426
rect 4852 63392 4880 63398
rect 2960 63364 4880 63392
rect 5159 63395 5171 63398
rect 5205 63395 5217 63429
rect 88325 63429 88383 63435
rect 88325 63426 88337 63429
rect 5159 63389 5217 63395
rect 2960 63352 2966 63364
rect 84322 63352 84328 63404
rect 84380 63392 84386 63404
rect 88020 63398 88337 63426
rect 88020 63392 88048 63398
rect 84380 63364 88048 63392
rect 88325 63395 88337 63398
rect 88371 63395 88383 63429
rect 88325 63389 88383 63395
rect 84380 63352 84386 63364
rect 5364 63259 5422 63265
rect 5364 63225 5376 63259
rect 5410 63256 5422 63259
rect 7226 63256 7232 63268
rect 5410 63228 7232 63256
rect 5410 63225 5422 63228
rect 5364 63219 5422 63225
rect 7226 63216 7232 63228
rect 7284 63216 7290 63268
rect 88554 63265 88560 63268
rect 88537 63259 88560 63265
rect 88537 63225 88549 63259
rect 88537 63219 88560 63225
rect 88554 63216 88560 63219
rect 88612 63216 88618 63268
rect 4876 63130 7912 63152
rect 4876 63078 5954 63130
rect 6006 63078 6018 63130
rect 6070 63078 6082 63130
rect 6134 63078 6146 63130
rect 6198 63078 6210 63130
rect 6262 63078 7912 63130
rect 4876 63056 7912 63078
rect 86020 63130 88964 63152
rect 86020 63078 87098 63130
rect 87150 63078 87162 63130
rect 87214 63078 87226 63130
rect 87278 63078 87290 63130
rect 87342 63078 87354 63130
rect 87406 63078 88964 63130
rect 86020 63056 88964 63078
rect 4876 62586 7912 62608
rect 4876 62534 6690 62586
rect 6742 62534 6754 62586
rect 6806 62534 6818 62586
rect 6870 62534 6882 62586
rect 6934 62534 6946 62586
rect 6998 62534 7912 62586
rect 4876 62512 7912 62534
rect 86020 62586 88964 62608
rect 86020 62534 87834 62586
rect 87886 62534 87898 62586
rect 87950 62534 87962 62586
rect 88014 62534 88026 62586
rect 88078 62534 88090 62586
rect 88142 62534 88964 62586
rect 86020 62512 88964 62534
rect 5364 62375 5422 62381
rect 5202 62298 5208 62350
rect 5260 62298 5266 62350
rect 5364 62341 5376 62375
rect 5410 62372 5422 62375
rect 9618 62372 9624 62384
rect 5410 62344 9624 62372
rect 5410 62341 5422 62344
rect 5364 62335 5422 62341
rect 9618 62332 9624 62344
rect 9676 62332 9682 62384
rect 88537 62375 88595 62381
rect 88370 62298 88376 62350
rect 88428 62298 88434 62350
rect 88537 62341 88549 62375
rect 88583 62372 88595 62375
rect 89934 62372 89940 62384
rect 88583 62344 89940 62372
rect 88583 62341 88595 62344
rect 88537 62335 88595 62341
rect 89934 62332 89940 62344
rect 89992 62332 89998 62384
rect 4876 62042 7912 62064
rect 4876 61990 5954 62042
rect 6006 61990 6018 62042
rect 6070 61990 6082 62042
rect 6134 61990 6146 62042
rect 6198 61990 6210 62042
rect 6262 61990 7912 62042
rect 4876 61968 7912 61990
rect 86020 62042 88964 62064
rect 86020 61990 87098 62042
rect 87150 61990 87162 62042
rect 87214 61990 87226 62042
rect 87278 61990 87290 62042
rect 87342 61990 87354 62042
rect 87406 61990 88964 62042
rect 86020 61968 88964 61990
rect 4876 61498 7912 61520
rect 4876 61446 6690 61498
rect 6742 61446 6754 61498
rect 6806 61446 6818 61498
rect 6870 61446 6882 61498
rect 6934 61446 6946 61498
rect 6998 61446 7912 61498
rect 4876 61424 7912 61446
rect 86020 61498 88964 61520
rect 86020 61446 87834 61498
rect 87886 61446 87898 61498
rect 87950 61446 87962 61498
rect 88014 61446 88026 61498
rect 88078 61446 88090 61498
rect 88142 61446 88964 61498
rect 86020 61424 88964 61446
rect 5202 61210 5208 61262
rect 5260 61210 5266 61262
rect 88370 61210 88376 61262
rect 88428 61210 88434 61262
rect 5364 61083 5422 61089
rect 5364 61049 5376 61083
rect 5410 61080 5422 61083
rect 9618 61080 9624 61092
rect 5410 61052 9624 61080
rect 5410 61049 5422 61052
rect 5364 61043 5422 61049
rect 9618 61040 9624 61052
rect 9676 61040 9682 61092
rect 88537 61083 88595 61089
rect 88537 61049 88549 61083
rect 88583 61080 88595 61083
rect 89934 61080 89940 61092
rect 88583 61052 89940 61080
rect 88583 61049 88595 61052
rect 88537 61043 88595 61049
rect 89934 61040 89940 61052
rect 89992 61040 89998 61092
rect 4876 60954 7912 60976
rect 4876 60902 5954 60954
rect 6006 60902 6018 60954
rect 6070 60902 6082 60954
rect 6134 60902 6146 60954
rect 6198 60902 6210 60954
rect 6262 60902 7912 60954
rect 4876 60880 7912 60902
rect 86020 60954 88964 60976
rect 86020 60902 87098 60954
rect 87150 60902 87162 60954
rect 87214 60902 87226 60954
rect 87278 60902 87290 60954
rect 87342 60902 87354 60954
rect 87406 60902 88964 60954
rect 86020 60880 88964 60902
rect 4876 60410 7912 60432
rect 4876 60358 6690 60410
rect 6742 60358 6754 60410
rect 6806 60358 6818 60410
rect 6870 60358 6882 60410
rect 6934 60358 6946 60410
rect 6998 60358 7912 60410
rect 4876 60336 7912 60358
rect 86020 60410 88964 60432
rect 86020 60358 87834 60410
rect 87886 60358 87898 60410
rect 87950 60358 87962 60410
rect 88014 60358 88026 60410
rect 88078 60358 88090 60410
rect 88142 60358 88964 60410
rect 86020 60336 88964 60358
rect 4876 59866 7912 59888
rect 4876 59814 5954 59866
rect 6006 59814 6018 59866
rect 6070 59814 6082 59866
rect 6134 59814 6146 59866
rect 6198 59814 6210 59866
rect 6262 59814 7912 59866
rect 4876 59792 7912 59814
rect 86020 59866 88964 59888
rect 86020 59814 87098 59866
rect 87150 59814 87162 59866
rect 87214 59814 87226 59866
rect 87278 59814 87290 59866
rect 87342 59814 87354 59866
rect 87406 59814 88964 59866
rect 86020 59792 88964 59814
rect 5159 59553 5217 59559
rect 5159 59550 5171 59553
rect 2902 59476 2908 59528
rect 2960 59516 2966 59528
rect 4852 59522 5171 59550
rect 4852 59516 4880 59522
rect 2960 59488 4880 59516
rect 5159 59519 5171 59522
rect 5205 59519 5217 59553
rect 88233 59553 88291 59559
rect 88233 59550 88245 59553
rect 5159 59513 5217 59519
rect 5364 59519 5422 59525
rect 2960 59476 2966 59488
rect 5364 59485 5376 59519
rect 5410 59516 5422 59519
rect 5662 59516 5668 59528
rect 5410 59488 5668 59516
rect 5410 59485 5422 59488
rect 5364 59479 5422 59485
rect 5662 59476 5668 59488
rect 5720 59476 5726 59528
rect 84322 59476 84328 59528
rect 84380 59516 84386 59528
rect 87928 59522 88245 59550
rect 87928 59516 87956 59522
rect 84380 59488 87956 59516
rect 88233 59519 88245 59522
rect 88279 59519 88291 59553
rect 88233 59513 88291 59519
rect 84380 59476 84386 59488
rect 88445 59451 88503 59457
rect 88445 59417 88457 59451
rect 88491 59448 88503 59451
rect 89934 59448 89940 59460
rect 88491 59420 89940 59448
rect 88491 59417 88503 59420
rect 88445 59411 88503 59417
rect 89934 59408 89940 59420
rect 89992 59408 89998 59460
rect 4876 59322 7912 59344
rect 4876 59270 6690 59322
rect 6742 59270 6754 59322
rect 6806 59270 6818 59322
rect 6870 59270 6882 59322
rect 6934 59270 6946 59322
rect 6998 59270 7912 59322
rect 4876 59248 7912 59270
rect 86020 59322 88964 59344
rect 86020 59270 87834 59322
rect 87886 59270 87898 59322
rect 87950 59270 87962 59322
rect 88014 59270 88026 59322
rect 88078 59270 88090 59322
rect 88142 59270 88964 59322
rect 86020 59248 88964 59270
rect 5159 59077 5217 59083
rect 5159 59074 5171 59077
rect 2902 59000 2908 59052
rect 2960 59040 2966 59052
rect 4852 59046 5171 59074
rect 4852 59040 4880 59046
rect 2960 59012 4880 59040
rect 5159 59043 5171 59046
rect 5205 59043 5217 59077
rect 88325 59077 88383 59083
rect 88325 59074 88337 59077
rect 5159 59037 5217 59043
rect 2960 59000 2966 59012
rect 84322 59000 84328 59052
rect 84380 59040 84386 59052
rect 88020 59046 88337 59074
rect 88020 59040 88048 59046
rect 84380 59012 88048 59040
rect 88325 59043 88337 59046
rect 88371 59043 88383 59077
rect 88325 59037 88383 59043
rect 84380 59000 84386 59012
rect 5364 58907 5422 58913
rect 5364 58873 5376 58907
rect 5410 58904 5422 58907
rect 7226 58904 7232 58916
rect 5410 58876 7232 58904
rect 5410 58873 5422 58876
rect 5364 58867 5422 58873
rect 7226 58864 7232 58876
rect 7284 58864 7290 58916
rect 88554 58913 88560 58916
rect 88537 58907 88560 58913
rect 88537 58873 88549 58907
rect 88537 58867 88560 58873
rect 88554 58864 88560 58867
rect 88612 58864 88618 58916
rect 4876 58778 7912 58800
rect 4876 58726 5954 58778
rect 6006 58726 6018 58778
rect 6070 58726 6082 58778
rect 6134 58726 6146 58778
rect 6198 58726 6210 58778
rect 6262 58726 7912 58778
rect 4876 58704 7912 58726
rect 86020 58778 88964 58800
rect 86020 58726 87098 58778
rect 87150 58726 87162 58778
rect 87214 58726 87226 58778
rect 87278 58726 87290 58778
rect 87342 58726 87354 58778
rect 87406 58726 88964 58778
rect 86020 58704 88964 58726
rect 4876 58234 7912 58256
rect 4876 58182 6690 58234
rect 6742 58182 6754 58234
rect 6806 58182 6818 58234
rect 6870 58182 6882 58234
rect 6934 58182 6946 58234
rect 6998 58182 7912 58234
rect 4876 58160 7912 58182
rect 86020 58234 88964 58256
rect 86020 58182 87834 58234
rect 87886 58182 87898 58234
rect 87950 58182 87962 58234
rect 88014 58182 88026 58234
rect 88078 58182 88090 58234
rect 88142 58182 88964 58234
rect 86020 58160 88964 58182
rect 5159 57989 5217 57995
rect 5159 57986 5171 57989
rect 2902 57912 2908 57964
rect 2960 57952 2966 57964
rect 4852 57958 5171 57986
rect 4852 57952 4880 57958
rect 2960 57924 4880 57952
rect 5159 57955 5171 57958
rect 5205 57955 5217 57989
rect 88325 57989 88383 57995
rect 88325 57986 88337 57989
rect 5159 57949 5217 57955
rect 2960 57912 2966 57924
rect 84322 57912 84328 57964
rect 84380 57952 84386 57964
rect 88020 57958 88337 57986
rect 88020 57952 88048 57958
rect 84380 57924 88048 57952
rect 88325 57955 88337 57958
rect 88371 57955 88383 57989
rect 88325 57949 88383 57955
rect 84380 57912 84386 57924
rect 5364 57819 5422 57825
rect 5364 57785 5376 57819
rect 5410 57816 5422 57819
rect 7226 57816 7232 57828
rect 5410 57788 7232 57816
rect 5410 57785 5422 57788
rect 5364 57779 5422 57785
rect 7226 57776 7232 57788
rect 7284 57776 7290 57828
rect 88554 57825 88560 57828
rect 88537 57819 88560 57825
rect 88537 57785 88549 57819
rect 88537 57779 88560 57785
rect 88554 57776 88560 57779
rect 88612 57776 88618 57828
rect 4876 57690 7912 57712
rect 4876 57638 5954 57690
rect 6006 57638 6018 57690
rect 6070 57638 6082 57690
rect 6134 57638 6146 57690
rect 6198 57638 6210 57690
rect 6262 57638 7912 57690
rect 4876 57616 7912 57638
rect 86020 57690 88964 57712
rect 86020 57638 87098 57690
rect 87150 57638 87162 57690
rect 87214 57638 87226 57690
rect 87278 57638 87290 57690
rect 87342 57638 87354 57690
rect 87406 57638 88964 57690
rect 86020 57616 88964 57638
rect 4876 57146 7912 57168
rect 4876 57094 6690 57146
rect 6742 57094 6754 57146
rect 6806 57094 6818 57146
rect 6870 57094 6882 57146
rect 6934 57094 6946 57146
rect 6998 57094 7912 57146
rect 4876 57072 7912 57094
rect 86020 57146 88964 57168
rect 86020 57094 87834 57146
rect 87886 57094 87898 57146
rect 87950 57094 87962 57146
rect 88014 57094 88026 57146
rect 88078 57094 88090 57146
rect 88142 57094 88964 57146
rect 86020 57072 88964 57094
rect 4926 56858 4932 56910
rect 4984 56898 4990 56910
rect 5159 56901 5217 56907
rect 5159 56898 5171 56901
rect 4984 56870 5171 56898
rect 4984 56858 4990 56870
rect 5159 56867 5171 56870
rect 5205 56867 5217 56901
rect 5386 56873 5392 56876
rect 5159 56861 5217 56867
rect 5364 56867 5392 56873
rect 5364 56833 5376 56867
rect 5364 56827 5392 56833
rect 5386 56824 5392 56827
rect 5444 56824 5450 56876
rect 88278 56858 88284 56910
rect 88336 56898 88342 56910
rect 88373 56901 88431 56907
rect 88373 56898 88385 56901
rect 88336 56870 88385 56898
rect 88336 56858 88342 56870
rect 88373 56867 88385 56870
rect 88419 56867 88431 56901
rect 88373 56861 88431 56867
rect 88537 56867 88595 56873
rect 88537 56833 88549 56867
rect 88583 56864 88595 56867
rect 89934 56864 89940 56876
rect 88583 56836 89940 56864
rect 88583 56833 88595 56836
rect 88537 56827 88595 56833
rect 89934 56824 89940 56836
rect 89992 56824 89998 56876
rect 4876 56602 7912 56624
rect 4876 56550 5954 56602
rect 6006 56550 6018 56602
rect 6070 56550 6082 56602
rect 6134 56550 6146 56602
rect 6198 56550 6210 56602
rect 6262 56550 7912 56602
rect 4876 56528 7912 56550
rect 86020 56602 88964 56624
rect 86020 56550 87098 56602
rect 87150 56550 87162 56602
rect 87214 56550 87226 56602
rect 87278 56550 87290 56602
rect 87342 56550 87354 56602
rect 87406 56550 88964 56602
rect 86020 56528 88964 56550
rect 4876 56058 7912 56080
rect 4876 56006 6690 56058
rect 6742 56006 6754 56058
rect 6806 56006 6818 56058
rect 6870 56006 6882 56058
rect 6934 56006 6946 56058
rect 6998 56006 7912 56058
rect 4876 55984 7912 56006
rect 86020 56058 88964 56080
rect 86020 56006 87834 56058
rect 87886 56006 87898 56058
rect 87950 56006 87962 56058
rect 88014 56006 88026 56058
rect 88078 56006 88090 56058
rect 88142 56006 88964 56058
rect 86020 55984 88964 56006
rect 5018 55770 5024 55822
rect 5076 55810 5082 55822
rect 5159 55813 5217 55819
rect 5159 55810 5171 55813
rect 5076 55782 5171 55810
rect 5076 55770 5082 55782
rect 5159 55779 5171 55782
rect 5205 55779 5217 55813
rect 5159 55773 5217 55779
rect 88370 55770 88376 55822
rect 88428 55770 88434 55822
rect 5364 55643 5422 55649
rect 5364 55609 5376 55643
rect 5410 55640 5422 55643
rect 5662 55640 5668 55652
rect 5410 55612 5668 55640
rect 5410 55609 5422 55612
rect 5364 55603 5422 55609
rect 5662 55600 5668 55612
rect 5720 55600 5726 55652
rect 88537 55643 88595 55649
rect 88537 55609 88549 55643
rect 88583 55640 88595 55643
rect 89934 55640 89940 55652
rect 88583 55612 89940 55640
rect 88583 55609 88595 55612
rect 88537 55603 88595 55609
rect 89934 55600 89940 55612
rect 89992 55600 89998 55652
rect 4876 55514 7912 55536
rect 4876 55462 5954 55514
rect 6006 55462 6018 55514
rect 6070 55462 6082 55514
rect 6134 55462 6146 55514
rect 6198 55462 6210 55514
rect 6262 55462 7912 55514
rect 4876 55440 7912 55462
rect 86020 55514 88964 55536
rect 86020 55462 87098 55514
rect 87150 55462 87162 55514
rect 87214 55462 87226 55514
rect 87278 55462 87290 55514
rect 87342 55462 87354 55514
rect 87406 55462 88964 55514
rect 86020 55440 88964 55462
rect 2534 55124 2540 55176
rect 2592 55164 2598 55176
rect 5205 55167 5263 55173
rect 5205 55164 5217 55167
rect 2592 55136 5217 55164
rect 2592 55124 2598 55136
rect 5205 55133 5217 55136
rect 5251 55133 5263 55167
rect 5205 55127 5263 55133
rect 4876 54970 7912 54992
rect 4876 54918 6690 54970
rect 6742 54918 6754 54970
rect 6806 54918 6818 54970
rect 6870 54918 6882 54970
rect 6934 54918 6946 54970
rect 6998 54918 7912 54970
rect 4876 54896 7912 54918
rect 86020 54970 88964 54992
rect 86020 54918 87834 54970
rect 87886 54918 87898 54970
rect 87950 54918 87962 54970
rect 88014 54918 88026 54970
rect 88078 54918 88090 54970
rect 88142 54918 88964 54970
rect 86020 54896 88964 54918
rect 7594 54765 7600 54768
rect 7573 54759 7600 54765
rect 7573 54725 7585 54759
rect 7573 54719 7600 54725
rect 7594 54716 7600 54719
rect 7652 54716 7658 54768
rect 6953 54555 7011 54561
rect 6953 54521 6965 54555
rect 6999 54552 7011 54555
rect 7042 54552 7048 54564
rect 6999 54524 7048 54552
rect 6999 54521 7011 54524
rect 6953 54515 7011 54521
rect 7042 54512 7048 54524
rect 7100 54512 7106 54564
rect 4876 54426 7912 54448
rect 4876 54374 5954 54426
rect 6006 54374 6018 54426
rect 6070 54374 6082 54426
rect 6134 54374 6146 54426
rect 6198 54374 6210 54426
rect 6262 54374 7912 54426
rect 4876 54352 7912 54374
rect 86020 54426 88964 54448
rect 86020 54374 87098 54426
rect 87150 54374 87162 54426
rect 87214 54374 87226 54426
rect 87278 54374 87290 54426
rect 87342 54374 87354 54426
rect 87406 54374 88964 54426
rect 86020 54352 88964 54374
rect 84322 54104 84328 54156
rect 84380 54144 84386 54156
rect 84380 54116 87956 54144
rect 84380 54104 84386 54116
rect 87928 54110 87956 54116
rect 88233 54113 88291 54119
rect 88233 54110 88245 54113
rect 5202 54036 5208 54088
rect 5260 54036 5266 54088
rect 87928 54082 88245 54110
rect 88233 54079 88245 54082
rect 88279 54079 88291 54113
rect 88233 54073 88291 54079
rect 88445 54079 88503 54085
rect 88445 54045 88457 54079
rect 88491 54076 88503 54079
rect 89934 54076 89940 54088
rect 88491 54048 89940 54076
rect 88491 54045 88503 54048
rect 88445 54039 88503 54045
rect 89934 54036 89940 54048
rect 89992 54036 89998 54088
rect 4876 53882 7912 53904
rect 4876 53830 6690 53882
rect 6742 53830 6754 53882
rect 6806 53830 6818 53882
rect 6870 53830 6882 53882
rect 6934 53830 6946 53882
rect 6998 53830 7912 53882
rect 4876 53808 7912 53830
rect 86020 53882 88964 53904
rect 86020 53830 87834 53882
rect 87886 53830 87898 53882
rect 87950 53830 87962 53882
rect 88014 53830 88026 53882
rect 88078 53830 88090 53882
rect 88142 53830 88964 53882
rect 86020 53808 88964 53830
rect 5364 53739 5422 53745
rect 5364 53705 5376 53739
rect 5410 53736 5422 53739
rect 5662 53736 5668 53748
rect 5410 53708 5668 53736
rect 5410 53705 5422 53708
rect 5364 53699 5422 53705
rect 5662 53696 5668 53708
rect 5720 53696 5726 53748
rect 5159 53637 5217 53643
rect 2902 53560 2908 53612
rect 2960 53600 2966 53612
rect 5159 53603 5171 53637
rect 5205 53603 5217 53637
rect 88325 53637 88383 53643
rect 88325 53634 88337 53637
rect 5159 53600 5217 53603
rect 2960 53597 5217 53600
rect 2960 53572 5202 53597
rect 2960 53560 2966 53572
rect 84322 53560 84328 53612
rect 84380 53600 84386 53612
rect 88020 53606 88337 53634
rect 88020 53600 88048 53606
rect 84380 53572 88048 53600
rect 88325 53603 88337 53606
rect 88371 53603 88383 53637
rect 88325 53597 88383 53603
rect 84380 53560 84386 53572
rect 88554 53473 88560 53476
rect 88537 53467 88560 53473
rect 88537 53433 88549 53467
rect 88537 53427 88560 53433
rect 88554 53424 88560 53427
rect 88612 53424 88618 53476
rect 4876 53338 7912 53360
rect 4876 53286 5954 53338
rect 6006 53286 6018 53338
rect 6070 53286 6082 53338
rect 6134 53286 6146 53338
rect 6198 53286 6210 53338
rect 6262 53286 7912 53338
rect 4876 53264 7912 53286
rect 86020 53338 88964 53360
rect 86020 53286 87098 53338
rect 87150 53286 87162 53338
rect 87214 53286 87226 53338
rect 87278 53286 87290 53338
rect 87342 53286 87354 53338
rect 87406 53286 88964 53338
rect 86020 53264 88964 53286
rect 5365 53195 5423 53201
rect 5365 53161 5377 53195
rect 5411 53192 5423 53195
rect 7134 53192 7140 53204
rect 5411 53164 7140 53192
rect 5411 53161 5423 53164
rect 5365 53155 5423 53161
rect 7134 53152 7140 53164
rect 7192 53152 7198 53204
rect 5159 53025 5217 53031
rect 2902 52948 2908 53000
rect 2960 52988 2966 53000
rect 5159 52991 5171 53025
rect 5205 52991 5217 53025
rect 5159 52988 5217 52991
rect 2960 52985 5217 52988
rect 88465 52991 88523 52997
rect 2960 52960 5202 52985
rect 2960 52948 2966 52960
rect 88465 52957 88477 52991
rect 88511 52988 88523 52991
rect 89934 52988 89940 53000
rect 88511 52960 89940 52988
rect 88511 52957 88523 52960
rect 88465 52951 88523 52957
rect 89934 52948 89940 52960
rect 89992 52948 89998 53000
rect 4876 52794 7912 52816
rect 4876 52742 6690 52794
rect 6742 52742 6754 52794
rect 6806 52742 6818 52794
rect 6870 52742 6882 52794
rect 6934 52742 6946 52794
rect 6998 52742 7912 52794
rect 4876 52720 7912 52742
rect 86020 52794 88964 52816
rect 86020 52742 87834 52794
rect 87886 52742 87898 52794
rect 87950 52742 87962 52794
rect 88014 52742 88026 52794
rect 88078 52742 88090 52794
rect 88142 52742 88964 52794
rect 86020 52720 88964 52742
rect 5159 52549 5217 52555
rect 2902 52472 2908 52524
rect 2960 52512 2966 52524
rect 5159 52515 5171 52549
rect 5205 52515 5217 52549
rect 88325 52549 88383 52555
rect 88325 52546 88337 52549
rect 5159 52512 5217 52515
rect 2960 52509 5217 52512
rect 2960 52484 5202 52509
rect 2960 52472 2966 52484
rect 84322 52472 84328 52524
rect 84380 52512 84386 52524
rect 88020 52518 88337 52546
rect 88020 52512 88048 52518
rect 84380 52484 88048 52512
rect 88325 52515 88337 52518
rect 88371 52515 88383 52549
rect 88325 52509 88383 52515
rect 84380 52472 84386 52484
rect 5365 52379 5423 52385
rect 5365 52345 5377 52379
rect 5411 52376 5423 52379
rect 7134 52376 7140 52388
rect 5411 52348 7140 52376
rect 5411 52345 5423 52348
rect 5365 52339 5423 52345
rect 7134 52336 7140 52348
rect 7192 52336 7198 52388
rect 88554 52385 88560 52388
rect 88537 52379 88560 52385
rect 88537 52345 88549 52379
rect 88537 52339 88560 52345
rect 88554 52336 88560 52339
rect 88612 52336 88618 52388
rect 4876 52250 7912 52272
rect 4876 52198 5954 52250
rect 6006 52198 6018 52250
rect 6070 52198 6082 52250
rect 6134 52198 6146 52250
rect 6198 52198 6210 52250
rect 6262 52198 7912 52250
rect 4876 52176 7912 52198
rect 86020 52250 88964 52272
rect 86020 52198 87098 52250
rect 87150 52198 87162 52250
rect 87214 52198 87226 52250
rect 87278 52198 87290 52250
rect 87342 52198 87354 52250
rect 87406 52198 88964 52250
rect 86020 52176 88964 52198
rect 4876 51706 7912 51728
rect 4876 51654 6690 51706
rect 6742 51654 6754 51706
rect 6806 51654 6818 51706
rect 6870 51654 6882 51706
rect 6934 51654 6946 51706
rect 6998 51654 7912 51706
rect 4876 51632 7912 51654
rect 86020 51706 88964 51728
rect 86020 51654 87834 51706
rect 87886 51654 87898 51706
rect 87950 51654 87962 51706
rect 88014 51654 88026 51706
rect 88078 51654 88090 51706
rect 88142 51654 88964 51706
rect 86020 51632 88964 51654
rect 5159 51461 5217 51467
rect 2902 51384 2908 51436
rect 2960 51424 2966 51436
rect 5159 51427 5171 51461
rect 5205 51427 5217 51461
rect 5159 51424 5217 51427
rect 2960 51421 5217 51424
rect 2960 51396 5202 51421
rect 88370 51418 88376 51470
rect 88428 51418 88434 51470
rect 2960 51384 2966 51396
rect 5364 51359 5422 51365
rect 5364 51325 5376 51359
rect 5410 51356 5422 51359
rect 5662 51356 5668 51368
rect 5410 51328 5668 51356
rect 5410 51325 5422 51328
rect 5364 51319 5422 51325
rect 5662 51316 5668 51328
rect 5720 51316 5726 51368
rect 88554 51365 88560 51368
rect 88537 51359 88560 51365
rect 88537 51325 88549 51359
rect 88537 51319 88560 51325
rect 88554 51316 88560 51319
rect 88612 51316 88618 51368
rect 4876 51162 7912 51184
rect 4876 51110 5954 51162
rect 6006 51110 6018 51162
rect 6070 51110 6082 51162
rect 6134 51110 6146 51162
rect 6198 51110 6210 51162
rect 6262 51110 7912 51162
rect 4876 51088 7912 51110
rect 86020 51162 88964 51184
rect 86020 51110 87098 51162
rect 87150 51110 87162 51162
rect 87214 51110 87226 51162
rect 87278 51110 87290 51162
rect 87342 51110 87354 51162
rect 87406 51110 88964 51162
rect 86020 51088 88964 51110
rect 4876 50618 7912 50640
rect 4876 50566 6690 50618
rect 6742 50566 6754 50618
rect 6806 50566 6818 50618
rect 6870 50566 6882 50618
rect 6934 50566 6946 50618
rect 6998 50566 7912 50618
rect 4876 50544 7912 50566
rect 86020 50618 88964 50640
rect 86020 50566 87834 50618
rect 87886 50566 87898 50618
rect 87950 50566 87962 50618
rect 88014 50566 88026 50618
rect 88078 50566 88090 50618
rect 88142 50566 88964 50618
rect 86020 50544 88964 50566
rect 4876 50074 7912 50096
rect 4876 50022 5954 50074
rect 6006 50022 6018 50074
rect 6070 50022 6082 50074
rect 6134 50022 6146 50074
rect 6198 50022 6210 50074
rect 6262 50022 7912 50074
rect 4876 50000 7912 50022
rect 86020 50074 88964 50096
rect 86020 50022 87098 50074
rect 87150 50022 87162 50074
rect 87214 50022 87226 50074
rect 87278 50022 87290 50074
rect 87342 50022 87354 50074
rect 87406 50022 88964 50074
rect 86020 50000 88964 50022
rect 2902 49684 2908 49736
rect 2960 49724 2966 49736
rect 5205 49727 5263 49733
rect 5205 49724 5217 49727
rect 2960 49696 5217 49724
rect 2960 49684 2966 49696
rect 5205 49693 5217 49696
rect 5251 49693 5263 49727
rect 5205 49687 5263 49693
rect 88465 49727 88523 49733
rect 88465 49693 88477 49727
rect 88511 49724 88523 49727
rect 89934 49724 89940 49736
rect 88511 49696 89940 49724
rect 88511 49693 88523 49696
rect 88465 49687 88523 49693
rect 89934 49684 89940 49696
rect 89992 49684 89998 49736
rect 4876 49530 7912 49552
rect 4876 49478 6690 49530
rect 6742 49478 6754 49530
rect 6806 49478 6818 49530
rect 6870 49478 6882 49530
rect 6934 49478 6946 49530
rect 6998 49478 7912 49530
rect 4876 49456 7912 49478
rect 86020 49530 88964 49552
rect 86020 49478 87834 49530
rect 87886 49478 87898 49530
rect 87950 49478 87962 49530
rect 88014 49478 88026 49530
rect 88078 49478 88090 49530
rect 88142 49478 88964 49530
rect 86020 49456 88964 49478
rect 4876 48986 7912 49008
rect 4876 48934 5954 48986
rect 6006 48934 6018 48986
rect 6070 48934 6082 48986
rect 6134 48934 6146 48986
rect 6198 48934 6210 48986
rect 6262 48934 7912 48986
rect 4876 48912 7912 48934
rect 86020 48986 88964 49008
rect 86020 48934 87098 48986
rect 87150 48934 87162 48986
rect 87214 48934 87226 48986
rect 87278 48934 87290 48986
rect 87342 48934 87354 48986
rect 87406 48934 88964 48986
rect 86020 48912 88964 48934
rect 88465 48639 88523 48645
rect 88465 48605 88477 48639
rect 88511 48636 88523 48639
rect 89934 48636 89940 48648
rect 88511 48608 89940 48636
rect 88511 48605 88523 48608
rect 88465 48599 88523 48605
rect 89934 48596 89940 48608
rect 89992 48596 89998 48648
rect 4876 48442 7912 48464
rect 4876 48390 6690 48442
rect 6742 48390 6754 48442
rect 6806 48390 6818 48442
rect 6870 48390 6882 48442
rect 6934 48390 6946 48442
rect 6998 48390 7912 48442
rect 4876 48368 7912 48390
rect 86020 48442 88964 48464
rect 86020 48390 87834 48442
rect 87886 48390 87898 48442
rect 87950 48390 87962 48442
rect 88014 48390 88026 48442
rect 88078 48390 88090 48442
rect 88142 48390 88964 48442
rect 86020 48368 88964 48390
rect 88325 48197 88383 48203
rect 88325 48194 88337 48197
rect 88204 48166 88337 48194
rect 88204 48033 88232 48166
rect 88325 48163 88337 48166
rect 88371 48163 88383 48197
rect 88325 48157 88383 48163
rect 88554 48033 88560 48036
rect 88189 48027 88247 48033
rect 88189 48024 88201 48027
rect 85766 47996 88201 48024
rect 4876 47898 7912 47920
rect 4876 47846 5954 47898
rect 6006 47846 6018 47898
rect 6070 47846 6082 47898
rect 6134 47846 6146 47898
rect 6198 47846 6210 47898
rect 6262 47846 7912 47898
rect 4876 47824 7912 47846
rect 4876 47354 7912 47376
rect 4876 47302 6690 47354
rect 6742 47302 6754 47354
rect 6806 47302 6818 47354
rect 6870 47302 6882 47354
rect 6934 47302 6946 47354
rect 6998 47302 7912 47354
rect 12222 47304 12228 47356
rect 12280 47344 12286 47356
rect 49224 47344 49230 47356
rect 12280 47316 49230 47344
rect 12280 47304 12286 47316
rect 49224 47304 49230 47316
rect 49282 47304 49288 47356
rect 51432 47304 51438 47356
rect 51490 47344 51496 47356
rect 84414 47344 84420 47356
rect 51490 47316 84420 47344
rect 51490 47304 51496 47316
rect 84414 47304 84420 47316
rect 84472 47304 84478 47356
rect 4876 47280 7912 47302
rect 8146 47236 8152 47288
rect 8204 47276 8210 47288
rect 14430 47276 14436 47288
rect 8204 47248 14436 47276
rect 8204 47236 8210 47248
rect 14430 47236 14436 47248
rect 14488 47236 14494 47288
rect 7870 47168 7876 47220
rect 7928 47208 7934 47220
rect 12194 47208 12200 47220
rect 7928 47180 12200 47208
rect 7928 47168 7934 47180
rect 12194 47168 12200 47180
rect 12252 47168 12258 47220
rect 48166 47168 48172 47220
rect 48224 47208 48230 47220
rect 85766 47208 85794 47996
rect 88189 47993 88201 47996
rect 88235 47993 88247 48027
rect 88189 47987 88247 47993
rect 88537 48027 88560 48033
rect 88537 47993 88549 48027
rect 88537 47987 88560 47993
rect 88554 47984 88560 47987
rect 88612 47984 88618 48036
rect 86020 47898 88964 47920
rect 86020 47846 87098 47898
rect 87150 47846 87162 47898
rect 87214 47846 87226 47898
rect 87278 47846 87290 47898
rect 87342 47846 87354 47898
rect 87406 47846 88964 47898
rect 86020 47824 88964 47846
rect 86020 47354 88964 47376
rect 86020 47302 87834 47354
rect 87886 47302 87898 47354
rect 87950 47302 87962 47354
rect 88014 47302 88026 47354
rect 88078 47302 88090 47354
rect 88142 47302 88964 47354
rect 86020 47280 88964 47302
rect 48224 47180 85794 47208
rect 48224 47168 48230 47180
rect 2902 47100 2908 47152
rect 2960 47140 2966 47152
rect 5225 47143 5283 47149
rect 5225 47140 5237 47143
rect 2960 47112 5237 47140
rect 2960 47100 2966 47112
rect 5225 47109 5237 47112
rect 5271 47109 5283 47143
rect 5225 47103 5283 47109
rect 7042 47100 7048 47152
rect 7100 47140 7106 47152
rect 10998 47140 11004 47152
rect 7100 47112 11004 47140
rect 7100 47100 7106 47112
rect 10998 47100 11004 47112
rect 11056 47100 11062 47152
rect 5527 46939 5585 46945
rect 5527 46905 5539 46939
rect 5573 46936 5585 46939
rect 14126 46936 14132 46948
rect 5573 46908 14132 46936
rect 5573 46905 5585 46908
rect 5527 46899 5585 46905
rect 14126 46896 14132 46908
rect 14184 46896 14190 46948
rect 88554 46896 88560 46948
rect 88612 46896 88618 46948
rect 4876 46810 7912 46832
rect 13574 46828 13580 46880
rect 13632 46868 13638 46880
rect 50190 46868 50196 46880
rect 13632 46840 50196 46868
rect 13632 46828 13638 46840
rect 50190 46828 50196 46840
rect 50248 46828 50254 46880
rect 4876 46758 5954 46810
rect 6006 46758 6018 46810
rect 6070 46758 6082 46810
rect 6134 46758 6146 46810
rect 6198 46758 6210 46810
rect 6262 46758 7912 46810
rect 12470 46760 12476 46812
rect 12528 46800 12534 46812
rect 49086 46800 49092 46812
rect 12528 46772 49092 46800
rect 12528 46760 12534 46772
rect 49086 46760 49092 46772
rect 49144 46760 49150 46812
rect 50650 46760 50656 46812
rect 50708 46800 50714 46812
rect 84046 46800 84052 46812
rect 50708 46772 84052 46800
rect 50708 46760 50714 46772
rect 84046 46760 84052 46772
rect 84104 46760 84110 46812
rect 86020 46810 88964 46832
rect 4876 46736 7912 46758
rect 86020 46758 87098 46810
rect 87150 46758 87162 46810
rect 87214 46758 87226 46810
rect 87278 46758 87290 46810
rect 87342 46758 87354 46810
rect 87406 46758 88964 46810
rect 10998 46692 11004 46744
rect 11056 46732 11062 46744
rect 47798 46732 47804 46744
rect 11056 46704 47804 46732
rect 11056 46692 11062 46704
rect 47798 46692 47804 46704
rect 47856 46692 47862 46744
rect 49546 46692 49552 46744
rect 49604 46732 49610 46744
rect 83678 46732 83684 46744
rect 49604 46704 83684 46732
rect 49604 46692 49610 46704
rect 83678 46692 83684 46704
rect 83736 46692 83742 46744
rect 86020 46736 88964 46758
rect 4876 46266 7912 46288
rect 4876 46214 6690 46266
rect 6742 46214 6754 46266
rect 6806 46214 6818 46266
rect 6870 46214 6882 46266
rect 6934 46214 6946 46266
rect 6998 46214 7912 46266
rect 4876 46192 7912 46214
rect 86020 46266 88964 46288
rect 86020 46214 87834 46266
rect 87886 46214 87898 46266
rect 87950 46214 87962 46266
rect 88014 46214 88026 46266
rect 88078 46214 88090 46266
rect 88142 46214 88964 46266
rect 86020 46192 88964 46214
rect 2902 45808 2908 45860
rect 2960 45848 2966 45860
rect 5205 45851 5263 45857
rect 5205 45848 5217 45851
rect 2960 45820 5217 45848
rect 2960 45808 2966 45820
rect 5205 45817 5217 45820
rect 5251 45817 5263 45851
rect 5205 45811 5263 45817
rect 4876 45722 7912 45744
rect 4876 45670 5954 45722
rect 6006 45670 6018 45722
rect 6070 45670 6082 45722
rect 6134 45670 6146 45722
rect 6198 45670 6210 45722
rect 6262 45670 7912 45722
rect 4876 45648 7912 45670
rect 86020 45722 88964 45744
rect 86020 45670 87098 45722
rect 87150 45670 87162 45722
rect 87214 45670 87226 45722
rect 87278 45670 87290 45722
rect 87342 45670 87354 45722
rect 87406 45670 88964 45722
rect 86020 45648 88964 45670
rect 4876 45178 7912 45200
rect 4876 45126 6690 45178
rect 6742 45126 6754 45178
rect 6806 45126 6818 45178
rect 6870 45126 6882 45178
rect 6934 45126 6946 45178
rect 6998 45126 7912 45178
rect 4876 45104 7912 45126
rect 86020 45178 88964 45200
rect 86020 45126 87834 45178
rect 87886 45126 87898 45178
rect 87950 45126 87962 45178
rect 88014 45126 88026 45178
rect 88078 45126 88090 45178
rect 88142 45126 88964 45178
rect 86020 45104 88964 45126
rect 2534 44720 2540 44772
rect 2592 44760 2598 44772
rect 5205 44763 5263 44769
rect 5205 44760 5217 44763
rect 2592 44732 5217 44760
rect 2592 44720 2598 44732
rect 5205 44729 5217 44732
rect 5251 44729 5263 44763
rect 5205 44723 5263 44729
rect 4876 44634 7912 44656
rect 4876 44582 5954 44634
rect 6006 44582 6018 44634
rect 6070 44582 6082 44634
rect 6134 44582 6146 44634
rect 6198 44582 6210 44634
rect 6262 44582 7912 44634
rect 4876 44560 7912 44582
rect 86020 44634 88964 44656
rect 86020 44582 87098 44634
rect 87150 44582 87162 44634
rect 87214 44582 87226 44634
rect 87278 44582 87290 44634
rect 87342 44582 87354 44634
rect 87406 44582 88964 44634
rect 86020 44560 88964 44582
rect 5202 44380 5208 44432
rect 5260 44380 5266 44432
rect 4876 44090 7912 44112
rect 4876 44038 6690 44090
rect 6742 44038 6754 44090
rect 6806 44038 6818 44090
rect 6870 44038 6882 44090
rect 6934 44038 6946 44090
rect 6998 44038 7912 44090
rect 4876 44016 7912 44038
rect 86020 44090 88964 44112
rect 86020 44038 87834 44090
rect 87886 44038 87898 44090
rect 87950 44038 87962 44090
rect 88014 44038 88026 44090
rect 88078 44038 88090 44090
rect 88142 44038 88964 44090
rect 86020 44016 88964 44038
rect 4876 43546 7912 43568
rect 4876 43494 5954 43546
rect 6006 43494 6018 43546
rect 6070 43494 6082 43546
rect 6134 43494 6146 43546
rect 6198 43494 6210 43546
rect 6262 43494 7912 43546
rect 4876 43472 7912 43494
rect 86020 43546 88964 43568
rect 86020 43494 87098 43546
rect 87150 43494 87162 43546
rect 87214 43494 87226 43546
rect 87278 43494 87290 43546
rect 87342 43494 87354 43546
rect 87406 43494 88964 43546
rect 86020 43472 88964 43494
rect 88511 43267 88569 43273
rect 5457 43233 5515 43239
rect 5457 43199 5469 43233
rect 5503 43230 5515 43233
rect 88511 43233 88523 43267
rect 88557 43264 88569 43267
rect 89934 43264 89940 43276
rect 88557 43236 89940 43264
rect 88557 43233 88569 43236
rect 5503 43202 5800 43230
rect 88511 43227 88569 43233
rect 89934 43224 89940 43236
rect 89992 43224 89998 43276
rect 5503 43199 5515 43202
rect 5457 43193 5515 43199
rect 5772 43196 5800 43202
rect 7134 43196 7140 43208
rect 5772 43168 7140 43196
rect 7134 43156 7140 43168
rect 7192 43156 7198 43208
rect 2902 43088 2908 43140
rect 2960 43128 2966 43140
rect 5251 43131 5309 43137
rect 5251 43128 5263 43131
rect 2960 43100 5263 43128
rect 2960 43088 2966 43100
rect 5251 43097 5263 43100
rect 5297 43097 5309 43131
rect 5251 43091 5309 43097
rect 84322 43088 84328 43140
rect 84380 43128 84386 43140
rect 88281 43131 88339 43137
rect 88281 43128 88293 43131
rect 84380 43100 88293 43128
rect 84380 43088 84386 43100
rect 88281 43097 88293 43100
rect 88327 43097 88339 43131
rect 88281 43091 88339 43097
rect 4876 43002 7912 43024
rect 4876 42950 6690 43002
rect 6742 42950 6754 43002
rect 6806 42950 6818 43002
rect 6870 42950 6882 43002
rect 6934 42950 6946 43002
rect 6998 42950 7912 43002
rect 4876 42928 7912 42950
rect 86020 43002 88964 43024
rect 86020 42950 87834 43002
rect 87886 42950 87898 43002
rect 87950 42950 87962 43002
rect 88014 42950 88026 43002
rect 88078 42950 88090 43002
rect 88142 42950 88964 43002
rect 86020 42928 88964 42950
rect 2902 42544 2908 42596
rect 2960 42584 2966 42596
rect 5205 42587 5263 42593
rect 5205 42584 5217 42587
rect 2960 42556 5217 42584
rect 2960 42544 2966 42556
rect 5205 42553 5217 42556
rect 5251 42553 5263 42587
rect 5205 42547 5263 42553
rect 4876 42458 7912 42480
rect 4876 42406 5954 42458
rect 6006 42406 6018 42458
rect 6070 42406 6082 42458
rect 6134 42406 6146 42458
rect 6198 42406 6210 42458
rect 6262 42406 7912 42458
rect 4876 42384 7912 42406
rect 86020 42458 88964 42480
rect 86020 42406 87098 42458
rect 87150 42406 87162 42458
rect 87214 42406 87226 42458
rect 87278 42406 87290 42458
rect 87342 42406 87354 42458
rect 87406 42406 88964 42458
rect 86020 42384 88964 42406
rect 88554 42151 88560 42154
rect 5457 42145 5515 42151
rect 5457 42111 5469 42145
rect 5503 42142 5515 42145
rect 88533 42145 88560 42151
rect 5503 42114 5800 42142
rect 5503 42111 5515 42114
rect 5457 42105 5515 42111
rect 5772 42108 5800 42114
rect 7134 42108 7140 42120
rect 5772 42080 7140 42108
rect 7134 42068 7140 42080
rect 7192 42068 7198 42120
rect 88533 42111 88545 42145
rect 88533 42105 88560 42111
rect 88554 42102 88560 42105
rect 88612 42102 88618 42154
rect 2902 42000 2908 42052
rect 2960 42040 2966 42052
rect 5251 42043 5309 42049
rect 5251 42040 5263 42043
rect 2960 42012 5263 42040
rect 2960 42000 2966 42012
rect 5251 42009 5263 42012
rect 5297 42009 5309 42043
rect 5251 42003 5309 42009
rect 84322 42000 84328 42052
rect 84380 42040 84386 42052
rect 88327 42043 88385 42049
rect 88327 42040 88339 42043
rect 84380 42012 88339 42040
rect 84380 42000 84386 42012
rect 88327 42009 88339 42012
rect 88373 42009 88385 42043
rect 88327 42003 88385 42009
rect 4876 41914 7912 41936
rect 4876 41862 6690 41914
rect 6742 41862 6754 41914
rect 6806 41862 6818 41914
rect 6870 41862 6882 41914
rect 6934 41862 6946 41914
rect 6998 41862 7912 41914
rect 4876 41840 7912 41862
rect 86020 41914 88964 41936
rect 86020 41862 87834 41914
rect 87886 41862 87898 41914
rect 87950 41862 87962 41914
rect 88014 41862 88026 41914
rect 88078 41862 88090 41914
rect 88142 41862 88964 41914
rect 86020 41840 88964 41862
rect 4374 41728 4380 41780
rect 4432 41768 4438 41780
rect 5251 41771 5309 41777
rect 5251 41768 5263 41771
rect 4432 41740 5263 41768
rect 4432 41728 4438 41740
rect 5251 41737 5263 41740
rect 5297 41737 5309 41771
rect 5251 41731 5309 41737
rect 87450 41728 87456 41780
rect 87508 41768 87514 41780
rect 88419 41771 88477 41777
rect 88419 41768 88431 41771
rect 87508 41740 88431 41768
rect 87508 41728 87514 41740
rect 88419 41737 88431 41740
rect 88465 41737 88477 41771
rect 88419 41731 88477 41737
rect 89934 41700 89940 41712
rect 5457 41669 5515 41675
rect 5457 41635 5469 41669
rect 5503 41666 5515 41669
rect 5662 41666 5668 41678
rect 5503 41638 5668 41666
rect 5503 41635 5515 41638
rect 5457 41629 5515 41635
rect 5662 41626 5668 41638
rect 5720 41626 5726 41678
rect 88625 41669 88683 41675
rect 88625 41635 88637 41669
rect 88671 41666 88683 41669
rect 88940 41672 89940 41700
rect 88940 41666 88968 41672
rect 88671 41638 88968 41666
rect 89934 41660 89940 41672
rect 89992 41660 89998 41712
rect 88671 41635 88683 41638
rect 88625 41629 88683 41635
rect 4876 41370 7912 41392
rect 4876 41318 5954 41370
rect 6006 41318 6018 41370
rect 6070 41318 6082 41370
rect 6134 41318 6146 41370
rect 6198 41318 6210 41370
rect 6262 41318 7912 41370
rect 4876 41296 7912 41318
rect 86020 41370 88964 41392
rect 86020 41318 87098 41370
rect 87150 41318 87162 41370
rect 87214 41318 87226 41370
rect 87278 41318 87290 41370
rect 87342 41318 87354 41370
rect 87406 41318 88964 41370
rect 86020 41296 88964 41318
rect 4876 40826 7912 40848
rect 4876 40774 6690 40826
rect 6742 40774 6754 40826
rect 6806 40774 6818 40826
rect 6870 40774 6882 40826
rect 6934 40774 6946 40826
rect 6998 40774 7912 40826
rect 4876 40752 7912 40774
rect 86020 40826 88964 40848
rect 86020 40774 87834 40826
rect 87886 40774 87898 40826
rect 87950 40774 87962 40826
rect 88014 40774 88026 40826
rect 88078 40774 88090 40826
rect 88142 40774 88964 40826
rect 86020 40752 88964 40774
rect 4876 40282 7912 40304
rect 4876 40230 5954 40282
rect 6006 40230 6018 40282
rect 6070 40230 6082 40282
rect 6134 40230 6146 40282
rect 6198 40230 6210 40282
rect 6262 40230 7912 40282
rect 4876 40208 7912 40230
rect 86020 40282 88964 40304
rect 86020 40230 87098 40282
rect 87150 40230 87162 40282
rect 87214 40230 87226 40282
rect 87278 40230 87290 40282
rect 87342 40230 87354 40282
rect 87406 40230 88964 40282
rect 86020 40208 88964 40230
rect 5457 39969 5515 39975
rect 5457 39935 5469 39969
rect 5503 39966 5515 39969
rect 5503 39938 5800 39966
rect 5503 39935 5515 39938
rect 5457 39929 5515 39935
rect 5772 39932 5800 39938
rect 7134 39932 7140 39944
rect 5772 39904 7140 39932
rect 7134 39892 7140 39904
rect 7192 39892 7198 39944
rect 84322 39892 84328 39944
rect 84380 39932 84386 39944
rect 88097 39935 88155 39941
rect 88097 39932 88109 39935
rect 84380 39904 88109 39932
rect 84380 39892 84386 39904
rect 88097 39901 88109 39904
rect 88143 39901 88155 39935
rect 88097 39895 88155 39901
rect 88465 39935 88523 39941
rect 88465 39901 88477 39935
rect 88511 39932 88523 39935
rect 89934 39932 89940 39944
rect 88511 39904 89940 39932
rect 88511 39901 88523 39904
rect 88465 39895 88523 39901
rect 89934 39892 89940 39904
rect 89992 39892 89998 39944
rect 2902 39824 2908 39876
rect 2960 39864 2966 39876
rect 5251 39867 5309 39873
rect 5251 39864 5263 39867
rect 2960 39836 5263 39864
rect 2960 39824 2966 39836
rect 5251 39833 5263 39836
rect 5297 39833 5309 39867
rect 5251 39827 5309 39833
rect 4876 39738 7912 39760
rect 4876 39686 6690 39738
rect 6742 39686 6754 39738
rect 6806 39686 6818 39738
rect 6870 39686 6882 39738
rect 6934 39686 6946 39738
rect 6998 39686 7912 39738
rect 4876 39664 7912 39686
rect 86020 39738 88964 39760
rect 86020 39686 87834 39738
rect 87886 39686 87898 39738
rect 87950 39686 87962 39738
rect 88014 39686 88026 39738
rect 88078 39686 88090 39738
rect 88142 39686 88964 39738
rect 86020 39664 88964 39686
rect 4876 39194 7912 39216
rect 4876 39142 5954 39194
rect 6006 39142 6018 39194
rect 6070 39142 6082 39194
rect 6134 39142 6146 39194
rect 6198 39142 6210 39194
rect 6262 39142 7912 39194
rect 4876 39120 7912 39142
rect 86020 39194 88964 39216
rect 86020 39142 87098 39194
rect 87150 39142 87162 39194
rect 87214 39142 87226 39194
rect 87278 39142 87290 39194
rect 87342 39142 87354 39194
rect 87406 39142 88964 39194
rect 86020 39120 88964 39142
rect 4374 38940 4380 38992
rect 4432 38980 4438 38992
rect 5251 38983 5309 38989
rect 5251 38980 5263 38983
rect 4432 38952 5263 38980
rect 4432 38940 4438 38952
rect 5251 38949 5263 38952
rect 5297 38949 5309 38983
rect 5251 38943 5309 38949
rect 87174 38940 87180 38992
rect 87232 38980 87238 38992
rect 88327 38983 88385 38989
rect 88327 38980 88339 38983
rect 87232 38952 88339 38980
rect 87232 38940 87238 38952
rect 88327 38949 88339 38952
rect 88373 38949 88385 38983
rect 88327 38943 88385 38949
rect 5457 38881 5515 38887
rect 5457 38847 5469 38881
rect 5503 38878 5515 38881
rect 88533 38881 88591 38887
rect 5503 38847 5524 38878
rect 5457 38844 5524 38847
rect 7410 38844 7416 38856
rect 5457 38841 7416 38844
rect 5496 38816 7416 38841
rect 7410 38804 7416 38816
rect 7468 38804 7474 38856
rect 88533 38847 88545 38881
rect 88579 38878 88591 38881
rect 88579 38847 88600 38878
rect 88533 38844 88600 38847
rect 89290 38844 89296 38856
rect 88533 38841 89296 38844
rect 88572 38816 89296 38841
rect 89290 38804 89296 38816
rect 89348 38804 89354 38856
rect 4876 38650 7912 38672
rect 4876 38598 6690 38650
rect 6742 38598 6754 38650
rect 6806 38598 6818 38650
rect 6870 38598 6882 38650
rect 6934 38598 6946 38650
rect 6998 38598 7912 38650
rect 4876 38576 7912 38598
rect 86020 38650 88964 38672
rect 86020 38598 87834 38650
rect 87886 38598 87898 38650
rect 87950 38598 87962 38650
rect 88014 38598 88026 38650
rect 88078 38598 88090 38650
rect 88142 38598 88964 38650
rect 86020 38576 88964 38598
rect 4876 38106 7912 38128
rect 4876 38054 5954 38106
rect 6006 38054 6018 38106
rect 6070 38054 6082 38106
rect 6134 38054 6146 38106
rect 6198 38054 6210 38106
rect 6262 38054 7912 38106
rect 4876 38032 7912 38054
rect 86020 38106 88964 38128
rect 86020 38054 87098 38106
rect 87150 38054 87162 38106
rect 87214 38054 87226 38106
rect 87278 38054 87290 38106
rect 87342 38054 87354 38106
rect 87406 38054 88964 38106
rect 86020 38032 88964 38054
rect 5457 37793 5515 37799
rect 5457 37759 5469 37793
rect 5503 37790 5515 37793
rect 5503 37762 5800 37790
rect 5503 37759 5515 37762
rect 5457 37753 5515 37759
rect 5772 37756 5800 37762
rect 7134 37756 7140 37768
rect 5772 37728 7140 37756
rect 7134 37716 7140 37728
rect 7192 37716 7198 37768
rect 84322 37716 84328 37768
rect 84380 37756 84386 37768
rect 88235 37759 88293 37765
rect 88235 37756 88247 37759
rect 84380 37728 88247 37756
rect 84380 37716 84386 37728
rect 88235 37725 88247 37728
rect 88281 37725 88293 37759
rect 88235 37719 88293 37725
rect 88465 37759 88523 37765
rect 88465 37725 88477 37759
rect 88511 37756 88523 37759
rect 89934 37756 89940 37768
rect 88511 37728 89940 37756
rect 88511 37725 88523 37728
rect 88465 37719 88523 37725
rect 89934 37716 89940 37728
rect 89992 37716 89998 37768
rect 2902 37648 2908 37700
rect 2960 37688 2966 37700
rect 5251 37691 5309 37697
rect 5251 37688 5263 37691
rect 2960 37660 5263 37688
rect 2960 37648 2966 37660
rect 5251 37657 5263 37660
rect 5297 37657 5309 37691
rect 5251 37651 5309 37657
rect 4876 37562 7912 37584
rect 4876 37510 6690 37562
rect 6742 37510 6754 37562
rect 6806 37510 6818 37562
rect 6870 37510 6882 37562
rect 6934 37510 6946 37562
rect 6998 37510 7912 37562
rect 4876 37488 7912 37510
rect 86020 37562 88964 37584
rect 86020 37510 87834 37562
rect 87886 37510 87898 37562
rect 87950 37510 87962 37562
rect 88014 37510 88026 37562
rect 88078 37510 88090 37562
rect 88142 37510 88964 37562
rect 86020 37488 88964 37510
rect 4876 37018 7912 37040
rect 4876 36966 5954 37018
rect 6006 36966 6018 37018
rect 6070 36966 6082 37018
rect 6134 36966 6146 37018
rect 6198 36966 6210 37018
rect 6262 36966 7912 37018
rect 4876 36944 7912 36966
rect 86020 37018 88964 37040
rect 86020 36966 87098 37018
rect 87150 36966 87162 37018
rect 87214 36966 87226 37018
rect 87278 36966 87290 37018
rect 87342 36966 87354 37018
rect 87406 36966 88964 37018
rect 86020 36944 88964 36966
rect 5457 36705 5515 36711
rect 5457 36671 5469 36705
rect 5503 36671 5515 36705
rect 5457 36668 5515 36671
rect 7134 36668 7140 36680
rect 5457 36665 7140 36668
rect 5472 36640 7140 36665
rect 7134 36628 7140 36640
rect 7192 36628 7198 36680
rect 84322 36628 84328 36680
rect 84380 36668 84386 36680
rect 88235 36671 88293 36677
rect 88235 36668 88247 36671
rect 84380 36640 88247 36668
rect 84380 36628 84386 36640
rect 88235 36637 88247 36640
rect 88281 36637 88293 36671
rect 88235 36631 88293 36637
rect 88465 36671 88523 36677
rect 88465 36637 88477 36671
rect 88511 36668 88523 36671
rect 89934 36668 89940 36680
rect 88511 36640 89940 36668
rect 88511 36637 88523 36640
rect 88465 36631 88523 36637
rect 89934 36628 89940 36640
rect 89992 36628 89998 36680
rect 2902 36560 2908 36612
rect 2960 36600 2966 36612
rect 5251 36603 5309 36609
rect 5251 36600 5263 36603
rect 2960 36572 5263 36600
rect 2960 36560 2966 36572
rect 5251 36569 5263 36572
rect 5297 36569 5309 36603
rect 5251 36563 5309 36569
rect 4876 36474 7912 36496
rect 4876 36422 6690 36474
rect 6742 36422 6754 36474
rect 6806 36422 6818 36474
rect 6870 36422 6882 36474
rect 6934 36422 6946 36474
rect 6998 36422 7912 36474
rect 4876 36400 7912 36422
rect 86020 36474 88964 36496
rect 86020 36422 87834 36474
rect 87886 36422 87898 36474
rect 87950 36422 87962 36474
rect 88014 36422 88026 36474
rect 88078 36422 88090 36474
rect 88142 36422 88964 36474
rect 86020 36400 88964 36422
rect 5457 36229 5515 36235
rect 5457 36195 5469 36229
rect 5503 36226 5515 36229
rect 5662 36226 5668 36238
rect 5503 36198 5668 36226
rect 5503 36195 5515 36198
rect 5457 36189 5515 36195
rect 5662 36186 5668 36198
rect 5720 36186 5726 36238
rect 88603 36211 88661 36217
rect 88603 36177 88615 36211
rect 88649 36208 88661 36211
rect 88649 36192 88876 36208
rect 90118 36192 90124 36204
rect 88649 36180 90124 36192
rect 88649 36177 88661 36180
rect 88603 36171 88661 36177
rect 88848 36164 90124 36180
rect 90118 36152 90124 36164
rect 90176 36152 90182 36204
rect 4374 36084 4380 36136
rect 4432 36124 4438 36136
rect 5251 36127 5309 36133
rect 5251 36124 5263 36127
rect 4432 36096 5263 36124
rect 4432 36084 4438 36096
rect 5251 36093 5263 36096
rect 5297 36093 5309 36127
rect 5251 36087 5309 36093
rect 87450 36084 87456 36136
rect 87508 36124 87514 36136
rect 88419 36127 88477 36133
rect 88419 36124 88431 36127
rect 87508 36096 88431 36124
rect 87508 36084 87514 36096
rect 88419 36093 88431 36096
rect 88465 36093 88477 36127
rect 88419 36087 88477 36093
rect 4876 35930 7912 35952
rect 4876 35878 5954 35930
rect 6006 35878 6018 35930
rect 6070 35878 6082 35930
rect 6134 35878 6146 35930
rect 6198 35878 6210 35930
rect 6262 35878 7912 35930
rect 4876 35856 7912 35878
rect 86020 35930 88964 35952
rect 86020 35878 87098 35930
rect 87150 35878 87162 35930
rect 87214 35878 87226 35930
rect 87278 35878 87290 35930
rect 87342 35878 87354 35930
rect 87406 35878 88964 35930
rect 86020 35856 88964 35878
rect 4876 35386 7912 35408
rect 4876 35334 6690 35386
rect 6742 35334 6754 35386
rect 6806 35334 6818 35386
rect 6870 35334 6882 35386
rect 6934 35334 6946 35386
rect 6998 35334 7912 35386
rect 4876 35312 7912 35334
rect 86020 35386 88964 35408
rect 86020 35334 87834 35386
rect 87886 35334 87898 35386
rect 87950 35334 87962 35386
rect 88014 35334 88026 35386
rect 88078 35334 88090 35386
rect 88142 35334 88964 35386
rect 86020 35312 88964 35334
rect 4876 34842 7912 34864
rect 4876 34790 5954 34842
rect 6006 34790 6018 34842
rect 6070 34790 6082 34842
rect 6134 34790 6146 34842
rect 6198 34790 6210 34842
rect 6262 34790 7912 34842
rect 4876 34768 7912 34790
rect 86020 34842 88964 34864
rect 86020 34790 87098 34842
rect 87150 34790 87162 34842
rect 87214 34790 87226 34842
rect 87278 34790 87290 34842
rect 87342 34790 87354 34842
rect 87406 34790 88964 34842
rect 86020 34768 88964 34790
rect 5457 34529 5515 34535
rect 88554 34529 88560 34532
rect 5457 34495 5469 34529
rect 5503 34495 5515 34529
rect 88529 34523 88560 34529
rect 5457 34492 5515 34495
rect 7134 34492 7140 34504
rect 5457 34489 7140 34492
rect 5472 34464 7140 34489
rect 7134 34452 7140 34464
rect 7192 34452 7198 34504
rect 88529 34489 88541 34523
rect 88529 34483 88560 34489
rect 88554 34480 88560 34483
rect 88612 34480 88618 34532
rect 2902 34384 2908 34436
rect 2960 34424 2966 34436
rect 5251 34427 5309 34433
rect 5251 34424 5263 34427
rect 2960 34396 5263 34424
rect 2960 34384 2966 34396
rect 5251 34393 5263 34396
rect 5297 34393 5309 34427
rect 5251 34387 5309 34393
rect 84322 34384 84328 34436
rect 84380 34424 84386 34436
rect 88327 34427 88385 34433
rect 88327 34424 88339 34427
rect 84380 34396 88339 34424
rect 84380 34384 84386 34396
rect 88327 34393 88339 34396
rect 88373 34393 88385 34427
rect 88327 34387 88385 34393
rect 4876 34298 7912 34320
rect 4876 34246 6690 34298
rect 6742 34246 6754 34298
rect 6806 34246 6818 34298
rect 6870 34246 6882 34298
rect 6934 34246 6946 34298
rect 6998 34246 7912 34298
rect 4876 34224 7912 34246
rect 86020 34298 88964 34320
rect 86020 34246 87834 34298
rect 87886 34246 87898 34298
rect 87950 34246 87962 34298
rect 88014 34246 88026 34298
rect 88078 34246 88090 34298
rect 88142 34246 88964 34298
rect 86020 34224 88964 34246
rect 2902 33840 2908 33892
rect 2960 33880 2966 33892
rect 5205 33883 5263 33889
rect 5205 33880 5217 33883
rect 2960 33852 5217 33880
rect 2960 33840 2966 33852
rect 5205 33849 5217 33852
rect 5251 33849 5263 33883
rect 5205 33843 5263 33849
rect 4876 33754 7912 33776
rect 4876 33702 5954 33754
rect 6006 33702 6018 33754
rect 6070 33702 6082 33754
rect 6134 33702 6146 33754
rect 6198 33702 6210 33754
rect 6262 33702 7912 33754
rect 4876 33680 7912 33702
rect 86020 33754 88964 33776
rect 86020 33702 87098 33754
rect 87150 33702 87162 33754
rect 87214 33702 87226 33754
rect 87278 33702 87290 33754
rect 87342 33702 87354 33754
rect 87406 33702 88964 33754
rect 86020 33680 88964 33702
rect 4374 33500 4380 33552
rect 4432 33540 4438 33552
rect 5251 33543 5309 33549
rect 5251 33540 5263 33543
rect 4432 33512 5263 33540
rect 4432 33500 4438 33512
rect 5251 33509 5263 33512
rect 5297 33509 5309 33543
rect 5251 33503 5309 33509
rect 5457 33441 5515 33447
rect 5457 33407 5469 33441
rect 5503 33438 5515 33441
rect 5662 33438 5668 33450
rect 5503 33410 5668 33438
rect 5503 33407 5515 33410
rect 5457 33401 5515 33407
rect 5662 33398 5668 33410
rect 5720 33398 5726 33450
rect 87174 33364 87180 33416
rect 87232 33404 87238 33416
rect 88235 33407 88293 33413
rect 88235 33404 88247 33407
rect 87232 33376 88247 33404
rect 87232 33364 87238 33376
rect 88235 33373 88247 33376
rect 88281 33373 88293 33407
rect 88235 33367 88293 33373
rect 88465 33407 88523 33413
rect 88465 33373 88477 33407
rect 88511 33404 88523 33407
rect 89934 33404 89940 33416
rect 88511 33376 89940 33404
rect 88511 33373 88523 33376
rect 88465 33367 88523 33373
rect 89934 33364 89940 33376
rect 89992 33364 89998 33416
rect 4876 33210 7912 33232
rect 4876 33158 6690 33210
rect 6742 33158 6754 33210
rect 6806 33158 6818 33210
rect 6870 33158 6882 33210
rect 6934 33158 6946 33210
rect 6998 33158 7912 33210
rect 4876 33136 7912 33158
rect 86020 33210 88964 33232
rect 86020 33158 87834 33210
rect 87886 33158 87898 33210
rect 87950 33158 87962 33210
rect 88014 33158 88026 33210
rect 88078 33158 88090 33210
rect 88142 33158 88964 33210
rect 86020 33136 88964 33158
rect 4876 32666 7912 32688
rect 4876 32614 5954 32666
rect 6006 32614 6018 32666
rect 6070 32614 6082 32666
rect 6134 32614 6146 32666
rect 6198 32614 6210 32666
rect 6262 32614 7912 32666
rect 4876 32592 7912 32614
rect 86020 32666 88964 32688
rect 86020 32614 87098 32666
rect 87150 32614 87162 32666
rect 87214 32614 87226 32666
rect 87278 32614 87290 32666
rect 87342 32614 87354 32666
rect 87406 32614 88964 32666
rect 86020 32592 88964 32614
rect 5457 32353 5515 32359
rect 5457 32319 5469 32353
rect 5503 32319 5515 32353
rect 5457 32316 5515 32319
rect 7134 32316 7140 32328
rect 5457 32313 7140 32316
rect 5472 32288 7140 32313
rect 7134 32276 7140 32288
rect 7192 32276 7198 32328
rect 84322 32276 84328 32328
rect 84380 32316 84386 32328
rect 88235 32319 88293 32325
rect 88235 32316 88247 32319
rect 84380 32288 88247 32316
rect 84380 32276 84386 32288
rect 88235 32285 88247 32288
rect 88281 32285 88293 32319
rect 88235 32279 88293 32285
rect 88465 32319 88523 32325
rect 88465 32285 88477 32319
rect 88511 32316 88523 32319
rect 89934 32316 89940 32328
rect 88511 32288 89940 32316
rect 88511 32285 88523 32288
rect 88465 32279 88523 32285
rect 89934 32276 89940 32288
rect 89992 32276 89998 32328
rect 2902 32208 2908 32260
rect 2960 32248 2966 32260
rect 5251 32251 5309 32257
rect 5251 32248 5263 32251
rect 2960 32220 5263 32248
rect 2960 32208 2966 32220
rect 5251 32217 5263 32220
rect 5297 32217 5309 32251
rect 5251 32211 5309 32217
rect 4876 32122 7912 32144
rect 4876 32070 6690 32122
rect 6742 32070 6754 32122
rect 6806 32070 6818 32122
rect 6870 32070 6882 32122
rect 6934 32070 6946 32122
rect 6998 32070 7912 32122
rect 4876 32048 7912 32070
rect 86020 32122 88964 32144
rect 86020 32070 87834 32122
rect 87886 32070 87898 32122
rect 87950 32070 87962 32122
rect 88014 32070 88026 32122
rect 88078 32070 88090 32122
rect 88142 32070 88964 32122
rect 86020 32048 88964 32070
rect 4876 31578 7912 31600
rect 4876 31526 5954 31578
rect 6006 31526 6018 31578
rect 6070 31526 6082 31578
rect 6134 31526 6146 31578
rect 6198 31526 6210 31578
rect 6262 31526 7912 31578
rect 4876 31504 7912 31526
rect 86020 31578 88964 31600
rect 86020 31526 87098 31578
rect 87150 31526 87162 31578
rect 87214 31526 87226 31578
rect 87278 31526 87290 31578
rect 87342 31526 87354 31578
rect 87406 31526 88964 31578
rect 86020 31504 88964 31526
rect 5457 31265 5515 31271
rect 88554 31265 88560 31268
rect 5457 31231 5469 31265
rect 5503 31231 5515 31265
rect 88529 31259 88560 31265
rect 5457 31228 5515 31231
rect 7134 31228 7140 31240
rect 5457 31225 7140 31228
rect 5472 31200 7140 31225
rect 7134 31188 7140 31200
rect 7192 31188 7198 31240
rect 88529 31225 88541 31259
rect 88529 31219 88560 31225
rect 88554 31216 88560 31219
rect 88612 31216 88618 31268
rect 2902 31120 2908 31172
rect 2960 31160 2966 31172
rect 5251 31163 5309 31169
rect 5251 31160 5263 31163
rect 2960 31132 5263 31160
rect 2960 31120 2966 31132
rect 5251 31129 5263 31132
rect 5297 31129 5309 31163
rect 5251 31123 5309 31129
rect 84322 31120 84328 31172
rect 84380 31160 84386 31172
rect 88327 31163 88385 31169
rect 88327 31160 88339 31163
rect 84380 31132 88339 31160
rect 84380 31120 84386 31132
rect 88327 31129 88339 31132
rect 88373 31129 88385 31163
rect 88327 31123 88385 31129
rect 4876 31034 7912 31056
rect 4876 30982 6690 31034
rect 6742 30982 6754 31034
rect 6806 30982 6818 31034
rect 6870 30982 6882 31034
rect 6934 30982 6946 31034
rect 6998 30982 7912 31034
rect 4876 30960 7912 30982
rect 86020 31034 88964 31056
rect 86020 30982 87834 31034
rect 87886 30982 87898 31034
rect 87950 30982 87962 31034
rect 88014 30982 88026 31034
rect 88078 30982 88090 31034
rect 88142 30982 88964 31034
rect 86020 30960 88964 30982
rect 5457 30789 5515 30795
rect 5457 30755 5469 30789
rect 5503 30786 5515 30789
rect 5662 30786 5668 30798
rect 5503 30758 5668 30786
rect 5503 30755 5515 30758
rect 5457 30749 5515 30755
rect 5662 30746 5668 30758
rect 5720 30746 5726 30798
rect 88603 30771 88661 30777
rect 88603 30737 88615 30771
rect 88649 30768 88661 30771
rect 88649 30752 88876 30768
rect 89934 30752 89940 30764
rect 88649 30740 89940 30752
rect 88649 30737 88661 30740
rect 88603 30731 88661 30737
rect 88848 30724 89940 30740
rect 89934 30712 89940 30724
rect 89992 30712 89998 30764
rect 4374 30576 4380 30628
rect 4432 30616 4438 30628
rect 5251 30619 5309 30625
rect 5251 30616 5263 30619
rect 4432 30588 5263 30616
rect 4432 30576 4438 30588
rect 5251 30585 5263 30588
rect 5297 30585 5309 30619
rect 5251 30579 5309 30585
rect 87450 30576 87456 30628
rect 87508 30616 87514 30628
rect 88419 30619 88477 30625
rect 88419 30616 88431 30619
rect 87508 30588 88431 30616
rect 87508 30576 87514 30588
rect 88419 30585 88431 30588
rect 88465 30585 88477 30619
rect 88419 30579 88477 30585
rect 4876 30490 7912 30512
rect 4876 30438 5954 30490
rect 6006 30438 6018 30490
rect 6070 30438 6082 30490
rect 6134 30438 6146 30490
rect 6198 30438 6210 30490
rect 6262 30438 7912 30490
rect 4876 30416 7912 30438
rect 86020 30490 88964 30512
rect 86020 30438 87098 30490
rect 87150 30438 87162 30490
rect 87214 30438 87226 30490
rect 87278 30438 87290 30490
rect 87342 30438 87354 30490
rect 87406 30438 88964 30490
rect 86020 30416 88964 30438
rect 4876 29946 7912 29968
rect 4876 29894 6690 29946
rect 6742 29894 6754 29946
rect 6806 29894 6818 29946
rect 6870 29894 6882 29946
rect 6934 29894 6946 29946
rect 6998 29894 7912 29946
rect 4876 29872 7912 29894
rect 86020 29946 88964 29968
rect 86020 29894 87834 29946
rect 87886 29894 87898 29946
rect 87950 29894 87962 29946
rect 88014 29894 88026 29946
rect 88078 29894 88090 29946
rect 88142 29894 88964 29946
rect 86020 29872 88964 29894
rect 4876 29402 7912 29424
rect 4876 29350 5954 29402
rect 6006 29350 6018 29402
rect 6070 29350 6082 29402
rect 6134 29350 6146 29402
rect 6198 29350 6210 29402
rect 6262 29350 7912 29402
rect 4876 29328 7912 29350
rect 86020 29402 88964 29424
rect 86020 29350 87098 29402
rect 87150 29350 87162 29402
rect 87214 29350 87226 29402
rect 87278 29350 87290 29402
rect 87342 29350 87354 29402
rect 87406 29350 88964 29402
rect 86020 29328 88964 29350
rect 5457 29089 5515 29095
rect 88554 29089 88560 29092
rect 5457 29055 5469 29089
rect 5503 29055 5515 29089
rect 88529 29083 88560 29089
rect 5457 29052 5515 29055
rect 7134 29052 7140 29064
rect 5457 29049 7140 29052
rect 5472 29024 7140 29049
rect 7134 29012 7140 29024
rect 7192 29012 7198 29064
rect 88529 29049 88541 29083
rect 88529 29043 88560 29049
rect 88554 29040 88560 29043
rect 88612 29040 88618 29092
rect 2902 28944 2908 28996
rect 2960 28984 2966 28996
rect 5251 28987 5309 28993
rect 5251 28984 5263 28987
rect 2960 28956 5263 28984
rect 2960 28944 2966 28956
rect 5251 28953 5263 28956
rect 5297 28953 5309 28987
rect 5251 28947 5309 28953
rect 84322 28944 84328 28996
rect 84380 28984 84386 28996
rect 88327 28987 88385 28993
rect 88327 28984 88339 28987
rect 84380 28956 88339 28984
rect 84380 28944 84386 28956
rect 88327 28953 88339 28956
rect 88373 28953 88385 28987
rect 88327 28947 88385 28953
rect 4876 28858 7912 28880
rect 4876 28806 6690 28858
rect 6742 28806 6754 28858
rect 6806 28806 6818 28858
rect 6870 28806 6882 28858
rect 6934 28806 6946 28858
rect 6998 28806 7912 28858
rect 4876 28784 7912 28806
rect 86020 28858 88964 28880
rect 86020 28806 87834 28858
rect 87886 28806 87898 28858
rect 87950 28806 87962 28858
rect 88014 28806 88026 28858
rect 88078 28806 88090 28858
rect 88142 28806 88964 28858
rect 86020 28784 88964 28806
rect 4876 28314 7912 28336
rect 4876 28262 5954 28314
rect 6006 28262 6018 28314
rect 6070 28262 6082 28314
rect 6134 28262 6146 28314
rect 6198 28262 6210 28314
rect 6262 28262 7912 28314
rect 4876 28240 7912 28262
rect 86020 28314 88964 28336
rect 86020 28262 87098 28314
rect 87150 28262 87162 28314
rect 87214 28262 87226 28314
rect 87278 28262 87290 28314
rect 87342 28262 87354 28314
rect 87406 28262 88964 28314
rect 86020 28240 88964 28262
rect 5110 27958 5116 28010
rect 5168 27998 5174 28010
rect 5205 28001 5263 28007
rect 5205 27998 5217 28001
rect 5168 27970 5217 27998
rect 5168 27958 5174 27970
rect 5205 27967 5217 27970
rect 5251 27967 5263 28001
rect 88233 28001 88291 28007
rect 88233 27998 88245 28001
rect 5205 27961 5263 27967
rect 87542 27924 87548 27976
rect 87600 27964 87606 27976
rect 87928 27970 88245 27998
rect 87928 27964 87956 27970
rect 87600 27936 87956 27964
rect 88233 27967 88245 27970
rect 88279 27967 88291 28001
rect 88233 27961 88291 27967
rect 87600 27924 87606 27936
rect 5386 27905 5392 27908
rect 5364 27899 5392 27905
rect 5364 27865 5376 27899
rect 5364 27859 5392 27865
rect 5386 27856 5392 27859
rect 5444 27856 5450 27908
rect 88445 27899 88503 27905
rect 88445 27865 88457 27899
rect 88491 27896 88503 27899
rect 89934 27896 89940 27908
rect 88491 27868 89940 27896
rect 88491 27865 88503 27868
rect 88445 27859 88503 27865
rect 89934 27856 89940 27868
rect 89992 27856 89998 27908
rect 4876 27770 7912 27792
rect 4876 27718 6690 27770
rect 6742 27718 6754 27770
rect 6806 27718 6818 27770
rect 6870 27718 6882 27770
rect 6934 27718 6946 27770
rect 6998 27718 7912 27770
rect 4876 27696 7912 27718
rect 86020 27770 88964 27792
rect 86020 27718 87834 27770
rect 87886 27718 87898 27770
rect 87950 27718 87962 27770
rect 88014 27718 88026 27770
rect 88078 27718 88090 27770
rect 88142 27718 88964 27770
rect 86020 27696 88964 27718
rect 4876 27226 7912 27248
rect 4876 27174 5954 27226
rect 6006 27174 6018 27226
rect 6070 27174 6082 27226
rect 6134 27174 6146 27226
rect 6198 27174 6210 27226
rect 6262 27174 7912 27226
rect 4876 27152 7912 27174
rect 86020 27226 88964 27248
rect 86020 27174 87098 27226
rect 87150 27174 87162 27226
rect 87214 27174 87226 27226
rect 87278 27174 87290 27226
rect 87342 27174 87354 27226
rect 87406 27174 88964 27226
rect 86020 27152 88964 27174
rect 5159 26913 5217 26919
rect 2902 26836 2908 26888
rect 2960 26876 2966 26888
rect 5159 26879 5171 26913
rect 5205 26879 5217 26913
rect 88233 26913 88291 26919
rect 5159 26876 5217 26879
rect 2960 26873 5217 26876
rect 2960 26848 5202 26873
rect 2960 26836 2966 26848
rect 84322 26836 84328 26888
rect 84380 26876 84386 26888
rect 88233 26879 88245 26913
rect 88279 26879 88291 26913
rect 88233 26876 88291 26879
rect 84380 26873 88291 26876
rect 84380 26848 88276 26873
rect 84380 26836 84386 26848
rect 5364 26811 5422 26817
rect 5364 26777 5376 26811
rect 5410 26808 5422 26811
rect 7134 26808 7140 26820
rect 5410 26780 7140 26808
rect 5410 26777 5422 26780
rect 5364 26771 5422 26777
rect 7134 26768 7140 26780
rect 7192 26768 7198 26820
rect 88445 26811 88503 26817
rect 88445 26777 88457 26811
rect 88491 26808 88503 26811
rect 89934 26808 89940 26820
rect 88491 26780 89940 26808
rect 88491 26777 88503 26780
rect 88445 26771 88503 26777
rect 89934 26768 89940 26780
rect 89992 26768 89998 26820
rect 4876 26682 7912 26704
rect 4876 26630 6690 26682
rect 6742 26630 6754 26682
rect 6806 26630 6818 26682
rect 6870 26630 6882 26682
rect 6934 26630 6946 26682
rect 6998 26630 7912 26682
rect 4876 26608 7912 26630
rect 86020 26682 88964 26704
rect 86020 26630 87834 26682
rect 87886 26630 87898 26682
rect 87950 26630 87962 26682
rect 88014 26630 88026 26682
rect 88078 26630 88090 26682
rect 88142 26630 88964 26682
rect 86020 26608 88964 26630
rect 4876 26138 7912 26160
rect 4876 26086 5954 26138
rect 6006 26086 6018 26138
rect 6070 26086 6082 26138
rect 6134 26086 6146 26138
rect 6198 26086 6210 26138
rect 6262 26086 7912 26138
rect 4876 26064 7912 26086
rect 86020 26138 88964 26160
rect 86020 26086 87098 26138
rect 87150 26086 87162 26138
rect 87214 26086 87226 26138
rect 87278 26086 87290 26138
rect 87342 26086 87354 26138
rect 87406 26086 88964 26138
rect 86020 26064 88964 26086
rect 5159 25825 5217 25831
rect 2902 25748 2908 25800
rect 2960 25788 2966 25800
rect 5159 25791 5171 25825
rect 5205 25791 5217 25825
rect 88233 25825 88291 25831
rect 5159 25788 5217 25791
rect 2960 25785 5217 25788
rect 2960 25760 5202 25785
rect 2960 25748 2966 25760
rect 84322 25748 84328 25800
rect 84380 25788 84386 25800
rect 88233 25791 88245 25825
rect 88279 25791 88291 25825
rect 88233 25788 88291 25791
rect 84380 25785 88291 25788
rect 84380 25760 88276 25785
rect 84380 25748 84386 25760
rect 5364 25723 5422 25729
rect 5364 25689 5376 25723
rect 5410 25720 5422 25723
rect 7134 25720 7140 25732
rect 5410 25692 7140 25720
rect 5410 25689 5422 25692
rect 5364 25683 5422 25689
rect 7134 25680 7140 25692
rect 7192 25680 7198 25732
rect 88445 25723 88503 25729
rect 88445 25689 88457 25723
rect 88491 25720 88503 25723
rect 89934 25720 89940 25732
rect 88491 25692 89940 25720
rect 88491 25689 88503 25692
rect 88445 25683 88503 25689
rect 89934 25680 89940 25692
rect 89992 25680 89998 25732
rect 4876 25594 7912 25616
rect 4876 25542 6690 25594
rect 6742 25542 6754 25594
rect 6806 25542 6818 25594
rect 6870 25542 6882 25594
rect 6934 25542 6946 25594
rect 6998 25542 7912 25594
rect 4876 25520 7912 25542
rect 86020 25594 88964 25616
rect 86020 25542 87834 25594
rect 87886 25542 87898 25594
rect 87950 25542 87962 25594
rect 88014 25542 88026 25594
rect 88078 25542 88090 25594
rect 88142 25542 88964 25594
rect 86020 25520 88964 25542
rect 4926 25306 4932 25358
rect 4984 25346 4990 25358
rect 5159 25349 5217 25355
rect 5159 25346 5171 25349
rect 4984 25318 5171 25346
rect 4984 25306 4990 25318
rect 5159 25315 5171 25318
rect 5205 25315 5217 25349
rect 5159 25309 5217 25315
rect 88370 25306 88376 25358
rect 88428 25306 88434 25358
rect 5364 25179 5422 25185
rect 5364 25145 5376 25179
rect 5410 25176 5422 25179
rect 5662 25176 5668 25188
rect 5410 25148 5668 25176
rect 5410 25145 5422 25148
rect 5364 25139 5422 25145
rect 5662 25136 5668 25148
rect 5720 25136 5726 25188
rect 88537 25179 88595 25185
rect 88537 25145 88549 25179
rect 88583 25176 88595 25179
rect 89934 25176 89940 25188
rect 88583 25148 89940 25176
rect 88583 25145 88595 25148
rect 88537 25139 88595 25145
rect 89934 25136 89940 25148
rect 89992 25136 89998 25188
rect 4876 25050 7912 25072
rect 4876 24998 5954 25050
rect 6006 24998 6018 25050
rect 6070 24998 6082 25050
rect 6134 24998 6146 25050
rect 6198 24998 6210 25050
rect 6262 24998 7912 25050
rect 4876 24976 7912 24998
rect 86020 25050 88964 25072
rect 86020 24998 87098 25050
rect 87150 24998 87162 25050
rect 87214 24998 87226 25050
rect 87278 24998 87290 25050
rect 87342 24998 87354 25050
rect 87406 24998 88964 25050
rect 86020 24976 88964 24998
rect 4876 24506 7912 24528
rect 4876 24454 6690 24506
rect 6742 24454 6754 24506
rect 6806 24454 6818 24506
rect 6870 24454 6882 24506
rect 6934 24454 6946 24506
rect 6998 24454 7912 24506
rect 4876 24432 7912 24454
rect 86020 24506 88964 24528
rect 86020 24454 87834 24506
rect 87886 24454 87898 24506
rect 87950 24454 87962 24506
rect 88014 24454 88026 24506
rect 88078 24454 88090 24506
rect 88142 24454 88964 24506
rect 86020 24432 88964 24454
rect 4876 23962 7912 23984
rect 4876 23910 5954 23962
rect 6006 23910 6018 23962
rect 6070 23910 6082 23962
rect 6134 23910 6146 23962
rect 6198 23910 6210 23962
rect 6262 23910 7912 23962
rect 4876 23888 7912 23910
rect 86020 23962 88964 23984
rect 86020 23910 87098 23962
rect 87150 23910 87162 23962
rect 87214 23910 87226 23962
rect 87278 23910 87290 23962
rect 87342 23910 87354 23962
rect 87406 23910 88964 23962
rect 86020 23888 88964 23910
rect 5159 23649 5217 23655
rect 2902 23572 2908 23624
rect 2960 23612 2966 23624
rect 5159 23615 5171 23649
rect 5205 23615 5217 23649
rect 88233 23649 88291 23655
rect 5159 23612 5217 23615
rect 2960 23609 5217 23612
rect 2960 23584 5202 23609
rect 2960 23572 2966 23584
rect 84322 23572 84328 23624
rect 84380 23612 84386 23624
rect 88233 23615 88245 23649
rect 88279 23615 88291 23649
rect 88233 23612 88291 23615
rect 84380 23609 88291 23612
rect 84380 23584 88276 23609
rect 84380 23572 84386 23584
rect 5364 23547 5422 23553
rect 5364 23513 5376 23547
rect 5410 23544 5422 23547
rect 7134 23544 7140 23556
rect 5410 23516 7140 23544
rect 5410 23513 5422 23516
rect 5364 23507 5422 23513
rect 7134 23504 7140 23516
rect 7192 23504 7198 23556
rect 88445 23547 88503 23553
rect 88445 23513 88457 23547
rect 88491 23544 88503 23547
rect 89934 23544 89940 23556
rect 88491 23516 89940 23544
rect 88491 23513 88503 23516
rect 88445 23507 88503 23513
rect 89934 23504 89940 23516
rect 89992 23504 89998 23556
rect 4876 23418 7912 23440
rect 4876 23366 6690 23418
rect 6742 23366 6754 23418
rect 6806 23366 6818 23418
rect 6870 23366 6882 23418
rect 6934 23366 6946 23418
rect 6998 23366 7912 23418
rect 4876 23344 7912 23366
rect 86020 23418 88964 23440
rect 86020 23366 87834 23418
rect 87886 23366 87898 23418
rect 87950 23366 87962 23418
rect 88014 23366 88026 23418
rect 88078 23366 88090 23418
rect 88142 23366 88964 23418
rect 86020 23344 88964 23366
rect 4876 22874 7912 22896
rect 4876 22822 5954 22874
rect 6006 22822 6018 22874
rect 6070 22822 6082 22874
rect 6134 22822 6146 22874
rect 6198 22822 6210 22874
rect 6262 22822 7912 22874
rect 4876 22800 7912 22822
rect 86020 22874 88964 22896
rect 86020 22822 87098 22874
rect 87150 22822 87162 22874
rect 87214 22822 87226 22874
rect 87278 22822 87290 22874
rect 87342 22822 87354 22874
rect 87406 22822 88964 22874
rect 86020 22800 88964 22822
rect 5202 22518 5208 22570
rect 5260 22518 5266 22570
rect 88233 22561 88291 22567
rect 84322 22484 84328 22536
rect 84380 22524 84386 22536
rect 88233 22527 88245 22561
rect 88279 22527 88291 22561
rect 88233 22524 88291 22527
rect 84380 22521 88291 22524
rect 84380 22496 88276 22521
rect 84380 22484 84386 22496
rect 5364 22459 5422 22465
rect 5364 22425 5376 22459
rect 5410 22456 5422 22459
rect 7134 22456 7140 22468
rect 5410 22428 7140 22456
rect 5410 22425 5422 22428
rect 5364 22419 5422 22425
rect 7134 22416 7140 22428
rect 7192 22416 7198 22468
rect 88445 22459 88503 22465
rect 88445 22425 88457 22459
rect 88491 22456 88503 22459
rect 89934 22456 89940 22468
rect 88491 22428 89940 22456
rect 88491 22425 88503 22428
rect 88445 22419 88503 22425
rect 89934 22416 89940 22428
rect 89992 22416 89998 22468
rect 4876 22330 7912 22352
rect 4876 22278 6690 22330
rect 6742 22278 6754 22330
rect 6806 22278 6818 22330
rect 6870 22278 6882 22330
rect 6934 22278 6946 22330
rect 6998 22278 7912 22330
rect 4876 22256 7912 22278
rect 86020 22330 88964 22352
rect 86020 22278 87834 22330
rect 87886 22278 87898 22330
rect 87950 22278 87962 22330
rect 88014 22278 88026 22330
rect 88078 22278 88090 22330
rect 88142 22278 88964 22330
rect 86020 22256 88964 22278
rect 4876 21786 7912 21808
rect 4876 21734 5954 21786
rect 6006 21734 6018 21786
rect 6070 21734 6082 21786
rect 6134 21734 6146 21786
rect 6198 21734 6210 21786
rect 6262 21734 7912 21786
rect 4876 21712 7912 21734
rect 86020 21786 88964 21808
rect 86020 21734 87098 21786
rect 87150 21734 87162 21786
rect 87214 21734 87226 21786
rect 87278 21734 87290 21786
rect 87342 21734 87354 21786
rect 87406 21734 88964 21786
rect 86020 21712 88964 21734
rect 5159 21473 5217 21479
rect 2902 21396 2908 21448
rect 2960 21436 2966 21448
rect 5159 21439 5171 21473
rect 5205 21439 5217 21473
rect 88233 21473 88291 21479
rect 5159 21436 5217 21439
rect 2960 21433 5217 21436
rect 2960 21408 5202 21433
rect 2960 21396 2966 21408
rect 84322 21396 84328 21448
rect 84380 21436 84386 21448
rect 88233 21439 88245 21473
rect 88279 21439 88291 21473
rect 88233 21436 88291 21439
rect 84380 21433 88291 21436
rect 84380 21408 88276 21433
rect 84380 21396 84386 21408
rect 5364 21371 5422 21377
rect 5364 21337 5376 21371
rect 5410 21368 5422 21371
rect 7134 21368 7140 21380
rect 5410 21340 7140 21368
rect 5410 21337 5422 21340
rect 5364 21331 5422 21337
rect 7134 21328 7140 21340
rect 7192 21328 7198 21380
rect 88445 21371 88503 21377
rect 88445 21337 88457 21371
rect 88491 21368 88503 21371
rect 89934 21368 89940 21380
rect 88491 21340 89940 21368
rect 88491 21337 88503 21340
rect 88445 21331 88503 21337
rect 89934 21328 89940 21340
rect 89992 21328 89998 21380
rect 4876 21242 7912 21264
rect 4876 21190 6690 21242
rect 6742 21190 6754 21242
rect 6806 21190 6818 21242
rect 6870 21190 6882 21242
rect 6934 21190 6946 21242
rect 6998 21190 7912 21242
rect 4876 21168 7912 21190
rect 86020 21242 88964 21264
rect 86020 21190 87834 21242
rect 87886 21190 87898 21242
rect 87950 21190 87962 21242
rect 88014 21190 88026 21242
rect 88078 21190 88090 21242
rect 88142 21190 88964 21242
rect 86020 21168 88964 21190
rect 4876 20698 7912 20720
rect 4876 20646 5954 20698
rect 6006 20646 6018 20698
rect 6070 20646 6082 20698
rect 6134 20646 6146 20698
rect 6198 20646 6210 20698
rect 6262 20646 7912 20698
rect 4876 20624 7912 20646
rect 86020 20698 88964 20720
rect 86020 20646 87098 20698
rect 87150 20646 87162 20698
rect 87214 20646 87226 20698
rect 87278 20646 87290 20698
rect 87342 20646 87354 20698
rect 87406 20646 88964 20698
rect 86020 20624 88964 20646
rect 5159 20385 5217 20391
rect 2902 20308 2908 20360
rect 2960 20348 2966 20360
rect 5159 20351 5171 20385
rect 5205 20351 5217 20385
rect 88233 20385 88291 20391
rect 5159 20348 5217 20351
rect 2960 20345 5217 20348
rect 2960 20320 5202 20345
rect 2960 20308 2966 20320
rect 84322 20308 84328 20360
rect 84380 20348 84386 20360
rect 88233 20351 88245 20385
rect 88279 20351 88291 20385
rect 88233 20348 88291 20351
rect 84380 20345 88291 20348
rect 84380 20320 88276 20345
rect 84380 20308 84386 20320
rect 5364 20283 5422 20289
rect 5364 20249 5376 20283
rect 5410 20280 5422 20283
rect 7134 20280 7140 20292
rect 5410 20252 7140 20280
rect 5410 20249 5422 20252
rect 5364 20243 5422 20249
rect 7134 20240 7140 20252
rect 7192 20240 7198 20292
rect 88445 20283 88503 20289
rect 88445 20249 88457 20283
rect 88491 20280 88503 20283
rect 89934 20280 89940 20292
rect 88491 20252 89940 20280
rect 88491 20249 88503 20252
rect 88445 20243 88503 20249
rect 89934 20240 89940 20252
rect 89992 20240 89998 20292
rect 4876 20154 7912 20176
rect 4876 20102 6690 20154
rect 6742 20102 6754 20154
rect 6806 20102 6818 20154
rect 6870 20102 6882 20154
rect 6934 20102 6946 20154
rect 6998 20102 7912 20154
rect 4876 20080 7912 20102
rect 86020 20154 88964 20176
rect 86020 20102 87834 20154
rect 87886 20102 87898 20154
rect 87950 20102 87962 20154
rect 88014 20102 88026 20154
rect 88078 20102 88090 20154
rect 88142 20102 88964 20154
rect 86020 20080 88964 20102
rect 4926 19866 4932 19918
rect 4984 19906 4990 19918
rect 5159 19909 5217 19915
rect 5159 19906 5171 19909
rect 4984 19878 5171 19906
rect 4984 19866 4990 19878
rect 5159 19875 5171 19878
rect 5205 19875 5217 19909
rect 5159 19869 5217 19875
rect 88370 19866 88376 19918
rect 88428 19866 88434 19918
rect 5364 19739 5422 19745
rect 5364 19705 5376 19739
rect 5410 19736 5422 19739
rect 9618 19736 9624 19748
rect 5410 19708 9624 19736
rect 5410 19705 5422 19708
rect 5364 19699 5422 19705
rect 9618 19696 9624 19708
rect 9676 19696 9682 19748
rect 88537 19739 88595 19745
rect 88537 19705 88549 19739
rect 88583 19736 88595 19739
rect 90026 19736 90032 19748
rect 88583 19708 90032 19736
rect 88583 19705 88595 19708
rect 88537 19699 88595 19705
rect 90026 19696 90032 19708
rect 90084 19696 90090 19748
rect 4876 19610 7912 19632
rect 4876 19558 5954 19610
rect 6006 19558 6018 19610
rect 6070 19558 6082 19610
rect 6134 19558 6146 19610
rect 6198 19558 6210 19610
rect 6262 19558 7912 19610
rect 4876 19536 7912 19558
rect 86020 19610 88964 19632
rect 86020 19558 87098 19610
rect 87150 19558 87162 19610
rect 87214 19558 87226 19610
rect 87278 19558 87290 19610
rect 87342 19558 87354 19610
rect 87406 19558 88964 19610
rect 86020 19536 88964 19558
rect 4876 19066 7912 19088
rect 4876 19014 6690 19066
rect 6742 19014 6754 19066
rect 6806 19014 6818 19066
rect 6870 19014 6882 19066
rect 6934 19014 6946 19066
rect 6998 19014 7912 19066
rect 4876 18992 7912 19014
rect 86020 19066 88964 19088
rect 86020 19014 87834 19066
rect 87886 19014 87898 19066
rect 87950 19014 87962 19066
rect 88014 19014 88026 19066
rect 88078 19014 88090 19066
rect 88142 19014 88964 19066
rect 86020 18992 88964 19014
rect 4876 18522 7912 18544
rect 4876 18470 5954 18522
rect 6006 18470 6018 18522
rect 6070 18470 6082 18522
rect 6134 18470 6146 18522
rect 6198 18470 6210 18522
rect 6262 18470 7912 18522
rect 4876 18448 7912 18470
rect 86020 18522 88964 18544
rect 86020 18470 87098 18522
rect 87150 18470 87162 18522
rect 87214 18470 87226 18522
rect 87278 18470 87290 18522
rect 87342 18470 87354 18522
rect 87406 18470 88964 18522
rect 86020 18448 88964 18470
rect 5364 18243 5422 18249
rect 5110 18166 5116 18218
rect 5168 18206 5174 18218
rect 5205 18209 5263 18215
rect 5205 18206 5217 18209
rect 5168 18178 5217 18206
rect 5168 18166 5174 18178
rect 5205 18175 5217 18178
rect 5251 18175 5263 18209
rect 5364 18209 5376 18243
rect 5410 18240 5422 18243
rect 9618 18240 9624 18252
rect 5410 18212 9624 18240
rect 5410 18209 5422 18212
rect 5364 18203 5422 18209
rect 9618 18200 9624 18212
rect 9676 18200 9682 18252
rect 88445 18243 88503 18249
rect 5205 18169 5263 18175
rect 88186 18166 88192 18218
rect 88244 18206 88250 18218
rect 88281 18209 88339 18215
rect 88281 18206 88293 18209
rect 88244 18178 88293 18206
rect 88244 18166 88250 18178
rect 88281 18175 88293 18178
rect 88327 18175 88339 18209
rect 88445 18209 88457 18243
rect 88491 18240 88503 18243
rect 89934 18240 89940 18252
rect 88491 18212 89940 18240
rect 88491 18209 88503 18212
rect 88445 18203 88503 18209
rect 89934 18200 89940 18212
rect 89992 18200 89998 18252
rect 88281 18169 88339 18175
rect 4876 17978 7912 18000
rect 4876 17926 6690 17978
rect 6742 17926 6754 17978
rect 6806 17926 6818 17978
rect 6870 17926 6882 17978
rect 6934 17926 6946 17978
rect 6998 17926 7912 17978
rect 4876 17904 7912 17926
rect 86020 17978 88964 18000
rect 86020 17926 87834 17978
rect 87886 17926 87898 17978
rect 87950 17926 87962 17978
rect 88014 17926 88026 17978
rect 88078 17926 88090 17978
rect 88142 17926 88964 17978
rect 86020 17904 88964 17926
rect 4876 17434 7912 17456
rect 4876 17382 5954 17434
rect 6006 17382 6018 17434
rect 6070 17382 6082 17434
rect 6134 17382 6146 17434
rect 6198 17382 6210 17434
rect 6262 17382 7912 17434
rect 4876 17360 7912 17382
rect 86020 17434 88964 17456
rect 86020 17382 87098 17434
rect 87150 17382 87162 17434
rect 87214 17382 87226 17434
rect 87278 17382 87290 17434
rect 87342 17382 87354 17434
rect 87406 17382 88964 17434
rect 86020 17360 88964 17382
rect 5202 17078 5208 17130
rect 5260 17078 5266 17130
rect 88233 17121 88291 17127
rect 88233 17118 88245 17121
rect 84322 17044 84328 17096
rect 84380 17084 84386 17096
rect 87928 17090 88245 17118
rect 87928 17084 87956 17090
rect 84380 17056 87956 17084
rect 88233 17087 88245 17090
rect 88279 17087 88291 17121
rect 88233 17081 88291 17087
rect 84380 17044 84386 17056
rect 5364 17019 5422 17025
rect 5364 16985 5376 17019
rect 5410 17016 5422 17019
rect 7134 17016 7140 17028
rect 5410 16988 7140 17016
rect 5410 16985 5422 16988
rect 5364 16979 5422 16985
rect 7134 16976 7140 16988
rect 7192 16976 7198 17028
rect 88445 17019 88503 17025
rect 88445 16985 88457 17019
rect 88491 17016 88503 17019
rect 89934 17016 89940 17028
rect 88491 16988 89940 17016
rect 88491 16985 88503 16988
rect 88445 16979 88503 16985
rect 89934 16976 89940 16988
rect 89992 16976 89998 17028
rect 4876 16890 7912 16912
rect 4876 16838 6690 16890
rect 6742 16838 6754 16890
rect 6806 16838 6818 16890
rect 6870 16838 6882 16890
rect 6934 16838 6946 16890
rect 6998 16838 7912 16890
rect 4876 16816 7912 16838
rect 86020 16890 88964 16912
rect 86020 16838 87834 16890
rect 87886 16838 87898 16890
rect 87950 16838 87962 16890
rect 88014 16838 88026 16890
rect 88078 16838 88090 16890
rect 88142 16838 88964 16890
rect 86020 16816 88964 16838
rect 4876 16346 7912 16368
rect 4876 16294 5954 16346
rect 6006 16294 6018 16346
rect 6070 16294 6082 16346
rect 6134 16294 6146 16346
rect 6198 16294 6210 16346
rect 6262 16294 7912 16346
rect 4876 16272 7912 16294
rect 86020 16346 88964 16368
rect 86020 16294 87098 16346
rect 87150 16294 87162 16346
rect 87214 16294 87226 16346
rect 87278 16294 87290 16346
rect 87342 16294 87354 16346
rect 87406 16294 88964 16346
rect 86020 16272 88964 16294
rect 5159 16033 5217 16039
rect 5159 16030 5171 16033
rect 2902 15956 2908 16008
rect 2960 15996 2966 16008
rect 4852 16002 5171 16030
rect 4852 15996 4880 16002
rect 2960 15968 4880 15996
rect 5159 15999 5171 16002
rect 5205 15999 5217 16033
rect 88233 16033 88291 16039
rect 88233 16030 88245 16033
rect 5159 15993 5217 15999
rect 2960 15956 2966 15968
rect 84322 15956 84328 16008
rect 84380 15996 84386 16008
rect 87928 16002 88245 16030
rect 87928 15996 87956 16002
rect 84380 15968 87956 15996
rect 88233 15999 88245 16002
rect 88279 15999 88291 16033
rect 88233 15993 88291 15999
rect 84380 15956 84386 15968
rect 5365 15931 5423 15937
rect 5365 15897 5377 15931
rect 5411 15928 5423 15931
rect 7594 15928 7600 15940
rect 5411 15900 7600 15928
rect 5411 15897 5423 15900
rect 5365 15891 5423 15897
rect 7594 15888 7600 15900
rect 7652 15888 7658 15940
rect 88445 15931 88503 15937
rect 88445 15897 88457 15931
rect 88491 15928 88503 15931
rect 89934 15928 89940 15940
rect 88491 15900 89940 15928
rect 88491 15897 88503 15900
rect 88445 15891 88503 15897
rect 89934 15888 89940 15900
rect 89992 15888 89998 15940
rect 4876 15802 7912 15824
rect 4876 15750 6690 15802
rect 6742 15750 6754 15802
rect 6806 15750 6818 15802
rect 6870 15750 6882 15802
rect 6934 15750 6946 15802
rect 6998 15750 7912 15802
rect 4876 15728 7912 15750
rect 86020 15802 88964 15824
rect 86020 15750 87834 15802
rect 87886 15750 87898 15802
rect 87950 15750 87962 15802
rect 88014 15750 88026 15802
rect 88078 15750 88090 15802
rect 88142 15750 88964 15802
rect 86020 15728 88964 15750
rect 4876 15258 7912 15280
rect 4876 15206 5954 15258
rect 6006 15206 6018 15258
rect 6070 15206 6082 15258
rect 6134 15206 6146 15258
rect 6198 15206 6210 15258
rect 6262 15206 7912 15258
rect 4876 15184 7912 15206
rect 86020 15258 88964 15280
rect 86020 15206 87098 15258
rect 87150 15206 87162 15258
rect 87214 15206 87226 15258
rect 87278 15206 87290 15258
rect 87342 15206 87354 15258
rect 87406 15206 88964 15258
rect 86020 15184 88964 15206
rect 5159 14945 5217 14951
rect 5159 14942 5171 14945
rect 2902 14868 2908 14920
rect 2960 14908 2966 14920
rect 4852 14914 5171 14942
rect 4852 14908 4880 14914
rect 2960 14880 4880 14908
rect 5159 14911 5171 14914
rect 5205 14911 5217 14945
rect 88233 14945 88291 14951
rect 88233 14942 88245 14945
rect 5159 14905 5217 14911
rect 2960 14868 2966 14880
rect 84322 14868 84328 14920
rect 84380 14908 84386 14920
rect 87928 14914 88245 14942
rect 87928 14908 87956 14914
rect 84380 14880 87956 14908
rect 88233 14911 88245 14914
rect 88279 14911 88291 14945
rect 88233 14905 88291 14911
rect 84380 14868 84386 14880
rect 5365 14843 5423 14849
rect 5365 14809 5377 14843
rect 5411 14840 5423 14843
rect 7594 14840 7600 14852
rect 5411 14812 7600 14840
rect 5411 14809 5423 14812
rect 5365 14803 5423 14809
rect 7594 14800 7600 14812
rect 7652 14800 7658 14852
rect 88445 14843 88503 14849
rect 88445 14809 88457 14843
rect 88491 14840 88503 14843
rect 89934 14840 89940 14852
rect 88491 14812 89940 14840
rect 88491 14809 88503 14812
rect 88445 14803 88503 14809
rect 89934 14800 89940 14812
rect 89992 14800 89998 14852
rect 4876 14714 7912 14736
rect 4876 14662 6690 14714
rect 6742 14662 6754 14714
rect 6806 14662 6818 14714
rect 6870 14662 6882 14714
rect 6934 14662 6946 14714
rect 6998 14662 7912 14714
rect 4876 14640 7912 14662
rect 86020 14714 88964 14736
rect 86020 14662 87834 14714
rect 87886 14662 87898 14714
rect 87950 14662 87962 14714
rect 88014 14662 88026 14714
rect 88078 14662 88090 14714
rect 88142 14662 88964 14714
rect 86020 14640 88964 14662
rect 4926 14426 4932 14478
rect 4984 14466 4990 14478
rect 5159 14469 5217 14475
rect 5159 14466 5171 14469
rect 4984 14438 5171 14466
rect 4984 14426 4990 14438
rect 5159 14435 5171 14438
rect 5205 14435 5217 14469
rect 5159 14429 5217 14435
rect 88370 14426 88376 14478
rect 88428 14426 88434 14478
rect 5364 14299 5422 14305
rect 5364 14265 5376 14299
rect 5410 14296 5422 14299
rect 5662 14296 5668 14308
rect 5410 14268 5668 14296
rect 5410 14265 5422 14268
rect 5364 14259 5422 14265
rect 5662 14256 5668 14268
rect 5720 14256 5726 14308
rect 88537 14299 88595 14305
rect 88537 14265 88549 14299
rect 88583 14296 88595 14299
rect 89934 14296 89940 14308
rect 88583 14268 89940 14296
rect 88583 14265 88595 14268
rect 88537 14259 88595 14265
rect 89934 14256 89940 14268
rect 89992 14256 89998 14308
rect 4876 14170 7912 14192
rect 4876 14118 5954 14170
rect 6006 14118 6018 14170
rect 6070 14118 6082 14170
rect 6134 14118 6146 14170
rect 6198 14118 6210 14170
rect 6262 14118 7912 14170
rect 4876 14096 7912 14118
rect 86020 14170 88964 14192
rect 86020 14118 87098 14170
rect 87150 14118 87162 14170
rect 87214 14118 87226 14170
rect 87278 14118 87290 14170
rect 87342 14118 87354 14170
rect 87406 14118 88964 14170
rect 86020 14096 88964 14118
rect 4876 13626 7912 13648
rect 4876 13574 6690 13626
rect 6742 13574 6754 13626
rect 6806 13574 6818 13626
rect 6870 13574 6882 13626
rect 6934 13574 6946 13626
rect 6998 13574 7912 13626
rect 4876 13552 7912 13574
rect 86020 13626 88964 13648
rect 86020 13574 87834 13626
rect 87886 13574 87898 13626
rect 87950 13574 87962 13626
rect 88014 13574 88026 13626
rect 88078 13574 88090 13626
rect 88142 13574 88964 13626
rect 86020 13552 88964 13574
rect 4876 13082 7912 13104
rect 4876 13030 5954 13082
rect 6006 13030 6018 13082
rect 6070 13030 6082 13082
rect 6134 13030 6146 13082
rect 6198 13030 6210 13082
rect 6262 13030 7912 13082
rect 4876 13008 7912 13030
rect 86020 13082 88964 13104
rect 86020 13030 87098 13082
rect 87150 13030 87162 13082
rect 87214 13030 87226 13082
rect 87278 13030 87290 13082
rect 87342 13030 87354 13082
rect 87406 13030 88964 13082
rect 86020 13008 88964 13030
rect 4876 12538 7912 12560
rect 4876 12486 6690 12538
rect 6742 12486 6754 12538
rect 6806 12486 6818 12538
rect 6870 12486 6882 12538
rect 6934 12486 6946 12538
rect 6998 12486 7912 12538
rect 4876 12464 7912 12486
rect 86020 12538 88964 12560
rect 86020 12486 87834 12538
rect 87886 12486 87898 12538
rect 87950 12486 87962 12538
rect 88014 12486 88026 12538
rect 88078 12486 88090 12538
rect 88142 12486 88964 12538
rect 86020 12464 88964 12486
rect 4876 11994 7912 12016
rect 4876 11942 5954 11994
rect 6006 11942 6018 11994
rect 6070 11942 6082 11994
rect 6134 11942 6146 11994
rect 6198 11942 6210 11994
rect 6262 11942 7912 11994
rect 4876 11920 7912 11942
rect 86020 11994 88964 12016
rect 86020 11942 87098 11994
rect 87150 11942 87162 11994
rect 87214 11942 87226 11994
rect 87278 11942 87290 11994
rect 87342 11942 87354 11994
rect 87406 11942 88964 11994
rect 86020 11920 88964 11942
rect 4876 11450 7912 11472
rect 4876 11398 6690 11450
rect 6742 11398 6754 11450
rect 6806 11398 6818 11450
rect 6870 11398 6882 11450
rect 6934 11398 6946 11450
rect 6998 11398 7912 11450
rect 4876 11376 7912 11398
rect 86020 11450 88964 11472
rect 86020 11398 87834 11450
rect 87886 11398 87898 11450
rect 87950 11398 87962 11450
rect 88014 11398 88026 11450
rect 88078 11398 88090 11450
rect 88142 11398 88964 11450
rect 86020 11376 88964 11398
rect 4876 10906 7912 10928
rect 4876 10854 5954 10906
rect 6006 10854 6018 10906
rect 6070 10854 6082 10906
rect 6134 10854 6146 10906
rect 6198 10854 6210 10906
rect 6262 10854 7912 10906
rect 4876 10832 7912 10854
rect 86020 10906 88964 10928
rect 86020 10854 87098 10906
rect 87150 10854 87162 10906
rect 87214 10854 87226 10906
rect 87278 10854 87290 10906
rect 87342 10854 87354 10906
rect 87406 10854 88964 10906
rect 86020 10832 88964 10854
rect 4876 10362 7912 10384
rect 4876 10310 6690 10362
rect 6742 10310 6754 10362
rect 6806 10310 6818 10362
rect 6870 10310 6882 10362
rect 6934 10310 6946 10362
rect 6998 10310 7912 10362
rect 4876 10288 7912 10310
rect 86020 10362 88964 10384
rect 86020 10310 87834 10362
rect 87886 10310 87898 10362
rect 87950 10310 87962 10362
rect 88014 10310 88026 10362
rect 88078 10310 88090 10362
rect 88142 10310 88964 10362
rect 86020 10288 88964 10310
rect 4876 9818 7912 9840
rect 4876 9766 5954 9818
rect 6006 9766 6018 9818
rect 6070 9766 6082 9818
rect 6134 9766 6146 9818
rect 6198 9766 6210 9818
rect 6262 9766 7912 9818
rect 4876 9744 7912 9766
rect 86020 9818 88964 9840
rect 86020 9766 87098 9818
rect 87150 9766 87162 9818
rect 87214 9766 87226 9818
rect 87278 9766 87290 9818
rect 87342 9766 87354 9818
rect 87406 9766 88964 9818
rect 86020 9744 88964 9766
rect 4876 9274 7912 9296
rect 4876 9222 6690 9274
rect 6742 9222 6754 9274
rect 6806 9222 6818 9274
rect 6870 9222 6882 9274
rect 6934 9222 6946 9274
rect 6998 9222 7912 9274
rect 4876 9200 7912 9222
rect 86020 9274 88964 9296
rect 86020 9222 87834 9274
rect 87886 9222 87898 9274
rect 87950 9222 87962 9274
rect 88014 9222 88026 9274
rect 88078 9222 88090 9274
rect 88142 9222 88964 9274
rect 86020 9200 88964 9222
rect 4876 8730 7912 8752
rect 4876 8678 5954 8730
rect 6006 8678 6018 8730
rect 6070 8678 6082 8730
rect 6134 8678 6146 8730
rect 6198 8678 6210 8730
rect 6262 8678 7912 8730
rect 4876 8656 7912 8678
rect 86020 8730 88964 8752
rect 86020 8678 87098 8730
rect 87150 8678 87162 8730
rect 87214 8678 87226 8730
rect 87278 8678 87290 8730
rect 87342 8678 87354 8730
rect 87406 8678 88964 8730
rect 86020 8656 88964 8678
rect 4876 8186 7912 8208
rect 4876 8134 6690 8186
rect 6742 8134 6754 8186
rect 6806 8134 6818 8186
rect 6870 8134 6882 8186
rect 6934 8134 6946 8186
rect 6998 8134 7912 8186
rect 4876 8112 7912 8134
rect 86020 8186 88964 8208
rect 86020 8134 87834 8186
rect 87886 8134 87898 8186
rect 87950 8134 87962 8186
rect 88014 8134 88026 8186
rect 88078 8134 88090 8186
rect 88142 8134 88964 8186
rect 86020 8112 88964 8134
rect 4876 7642 88964 7664
rect 4876 7590 5954 7642
rect 6006 7590 6018 7642
rect 6070 7590 6082 7642
rect 6134 7590 6146 7642
rect 6198 7590 6210 7642
rect 6262 7590 18722 7642
rect 18774 7590 18786 7642
rect 18838 7590 18850 7642
rect 18902 7590 18914 7642
rect 18966 7590 18978 7642
rect 19030 7590 37722 7642
rect 37774 7590 37786 7642
rect 37838 7590 37850 7642
rect 37902 7590 37914 7642
rect 37966 7590 37978 7642
rect 38030 7590 56722 7642
rect 56774 7590 56786 7642
rect 56838 7590 56850 7642
rect 56902 7590 56914 7642
rect 56966 7590 56978 7642
rect 57030 7590 75722 7642
rect 75774 7590 75786 7642
rect 75838 7590 75850 7642
rect 75902 7590 75914 7642
rect 75966 7590 75978 7642
rect 76030 7590 87098 7642
rect 87150 7590 87162 7642
rect 87214 7590 87226 7642
rect 87278 7590 87290 7642
rect 87342 7590 87354 7642
rect 87406 7590 88964 7642
rect 4876 7568 88964 7590
rect 4876 7098 88964 7120
rect 4876 7046 6690 7098
rect 6742 7046 6754 7098
rect 6806 7046 6818 7098
rect 6870 7046 6882 7098
rect 6934 7046 6946 7098
rect 6998 7046 19382 7098
rect 19434 7046 19446 7098
rect 19498 7046 19510 7098
rect 19562 7046 19574 7098
rect 19626 7046 19638 7098
rect 19690 7046 38382 7098
rect 38434 7046 38446 7098
rect 38498 7046 38510 7098
rect 38562 7046 38574 7098
rect 38626 7046 38638 7098
rect 38690 7046 57382 7098
rect 57434 7046 57446 7098
rect 57498 7046 57510 7098
rect 57562 7046 57574 7098
rect 57626 7046 57638 7098
rect 57690 7046 76382 7098
rect 76434 7046 76446 7098
rect 76498 7046 76510 7098
rect 76562 7046 76574 7098
rect 76626 7046 76638 7098
rect 76690 7046 87834 7098
rect 87886 7046 87898 7098
rect 87950 7046 87962 7098
rect 88014 7046 88026 7098
rect 88078 7046 88090 7098
rect 88142 7046 88964 7098
rect 4876 7024 88964 7046
rect 4876 6554 88964 6576
rect 4876 6502 18722 6554
rect 18774 6502 18786 6554
rect 18838 6502 18850 6554
rect 18902 6502 18914 6554
rect 18966 6502 18978 6554
rect 19030 6502 37722 6554
rect 37774 6502 37786 6554
rect 37838 6502 37850 6554
rect 37902 6502 37914 6554
rect 37966 6502 37978 6554
rect 38030 6502 56722 6554
rect 56774 6502 56786 6554
rect 56838 6502 56850 6554
rect 56902 6502 56914 6554
rect 56966 6502 56978 6554
rect 57030 6502 75722 6554
rect 75774 6502 75786 6554
rect 75838 6502 75850 6554
rect 75902 6502 75914 6554
rect 75966 6502 75978 6554
rect 76030 6502 88964 6554
rect 4876 6480 88964 6502
rect 4876 6010 88964 6032
rect 4876 5958 19382 6010
rect 19434 5958 19446 6010
rect 19498 5958 19510 6010
rect 19562 5958 19574 6010
rect 19626 5958 19638 6010
rect 19690 5958 38382 6010
rect 38434 5958 38446 6010
rect 38498 5958 38510 6010
rect 38562 5958 38574 6010
rect 38626 5958 38638 6010
rect 38690 5958 57382 6010
rect 57434 5958 57446 6010
rect 57498 5958 57510 6010
rect 57562 5958 57574 6010
rect 57626 5958 57638 6010
rect 57690 5958 76382 6010
rect 76434 5958 76446 6010
rect 76498 5958 76510 6010
rect 76562 5958 76574 6010
rect 76626 5958 76638 6010
rect 76690 5958 88964 6010
rect 4876 5936 88964 5958
rect 82114 5688 82120 5740
rect 82172 5728 82178 5740
rect 82301 5731 82359 5737
rect 82301 5728 82313 5731
rect 82172 5700 82313 5728
rect 82172 5688 82178 5700
rect 82301 5697 82313 5700
rect 82347 5697 82359 5731
rect 82301 5691 82359 5697
rect 82390 5620 82396 5672
rect 82448 5660 82454 5672
rect 82485 5663 82543 5669
rect 82485 5660 82497 5663
rect 82448 5632 82497 5660
rect 82448 5620 82454 5632
rect 82485 5629 82497 5632
rect 82531 5629 82543 5663
rect 82485 5623 82543 5629
rect 4876 5466 88964 5488
rect 4876 5414 18722 5466
rect 18774 5414 18786 5466
rect 18838 5414 18850 5466
rect 18902 5414 18914 5466
rect 18966 5414 18978 5466
rect 19030 5414 37722 5466
rect 37774 5414 37786 5466
rect 37838 5414 37850 5466
rect 37902 5414 37914 5466
rect 37966 5414 37978 5466
rect 38030 5414 56722 5466
rect 56774 5414 56786 5466
rect 56838 5414 56850 5466
rect 56902 5414 56914 5466
rect 56966 5414 56978 5466
rect 57030 5414 75722 5466
rect 75774 5414 75786 5466
rect 75838 5414 75850 5466
rect 75902 5414 75914 5466
rect 75966 5414 75978 5466
rect 76030 5414 88964 5466
rect 4876 5392 88964 5414
rect 12654 5280 12660 5332
rect 12712 5320 12718 5332
rect 13485 5323 13543 5329
rect 13485 5320 13497 5323
rect 12712 5292 13497 5320
rect 12712 5280 12718 5292
rect 13485 5289 13497 5292
rect 13531 5289 13543 5323
rect 13485 5283 13543 5289
rect 14678 5280 14684 5332
rect 14736 5280 14742 5332
rect 30962 5280 30968 5332
rect 31020 5320 31026 5332
rect 31287 5323 31345 5329
rect 31287 5320 31299 5323
rect 31020 5292 31299 5320
rect 31020 5280 31026 5292
rect 31287 5289 31299 5292
rect 31333 5289 31345 5323
rect 31287 5283 31345 5289
rect 33170 5280 33176 5332
rect 33228 5320 33234 5332
rect 33311 5323 33369 5329
rect 33311 5320 33323 5323
rect 33228 5292 33323 5320
rect 33228 5280 33234 5292
rect 33311 5289 33323 5292
rect 33357 5289 33369 5323
rect 33311 5283 33369 5289
rect 34274 5280 34280 5332
rect 34332 5320 34338 5332
rect 35378 5329 35384 5332
rect 34507 5323 34565 5329
rect 34507 5320 34519 5323
rect 34332 5292 34519 5320
rect 34332 5280 34338 5292
rect 34507 5289 34519 5292
rect 34553 5289 34565 5323
rect 34507 5283 34565 5289
rect 35356 5323 35384 5329
rect 35356 5289 35368 5323
rect 35356 5283 35384 5289
rect 35378 5280 35384 5283
rect 35436 5280 35442 5332
rect 36482 5280 36488 5332
rect 36540 5320 36546 5332
rect 36635 5323 36693 5329
rect 36635 5320 36647 5323
rect 36540 5292 36647 5320
rect 36540 5280 36546 5292
rect 36635 5289 36647 5292
rect 36681 5289 36693 5323
rect 36635 5283 36693 5289
rect 37586 5280 37592 5332
rect 37644 5320 37650 5332
rect 37727 5323 37785 5329
rect 37727 5320 37739 5323
rect 37644 5292 37739 5320
rect 37644 5280 37650 5292
rect 37727 5289 37739 5292
rect 37773 5289 37785 5323
rect 37727 5283 37785 5289
rect 38782 5280 38788 5332
rect 38840 5320 38846 5332
rect 39015 5323 39073 5329
rect 39015 5320 39027 5323
rect 38840 5292 39027 5320
rect 38840 5280 38846 5292
rect 39015 5289 39027 5292
rect 39061 5289 39073 5323
rect 39015 5283 39073 5289
rect 40898 5280 40904 5332
rect 40956 5320 40962 5332
rect 41039 5323 41097 5329
rect 41039 5320 41051 5323
rect 40956 5292 41051 5320
rect 40956 5280 40962 5292
rect 41039 5289 41051 5292
rect 41085 5289 41097 5323
rect 41039 5283 41097 5289
rect 44210 5280 44216 5332
rect 44268 5320 44274 5332
rect 44397 5323 44455 5329
rect 44397 5320 44409 5323
rect 44268 5292 44409 5320
rect 44268 5280 44274 5292
rect 44397 5289 44409 5292
rect 44443 5289 44455 5323
rect 44397 5283 44455 5289
rect 45314 5280 45320 5332
rect 45372 5320 45378 5332
rect 68038 5329 68044 5332
rect 46421 5323 46479 5329
rect 46421 5320 46433 5323
rect 45372 5292 46433 5320
rect 45372 5280 45378 5292
rect 46421 5289 46433 5292
rect 46467 5289 46479 5323
rect 46421 5283 46479 5289
rect 67995 5323 68044 5329
rect 67995 5289 68007 5323
rect 68041 5289 68044 5323
rect 67995 5283 68044 5289
rect 68038 5280 68044 5283
rect 68096 5280 68102 5332
rect 69326 5280 69332 5332
rect 69384 5329 69390 5332
rect 70154 5329 70160 5332
rect 69384 5323 69433 5329
rect 69384 5289 69387 5323
rect 69421 5289 69433 5323
rect 69384 5283 69433 5289
rect 70132 5323 70160 5329
rect 70132 5289 70144 5323
rect 70132 5283 70160 5289
rect 69384 5280 69390 5283
rect 70154 5280 70160 5283
rect 70212 5280 70218 5332
rect 72454 5280 72460 5332
rect 72512 5329 72518 5332
rect 72512 5323 72561 5329
rect 72512 5289 72515 5323
rect 72549 5289 72561 5323
rect 72512 5283 72561 5289
rect 72512 5280 72518 5283
rect 73558 5280 73564 5332
rect 73616 5320 73622 5332
rect 74754 5329 74760 5332
rect 73791 5323 73849 5329
rect 73791 5320 73803 5323
rect 73616 5292 73803 5320
rect 73616 5280 73622 5292
rect 73791 5289 73803 5292
rect 73837 5289 73849 5323
rect 73791 5283 73849 5289
rect 74732 5323 74760 5329
rect 74732 5289 74744 5323
rect 74732 5283 74760 5289
rect 74754 5280 74760 5283
rect 74812 5280 74818 5332
rect 75582 5280 75588 5332
rect 75640 5320 75646 5332
rect 75723 5323 75781 5329
rect 75723 5320 75735 5323
rect 75640 5292 75735 5320
rect 75640 5280 75646 5292
rect 75723 5289 75735 5292
rect 75769 5289 75781 5323
rect 75723 5283 75781 5289
rect 76870 5280 76876 5332
rect 76928 5320 76934 5332
rect 77882 5329 77888 5332
rect 77103 5323 77161 5329
rect 77103 5320 77115 5323
rect 76928 5292 77115 5320
rect 76928 5280 76934 5292
rect 77103 5289 77115 5292
rect 77149 5289 77161 5323
rect 77103 5283 77161 5289
rect 77860 5323 77888 5329
rect 77860 5289 77872 5323
rect 77860 5283 77888 5289
rect 77882 5280 77888 5283
rect 77940 5280 77946 5332
rect 81654 5280 81660 5332
rect 81712 5320 81718 5332
rect 82485 5323 82543 5329
rect 82485 5320 82497 5323
rect 81712 5292 82497 5320
rect 81712 5280 81718 5292
rect 82485 5289 82497 5292
rect 82531 5289 82543 5323
rect 82485 5283 82543 5289
rect 32066 5212 32072 5264
rect 32124 5261 32130 5264
rect 32124 5255 32173 5261
rect 32124 5221 32127 5255
rect 32161 5221 32173 5255
rect 32124 5215 32173 5221
rect 32124 5212 32130 5215
rect 39794 5212 39800 5264
rect 39852 5261 39858 5264
rect 39852 5255 39901 5261
rect 39852 5221 39855 5255
rect 39889 5221 39901 5255
rect 39852 5215 39901 5221
rect 39852 5212 39858 5215
rect 42002 5212 42008 5264
rect 42060 5252 42066 5264
rect 42235 5255 42293 5261
rect 42235 5252 42247 5255
rect 42060 5224 42247 5252
rect 42060 5212 42066 5224
rect 42235 5221 42247 5224
rect 42281 5221 42293 5255
rect 42235 5215 42293 5221
rect 43106 5212 43112 5264
rect 43164 5261 43170 5264
rect 43164 5255 43213 5261
rect 43164 5221 43167 5255
rect 43201 5221 43213 5255
rect 43164 5215 43213 5221
rect 43164 5212 43170 5215
rect 71350 5212 71356 5264
rect 71408 5261 71414 5264
rect 71408 5255 71457 5261
rect 71408 5221 71411 5255
rect 71445 5221 71457 5255
rect 71408 5215 71457 5221
rect 71408 5212 71414 5215
rect 79078 5212 79084 5264
rect 79136 5252 79142 5264
rect 80274 5261 80280 5264
rect 79219 5255 79277 5261
rect 79219 5252 79231 5255
rect 79136 5224 79231 5252
rect 79136 5212 79142 5224
rect 79219 5221 79231 5224
rect 79265 5221 79277 5255
rect 79219 5215 79277 5221
rect 80231 5255 80280 5261
rect 80231 5221 80243 5255
rect 80277 5221 80280 5255
rect 80231 5215 80280 5221
rect 80274 5212 80280 5215
rect 80332 5212 80338 5264
rect 15278 5153 15336 5159
rect 15278 5150 15290 5153
rect 12562 5076 12568 5128
rect 12620 5116 12626 5128
rect 12701 5119 12759 5125
rect 12701 5116 12713 5119
rect 12620 5088 12713 5116
rect 12620 5076 12626 5088
rect 12701 5085 12713 5088
rect 12747 5085 12759 5119
rect 12701 5079 12759 5085
rect 13850 5076 13856 5128
rect 13908 5125 13914 5128
rect 13908 5119 13955 5125
rect 13908 5085 13909 5119
rect 13943 5085 13955 5119
rect 13908 5079 13955 5085
rect 13908 5076 13914 5079
rect 14494 5076 14500 5128
rect 14552 5116 14558 5128
rect 14972 5122 15290 5150
rect 14972 5116 15000 5122
rect 14552 5088 15000 5116
rect 15278 5119 15290 5122
rect 15324 5119 15336 5153
rect 15506 5144 15512 5196
rect 15564 5184 15570 5196
rect 15564 5156 15736 5184
rect 15564 5144 15570 5156
rect 15708 5150 15736 5156
rect 15829 5153 15887 5159
rect 15829 5150 15841 5153
rect 15278 5113 15336 5119
rect 14552 5076 14558 5088
rect 15414 5076 15420 5128
rect 15472 5116 15478 5128
rect 15601 5119 15659 5125
rect 15708 5122 15841 5150
rect 15601 5116 15613 5119
rect 15472 5088 15613 5116
rect 15472 5076 15478 5088
rect 15601 5085 15613 5088
rect 15647 5085 15659 5119
rect 15829 5119 15841 5122
rect 15875 5119 15887 5153
rect 15829 5113 15887 5119
rect 16610 5110 16616 5162
rect 16668 5150 16674 5162
rect 16736 5153 16794 5159
rect 16736 5150 16748 5153
rect 16668 5122 16748 5150
rect 16668 5110 16674 5122
rect 16736 5119 16748 5122
rect 16782 5119 16794 5153
rect 16736 5113 16794 5119
rect 17714 5110 17720 5162
rect 17772 5150 17778 5162
rect 17853 5153 17911 5159
rect 17853 5150 17865 5153
rect 17772 5122 17865 5150
rect 17772 5110 17778 5122
rect 17853 5119 17865 5122
rect 17899 5119 17911 5153
rect 17853 5113 17911 5119
rect 19094 5110 19100 5162
rect 19152 5110 19158 5162
rect 19922 5110 19928 5162
rect 19980 5159 19986 5162
rect 19980 5153 20014 5159
rect 20002 5119 20014 5153
rect 19980 5113 20014 5119
rect 19980 5110 19986 5113
rect 21026 5110 21032 5162
rect 21084 5110 21090 5162
rect 22130 5110 22136 5162
rect 22188 5150 22194 5162
rect 22271 5153 22329 5159
rect 22271 5150 22283 5153
rect 22188 5122 22283 5150
rect 22188 5110 22194 5122
rect 22271 5119 22283 5122
rect 22317 5119 22329 5153
rect 22271 5113 22329 5119
rect 23326 5110 23332 5162
rect 23384 5150 23390 5162
rect 23557 5153 23615 5159
rect 23557 5150 23569 5153
rect 23384 5122 23569 5150
rect 23384 5110 23390 5122
rect 23557 5119 23569 5122
rect 23603 5119 23615 5153
rect 23557 5113 23615 5119
rect 24338 5110 24344 5162
rect 24396 5150 24402 5162
rect 24464 5153 24522 5159
rect 24464 5150 24476 5153
rect 24396 5122 24476 5150
rect 24396 5110 24402 5122
rect 24464 5119 24476 5122
rect 24510 5119 24522 5153
rect 24464 5113 24522 5119
rect 25442 5110 25448 5162
rect 25500 5150 25506 5162
rect 25581 5153 25639 5159
rect 25581 5150 25593 5153
rect 25500 5122 25593 5150
rect 25500 5110 25506 5122
rect 25581 5119 25593 5122
rect 25627 5119 25639 5153
rect 25581 5113 25639 5119
rect 26546 5110 26552 5162
rect 26604 5150 26610 5162
rect 26777 5153 26835 5159
rect 26777 5150 26789 5153
rect 26604 5122 26789 5150
rect 26604 5110 26610 5122
rect 26777 5119 26789 5122
rect 26823 5119 26835 5153
rect 26777 5113 26835 5119
rect 27650 5110 27656 5162
rect 27708 5159 27714 5162
rect 27708 5153 27742 5159
rect 27730 5119 27742 5153
rect 27708 5113 27742 5119
rect 27708 5110 27714 5113
rect 28754 5110 28760 5162
rect 28812 5110 28818 5162
rect 29858 5110 29864 5162
rect 29916 5150 29922 5162
rect 29997 5153 30055 5159
rect 29997 5150 30009 5153
rect 29916 5122 30009 5150
rect 29916 5110 29922 5122
rect 29997 5119 30009 5122
rect 30043 5119 30055 5153
rect 29997 5113 30055 5119
rect 31238 5104 31244 5156
rect 31296 5144 31302 5156
rect 31455 5147 31513 5153
rect 31455 5144 31467 5147
rect 31296 5116 31467 5144
rect 31296 5104 31302 5116
rect 31455 5113 31467 5116
rect 31501 5113 31513 5147
rect 31455 5107 31513 5113
rect 31882 5110 31888 5162
rect 31940 5150 31946 5162
rect 31977 5153 32035 5159
rect 31977 5150 31989 5153
rect 31940 5122 31989 5150
rect 31940 5110 31946 5122
rect 31977 5119 31989 5122
rect 32023 5119 32035 5153
rect 31977 5113 32035 5119
rect 15601 5079 15659 5085
rect 33170 5076 33176 5128
rect 33228 5116 33234 5128
rect 33495 5127 33553 5133
rect 33495 5124 33507 5127
rect 33280 5116 33507 5124
rect 33228 5096 33507 5116
rect 33228 5088 33308 5096
rect 33495 5093 33507 5096
rect 33541 5093 33553 5127
rect 33228 5076 33234 5088
rect 33495 5087 33553 5093
rect 34458 5084 34464 5136
rect 34516 5124 34522 5136
rect 34691 5127 34749 5133
rect 34691 5124 34703 5127
rect 34516 5096 34703 5124
rect 34516 5084 34522 5096
rect 34691 5093 34703 5096
rect 34737 5093 34749 5127
rect 35102 5110 35108 5162
rect 35160 5150 35166 5162
rect 35197 5153 35255 5159
rect 35197 5150 35209 5153
rect 35160 5122 35209 5150
rect 35160 5110 35166 5122
rect 35197 5119 35209 5122
rect 35243 5119 35255 5153
rect 35197 5113 35255 5119
rect 36390 5110 36396 5162
rect 36448 5150 36454 5162
rect 36485 5153 36543 5159
rect 36485 5150 36497 5153
rect 36448 5122 36497 5150
rect 36448 5110 36454 5122
rect 36485 5119 36497 5122
rect 36531 5119 36543 5153
rect 36485 5113 36543 5119
rect 37678 5104 37684 5156
rect 37736 5144 37742 5156
rect 37895 5147 37953 5153
rect 37895 5144 37907 5147
rect 37736 5116 37907 5144
rect 37736 5104 37742 5116
rect 37895 5113 37907 5116
rect 37941 5113 37953 5147
rect 37895 5107 37953 5113
rect 38966 5104 38972 5156
rect 39024 5144 39030 5156
rect 39183 5147 39241 5153
rect 39183 5144 39195 5147
rect 39024 5116 39195 5144
rect 39024 5104 39030 5116
rect 39183 5113 39195 5116
rect 39229 5113 39241 5147
rect 39183 5107 39241 5113
rect 39610 5110 39616 5162
rect 39668 5150 39674 5162
rect 39705 5153 39763 5159
rect 39705 5150 39717 5153
rect 39668 5122 39717 5150
rect 39668 5110 39674 5122
rect 39705 5119 39717 5122
rect 39751 5119 39763 5153
rect 44118 5144 44124 5196
rect 44176 5184 44182 5196
rect 44213 5187 44271 5193
rect 44213 5184 44225 5187
rect 44176 5156 44225 5184
rect 44176 5144 44182 5156
rect 44213 5153 44225 5156
rect 44259 5153 44271 5187
rect 44213 5147 44271 5153
rect 45406 5144 45412 5196
rect 45464 5184 45470 5196
rect 46237 5187 46295 5193
rect 46237 5184 46249 5187
rect 45464 5156 46249 5184
rect 45464 5144 45470 5156
rect 46237 5153 46249 5156
rect 46283 5153 46295 5187
rect 46237 5147 46295 5153
rect 39705 5113 39763 5119
rect 34691 5087 34749 5093
rect 40898 5076 40904 5128
rect 40956 5116 40962 5128
rect 41223 5127 41281 5133
rect 41223 5124 41235 5127
rect 41008 5116 41235 5124
rect 40956 5096 41235 5116
rect 40956 5088 41036 5096
rect 41223 5093 41235 5096
rect 41269 5093 41281 5127
rect 40956 5076 40962 5088
rect 41223 5087 41281 5093
rect 42186 5076 42192 5128
rect 42244 5116 42250 5128
rect 42465 5119 42523 5125
rect 42465 5116 42477 5119
rect 42244 5088 42477 5116
rect 42244 5076 42250 5088
rect 42465 5085 42477 5088
rect 42511 5085 42523 5119
rect 42465 5079 42523 5085
rect 42830 5076 42836 5128
rect 42888 5116 42894 5128
rect 42945 5119 43003 5125
rect 42945 5116 42957 5119
rect 42888 5088 42957 5116
rect 42888 5076 42894 5088
rect 42945 5085 42957 5088
rect 42991 5085 43003 5119
rect 52582 5110 52588 5162
rect 52640 5110 52646 5162
rect 53686 5110 53692 5162
rect 53744 5150 53750 5162
rect 54790 5159 54796 5162
rect 53917 5153 53975 5159
rect 53917 5150 53929 5153
rect 53744 5122 53929 5150
rect 53744 5110 53750 5122
rect 53917 5119 53929 5122
rect 53963 5119 53975 5153
rect 53917 5113 53975 5119
rect 54769 5153 54796 5159
rect 54769 5119 54781 5153
rect 54769 5113 54796 5119
rect 54790 5110 54796 5113
rect 54848 5110 54854 5162
rect 55802 5110 55808 5162
rect 55860 5110 55866 5162
rect 57090 5110 57096 5162
rect 57148 5110 57154 5162
rect 58194 5110 58200 5162
rect 58252 5150 58258 5162
rect 58333 5153 58391 5159
rect 58333 5150 58345 5153
rect 58252 5122 58345 5150
rect 58252 5110 58258 5122
rect 58333 5119 58345 5122
rect 58379 5119 58391 5153
rect 58333 5113 58391 5119
rect 59114 5110 59120 5162
rect 59172 5110 59178 5162
rect 60310 5110 60316 5162
rect 60368 5110 60374 5162
rect 61414 5110 61420 5162
rect 61472 5150 61478 5162
rect 62518 5159 62524 5162
rect 61645 5153 61703 5159
rect 61645 5150 61657 5153
rect 61472 5122 61657 5150
rect 61472 5110 61478 5122
rect 61645 5119 61657 5122
rect 61691 5119 61703 5153
rect 61645 5113 61703 5119
rect 62497 5153 62524 5159
rect 62497 5119 62509 5153
rect 62497 5113 62524 5119
rect 62518 5110 62524 5113
rect 62576 5110 62582 5162
rect 63530 5110 63536 5162
rect 63588 5110 63594 5162
rect 64726 5110 64732 5162
rect 64784 5150 64790 5162
rect 64821 5153 64879 5159
rect 64821 5150 64833 5153
rect 64784 5122 64833 5150
rect 64784 5110 64790 5122
rect 64821 5119 64833 5122
rect 64867 5119 64879 5153
rect 64821 5113 64879 5119
rect 65830 5110 65836 5162
rect 65888 5150 65894 5162
rect 66061 5153 66119 5159
rect 66061 5150 66073 5153
rect 65888 5122 66073 5150
rect 65888 5110 65894 5122
rect 66061 5119 66073 5122
rect 66107 5119 66119 5153
rect 66061 5113 66119 5119
rect 66842 5110 66848 5162
rect 66900 5110 66906 5162
rect 42945 5079 43003 5085
rect 67946 5084 67952 5136
rect 68004 5124 68010 5136
rect 68179 5127 68237 5133
rect 68179 5124 68191 5127
rect 68004 5096 68191 5124
rect 68004 5084 68010 5096
rect 68179 5093 68191 5096
rect 68225 5093 68237 5127
rect 68179 5087 68237 5093
rect 69234 5076 69240 5128
rect 69292 5116 69298 5128
rect 69559 5127 69617 5133
rect 69559 5124 69571 5127
rect 69344 5116 69571 5124
rect 69292 5096 69571 5116
rect 69292 5088 69372 5096
rect 69559 5093 69571 5096
rect 69605 5093 69617 5127
rect 69878 5110 69884 5162
rect 69936 5150 69942 5162
rect 69973 5153 70031 5159
rect 69973 5150 69985 5153
rect 69936 5122 69985 5150
rect 69936 5110 69942 5122
rect 69973 5119 69985 5122
rect 70019 5119 70031 5153
rect 69973 5113 70031 5119
rect 71166 5110 71172 5162
rect 71224 5150 71230 5162
rect 71261 5153 71319 5159
rect 71261 5150 71273 5153
rect 71224 5122 71273 5150
rect 71224 5110 71230 5122
rect 71261 5119 71273 5122
rect 71307 5119 71319 5153
rect 71261 5113 71319 5119
rect 72454 5104 72460 5156
rect 72512 5144 72518 5156
rect 72671 5147 72729 5153
rect 72671 5144 72683 5147
rect 72512 5116 72683 5144
rect 72512 5104 72518 5116
rect 72671 5113 72683 5116
rect 72717 5113 72729 5147
rect 72671 5107 72729 5113
rect 73742 5104 73748 5156
rect 73800 5144 73806 5156
rect 73959 5147 74017 5153
rect 73959 5144 73971 5147
rect 73800 5116 73971 5144
rect 73800 5104 73806 5116
rect 73959 5113 73971 5116
rect 74005 5113 74017 5147
rect 73959 5107 74017 5113
rect 74386 5110 74392 5162
rect 74444 5150 74450 5162
rect 74527 5153 74585 5159
rect 74527 5150 74539 5153
rect 74444 5122 74539 5150
rect 74444 5110 74450 5122
rect 74527 5119 74539 5122
rect 74573 5119 74585 5153
rect 74527 5113 74585 5119
rect 69292 5076 69298 5088
rect 69559 5087 69617 5093
rect 75674 5084 75680 5136
rect 75732 5124 75738 5136
rect 75907 5127 75965 5133
rect 75907 5124 75919 5127
rect 75732 5096 75919 5124
rect 75732 5084 75738 5096
rect 75907 5093 75919 5096
rect 75953 5093 75965 5127
rect 75907 5087 75965 5093
rect 76962 5076 76968 5128
rect 77020 5116 77026 5128
rect 77287 5127 77345 5133
rect 77287 5124 77299 5127
rect 77072 5116 77299 5124
rect 77020 5096 77299 5116
rect 77020 5088 77100 5096
rect 77287 5093 77299 5096
rect 77333 5093 77345 5127
rect 77606 5110 77612 5162
rect 77664 5150 77670 5162
rect 77701 5153 77759 5159
rect 77701 5150 77713 5153
rect 77664 5122 77713 5150
rect 77664 5110 77670 5122
rect 77701 5119 77713 5122
rect 77747 5119 77759 5153
rect 81470 5144 81476 5196
rect 81528 5184 81534 5196
rect 82301 5187 82359 5193
rect 82301 5184 82313 5187
rect 81528 5156 82313 5184
rect 81528 5144 81534 5156
rect 82301 5153 82313 5156
rect 82347 5153 82359 5187
rect 82301 5147 82359 5153
rect 77701 5113 77759 5119
rect 77020 5076 77026 5088
rect 77287 5087 77345 5093
rect 78894 5076 78900 5128
rect 78952 5116 78958 5128
rect 79009 5119 79067 5125
rect 79009 5116 79021 5119
rect 78952 5088 79021 5116
rect 78952 5076 78958 5088
rect 79009 5085 79021 5088
rect 79055 5085 79067 5119
rect 79009 5079 79067 5085
rect 80182 5076 80188 5128
rect 80240 5116 80246 5128
rect 80461 5119 80519 5125
rect 80461 5116 80473 5119
rect 80240 5088 80473 5116
rect 80240 5076 80246 5088
rect 80461 5085 80473 5088
rect 80507 5085 80519 5119
rect 80461 5079 80519 5085
rect 15782 5008 15788 5060
rect 15840 5048 15846 5060
rect 16032 5051 16090 5057
rect 16032 5048 16044 5051
rect 15840 5020 16044 5048
rect 15840 5008 15846 5020
rect 16032 5017 16044 5020
rect 16078 5017 16090 5051
rect 16032 5011 16090 5017
rect 16426 5008 16432 5060
rect 16484 5048 16490 5060
rect 16567 5051 16625 5057
rect 16567 5048 16579 5051
rect 16484 5020 16579 5048
rect 16484 5008 16490 5020
rect 16567 5017 16579 5020
rect 16613 5017 16625 5051
rect 16567 5011 16625 5017
rect 17714 5008 17720 5060
rect 17772 5048 17778 5060
rect 18056 5051 18114 5057
rect 18056 5048 18068 5051
rect 17772 5020 18068 5048
rect 17772 5008 17778 5020
rect 18056 5017 18068 5020
rect 18102 5017 18114 5051
rect 18056 5011 18114 5017
rect 19002 5008 19008 5060
rect 19060 5048 19066 5060
rect 19252 5051 19310 5057
rect 19252 5048 19264 5051
rect 19060 5020 19264 5048
rect 19060 5008 19066 5020
rect 19252 5017 19264 5020
rect 19298 5017 19310 5051
rect 19252 5011 19310 5017
rect 19738 5008 19744 5060
rect 19796 5057 19802 5060
rect 19796 5051 19845 5057
rect 19796 5017 19799 5051
rect 19833 5017 19845 5051
rect 19796 5011 19845 5017
rect 19796 5008 19802 5011
rect 20934 5008 20940 5060
rect 20992 5048 20998 5060
rect 21184 5051 21242 5057
rect 21184 5048 21196 5051
rect 20992 5020 21196 5048
rect 20992 5008 20998 5020
rect 21184 5017 21196 5020
rect 21230 5017 21242 5051
rect 21184 5011 21242 5017
rect 22222 5008 22228 5060
rect 22280 5048 22286 5060
rect 22472 5051 22530 5057
rect 22472 5048 22484 5051
rect 22280 5020 22484 5048
rect 22280 5008 22286 5020
rect 22472 5017 22484 5020
rect 22518 5017 22530 5051
rect 22472 5011 22530 5017
rect 23510 5008 23516 5060
rect 23568 5048 23574 5060
rect 23760 5051 23818 5057
rect 23760 5048 23772 5051
rect 23568 5020 23772 5048
rect 23568 5008 23574 5020
rect 23760 5017 23772 5020
rect 23806 5017 23818 5051
rect 23760 5011 23818 5017
rect 24154 5008 24160 5060
rect 24212 5048 24218 5060
rect 24295 5051 24353 5057
rect 24295 5048 24307 5051
rect 24212 5020 24307 5048
rect 24212 5008 24218 5020
rect 24295 5017 24307 5020
rect 24341 5017 24353 5051
rect 24295 5011 24353 5017
rect 25442 5008 25448 5060
rect 25500 5048 25506 5060
rect 25784 5051 25842 5057
rect 25784 5048 25796 5051
rect 25500 5020 25796 5048
rect 25500 5008 25506 5020
rect 25784 5017 25796 5020
rect 25830 5017 25842 5051
rect 25784 5011 25842 5017
rect 26730 5008 26736 5060
rect 26788 5048 26794 5060
rect 26980 5051 27038 5057
rect 26980 5048 26992 5051
rect 26788 5020 26992 5048
rect 26788 5008 26794 5020
rect 26980 5017 26992 5020
rect 27026 5017 27038 5051
rect 26980 5011 27038 5017
rect 27374 5008 27380 5060
rect 27432 5048 27438 5060
rect 27515 5051 27573 5057
rect 27515 5048 27527 5051
rect 27432 5020 27527 5048
rect 27432 5008 27438 5020
rect 27515 5017 27527 5020
rect 27561 5017 27573 5051
rect 27515 5011 27573 5017
rect 28662 5008 28668 5060
rect 28720 5048 28726 5060
rect 28912 5051 28970 5057
rect 28912 5048 28924 5051
rect 28720 5020 28924 5048
rect 28720 5008 28726 5020
rect 28912 5017 28924 5020
rect 28958 5017 28970 5051
rect 28912 5011 28970 5017
rect 29950 5008 29956 5060
rect 30008 5048 30014 5060
rect 30200 5051 30258 5057
rect 30200 5048 30212 5051
rect 30008 5020 30212 5048
rect 30008 5008 30014 5020
rect 30200 5017 30212 5020
rect 30246 5017 30258 5051
rect 30200 5011 30258 5017
rect 52490 5008 52496 5060
rect 52548 5048 52554 5060
rect 52740 5051 52798 5057
rect 52740 5048 52752 5051
rect 52548 5020 52752 5048
rect 52548 5008 52554 5020
rect 52740 5017 52752 5020
rect 52786 5017 52798 5051
rect 52740 5011 52798 5017
rect 53778 5008 53784 5060
rect 53836 5048 53842 5060
rect 54120 5051 54178 5057
rect 54120 5048 54132 5051
rect 53836 5020 54132 5048
rect 53836 5008 53842 5020
rect 54120 5017 54132 5020
rect 54166 5017 54178 5051
rect 54120 5011 54178 5017
rect 54422 5008 54428 5060
rect 54480 5048 54486 5060
rect 54563 5051 54621 5057
rect 54563 5048 54575 5051
rect 54480 5020 54575 5048
rect 54480 5008 54486 5020
rect 54563 5017 54575 5020
rect 54609 5017 54621 5051
rect 54563 5011 54621 5017
rect 55710 5008 55716 5060
rect 55768 5048 55774 5060
rect 55960 5051 56018 5057
rect 55960 5048 55972 5051
rect 55768 5020 55972 5048
rect 55768 5008 55774 5020
rect 55960 5017 55972 5020
rect 56006 5017 56018 5051
rect 55960 5011 56018 5017
rect 56998 5008 57004 5060
rect 57056 5048 57062 5060
rect 57248 5051 57306 5057
rect 57248 5048 57260 5051
rect 57056 5020 57260 5048
rect 57056 5008 57062 5020
rect 57248 5017 57260 5020
rect 57294 5017 57306 5051
rect 57248 5011 57306 5017
rect 58286 5008 58292 5060
rect 58344 5048 58350 5060
rect 58536 5051 58594 5057
rect 58536 5048 58548 5051
rect 58344 5020 58548 5048
rect 58344 5008 58350 5020
rect 58536 5017 58548 5020
rect 58582 5017 58594 5051
rect 58536 5011 58594 5017
rect 58930 5008 58936 5060
rect 58988 5048 58994 5060
rect 59272 5051 59330 5057
rect 59272 5048 59284 5051
rect 58988 5020 59284 5048
rect 58988 5008 58994 5020
rect 59272 5017 59284 5020
rect 59318 5017 59330 5051
rect 59272 5011 59330 5017
rect 60218 5008 60224 5060
rect 60276 5048 60282 5060
rect 60468 5051 60526 5057
rect 60468 5048 60480 5051
rect 60276 5020 60480 5048
rect 60276 5008 60282 5020
rect 60468 5017 60480 5020
rect 60514 5017 60526 5051
rect 60468 5011 60526 5017
rect 61506 5008 61512 5060
rect 61564 5048 61570 5060
rect 61848 5051 61906 5057
rect 61848 5048 61860 5051
rect 61564 5020 61860 5048
rect 61564 5008 61570 5020
rect 61848 5017 61860 5020
rect 61894 5017 61906 5051
rect 61848 5011 61906 5017
rect 62150 5008 62156 5060
rect 62208 5048 62214 5060
rect 62291 5051 62349 5057
rect 62291 5048 62303 5051
rect 62208 5020 62303 5048
rect 62208 5008 62214 5020
rect 62291 5017 62303 5020
rect 62337 5017 62349 5051
rect 62291 5011 62349 5017
rect 63438 5008 63444 5060
rect 63496 5048 63502 5060
rect 63688 5051 63746 5057
rect 63688 5048 63700 5051
rect 63496 5020 63700 5048
rect 63496 5008 63502 5020
rect 63688 5017 63700 5020
rect 63734 5017 63746 5051
rect 63688 5011 63746 5017
rect 64726 5008 64732 5060
rect 64784 5048 64790 5060
rect 64976 5051 65034 5057
rect 64976 5048 64988 5051
rect 64784 5020 64988 5048
rect 64784 5008 64790 5020
rect 64976 5017 64988 5020
rect 65022 5017 65034 5051
rect 64976 5011 65034 5017
rect 66014 5008 66020 5060
rect 66072 5048 66078 5060
rect 66264 5051 66322 5057
rect 66264 5048 66276 5051
rect 66072 5020 66276 5048
rect 66072 5008 66078 5020
rect 66264 5017 66276 5020
rect 66310 5017 66322 5051
rect 66264 5011 66322 5017
rect 66658 5008 66664 5060
rect 66716 5048 66722 5060
rect 67000 5051 67058 5057
rect 67000 5048 67012 5051
rect 66716 5020 67012 5048
rect 66716 5008 66722 5020
rect 67000 5017 67012 5020
rect 67046 5017 67058 5051
rect 67000 5011 67058 5017
rect 4876 4922 88964 4944
rect 4876 4870 19382 4922
rect 19434 4870 19446 4922
rect 19498 4870 19510 4922
rect 19562 4870 19574 4922
rect 19626 4870 19638 4922
rect 19690 4870 38382 4922
rect 38434 4870 38446 4922
rect 38498 4870 38510 4922
rect 38562 4870 38574 4922
rect 38626 4870 38638 4922
rect 38690 4870 57382 4922
rect 57434 4870 57446 4922
rect 57498 4870 57510 4922
rect 57562 4870 57574 4922
rect 57626 4870 57638 4922
rect 57690 4870 76382 4922
rect 76434 4870 76446 4922
rect 76498 4870 76510 4922
rect 76562 4870 76574 4922
rect 76626 4870 76638 4922
rect 76690 4870 88964 4922
rect 4876 4848 88964 4870
<< via1 >>
rect 18722 89190 18774 89242
rect 18786 89190 18838 89242
rect 18850 89190 18902 89242
rect 18914 89190 18966 89242
rect 18978 89190 19030 89242
rect 37722 89190 37774 89242
rect 37786 89190 37838 89242
rect 37850 89190 37902 89242
rect 37914 89190 37966 89242
rect 37978 89190 38030 89242
rect 56722 89190 56774 89242
rect 56786 89190 56838 89242
rect 56850 89190 56902 89242
rect 56914 89190 56966 89242
rect 56978 89190 57030 89242
rect 75722 89190 75774 89242
rect 75786 89190 75838 89242
rect 75850 89190 75902 89242
rect 75914 89190 75966 89242
rect 75978 89190 76030 89242
rect 31244 89056 31296 89108
rect 31888 89056 31940 89108
rect 33176 89056 33228 89108
rect 34464 89056 34516 89108
rect 35108 89056 35160 89108
rect 36396 89056 36448 89108
rect 37592 89056 37644 89108
rect 38972 89056 39024 89108
rect 39616 89056 39668 89108
rect 40904 89056 40956 89108
rect 42192 89056 42244 89108
rect 42836 89056 42888 89108
rect 44124 89056 44176 89108
rect 45412 89056 45464 89108
rect 46700 89056 46752 89108
rect 56360 89056 56412 89108
rect 57648 89056 57700 89108
rect 67952 89056 68004 89108
rect 69240 89056 69292 89108
rect 69884 89056 69936 89108
rect 71172 89056 71224 89108
rect 72460 89056 72512 89108
rect 73748 89056 73800 89108
rect 74392 89056 74444 89108
rect 75588 89056 75640 89108
rect 76968 89056 77020 89108
rect 77612 89056 77664 89108
rect 78900 89056 78952 89108
rect 80188 89056 80240 89108
rect 81476 89056 81528 89108
rect 82120 89056 82172 89108
rect 15788 88886 15840 88938
rect 16432 88886 16484 88938
rect 17720 88852 17772 88904
rect 19100 88929 19152 88938
rect 19100 88895 19109 88929
rect 19109 88895 19143 88929
rect 19143 88895 19152 88929
rect 19100 88886 19152 88895
rect 19652 88886 19704 88938
rect 20940 88852 20992 88904
rect 22228 88886 22280 88938
rect 23516 88886 23568 88938
rect 24160 88886 24212 88938
rect 25448 88920 25500 88972
rect 24344 88852 24396 88904
rect 26736 88852 26788 88904
rect 27380 88852 27432 88904
rect 28668 88886 28720 88938
rect 29956 88886 30008 88938
rect 30968 88852 31020 88904
rect 32072 88886 32124 88938
rect 33176 88886 33228 88938
rect 34280 88886 34332 88938
rect 35384 88929 35436 88938
rect 35384 88895 35424 88929
rect 35424 88895 35436 88929
rect 35384 88886 35436 88895
rect 36488 88929 36540 88938
rect 36488 88895 36497 88929
rect 36497 88895 36531 88929
rect 36531 88895 36540 88929
rect 36488 88886 36540 88895
rect 37592 88886 37644 88938
rect 38788 88886 38840 88938
rect 39800 88886 39852 88938
rect 40904 88886 40956 88938
rect 42008 88886 42060 88938
rect 43112 88929 43164 88938
rect 43112 88895 43152 88929
rect 43152 88895 43164 88929
rect 43112 88886 43164 88895
rect 44216 88929 44268 88938
rect 44216 88895 44225 88929
rect 44225 88895 44259 88929
rect 44259 88895 44268 88929
rect 44216 88886 44268 88895
rect 45320 88886 45372 88938
rect 49920 88924 49972 88933
rect 49920 88890 49929 88924
rect 49929 88890 49963 88924
rect 49963 88890 49972 88924
rect 49920 88881 49972 88890
rect 50012 88852 50064 88904
rect 52496 88886 52548 88938
rect 53784 88886 53836 88938
rect 54428 88852 54480 88904
rect 55716 88886 55768 88938
rect 57096 88929 57148 88938
rect 57096 88895 57105 88929
rect 57105 88895 57139 88929
rect 57139 88895 57148 88929
rect 57096 88886 57148 88895
rect 58292 88852 58344 88904
rect 58936 88886 58988 88938
rect 60224 88886 60276 88938
rect 61512 88886 61564 88938
rect 62156 88920 62208 88972
rect 15512 88784 15564 88836
rect 16708 88827 16760 88836
rect 16708 88793 16731 88827
rect 16731 88793 16760 88827
rect 16708 88784 16760 88793
rect 17812 88784 17864 88836
rect 18640 88784 18692 88836
rect 19928 88827 19980 88836
rect 19928 88793 19951 88827
rect 19951 88793 19980 88827
rect 19928 88784 19980 88793
rect 21032 88784 21084 88836
rect 22136 88784 22188 88836
rect 23240 88784 23292 88836
rect 25448 88784 25500 88836
rect 26552 88784 26604 88836
rect 27656 88784 27708 88836
rect 28760 88784 28812 88836
rect 29864 88784 29916 88836
rect 52772 88827 52824 88836
rect 52772 88793 52795 88827
rect 52795 88793 52824 88827
rect 52772 88784 52824 88793
rect 54152 88827 54204 88836
rect 54152 88793 54175 88827
rect 54175 88793 54204 88827
rect 54152 88784 54204 88793
rect 54796 88784 54848 88836
rect 55992 88827 56044 88836
rect 55992 88793 56015 88827
rect 56015 88793 56044 88827
rect 55992 88784 56044 88793
rect 57096 88784 57148 88836
rect 58384 88784 58436 88836
rect 59304 88827 59356 88836
rect 59304 88793 59327 88827
rect 59327 88793 59356 88827
rect 59304 88784 59356 88793
rect 60316 88784 60368 88836
rect 61420 88784 61472 88836
rect 63444 88852 63496 88904
rect 64732 88852 64784 88904
rect 66020 88886 66072 88938
rect 66664 88886 66716 88938
rect 68044 88929 68096 88938
rect 68044 88895 68053 88929
rect 68053 88895 68087 88929
rect 68087 88895 68096 88929
rect 68044 88886 68096 88895
rect 69424 88929 69476 88938
rect 69424 88895 69433 88929
rect 69433 88895 69467 88929
rect 69467 88895 69476 88929
rect 69424 88886 69476 88895
rect 70252 88929 70304 88938
rect 70252 88895 70271 88929
rect 70271 88895 70304 88929
rect 70252 88886 70304 88895
rect 71356 88886 71408 88938
rect 72460 88886 72512 88938
rect 73564 88886 73616 88938
rect 74668 88886 74720 88938
rect 75496 88886 75548 88938
rect 76876 88886 76928 88938
rect 77980 88929 78032 88938
rect 77980 88895 77999 88929
rect 77999 88895 78032 88929
rect 77980 88886 78032 88895
rect 79084 88886 79136 88938
rect 80280 88929 80332 88938
rect 80280 88895 80289 88929
rect 80289 88895 80323 88929
rect 80323 88895 80332 88929
rect 80280 88886 80332 88895
rect 81292 88886 81344 88938
rect 82396 88886 82448 88938
rect 62524 88784 62576 88836
rect 63720 88784 63772 88836
rect 65100 88784 65152 88836
rect 65836 88784 65888 88836
rect 66940 88784 66992 88836
rect 19382 88646 19434 88698
rect 19446 88646 19498 88698
rect 19510 88646 19562 88698
rect 19574 88646 19626 88698
rect 19638 88646 19690 88698
rect 38382 88646 38434 88698
rect 38446 88646 38498 88698
rect 38510 88646 38562 88698
rect 38574 88646 38626 88698
rect 38638 88646 38690 88698
rect 57382 88646 57434 88698
rect 57446 88646 57498 88698
rect 57510 88646 57562 88698
rect 57574 88646 57626 88698
rect 57638 88646 57690 88698
rect 76382 88646 76434 88698
rect 76446 88646 76498 88698
rect 76510 88646 76562 88698
rect 76574 88646 76626 88698
rect 76638 88646 76690 88698
rect 48632 88410 48684 88462
rect 49644 88419 49696 88428
rect 49644 88385 49653 88419
rect 49653 88385 49687 88419
rect 49687 88385 49696 88419
rect 49644 88376 49696 88385
rect 18722 88102 18774 88154
rect 18786 88102 18838 88154
rect 18850 88102 18902 88154
rect 18914 88102 18966 88154
rect 18978 88102 19030 88154
rect 37722 88102 37774 88154
rect 37786 88102 37838 88154
rect 37850 88102 37902 88154
rect 37914 88102 37966 88154
rect 37978 88102 38030 88154
rect 56722 88102 56774 88154
rect 56786 88102 56838 88154
rect 56850 88102 56902 88154
rect 56914 88102 56966 88154
rect 56978 88102 57030 88154
rect 75722 88102 75774 88154
rect 75786 88102 75838 88154
rect 75850 88102 75902 88154
rect 75914 88102 75966 88154
rect 75978 88102 76030 88154
rect 19382 87558 19434 87610
rect 19446 87558 19498 87610
rect 19510 87558 19562 87610
rect 19574 87558 19626 87610
rect 19638 87558 19690 87610
rect 38382 87558 38434 87610
rect 38446 87558 38498 87610
rect 38510 87558 38562 87610
rect 38574 87558 38626 87610
rect 38638 87558 38690 87610
rect 57382 87558 57434 87610
rect 57446 87558 57498 87610
rect 57510 87558 57562 87610
rect 57574 87558 57626 87610
rect 57638 87558 57690 87610
rect 76382 87558 76434 87610
rect 76446 87558 76498 87610
rect 76510 87558 76562 87610
rect 76574 87558 76626 87610
rect 76638 87558 76690 87610
rect 49276 87322 49328 87374
rect 49644 87322 49696 87374
rect 83684 87288 83736 87340
rect 5954 87014 6006 87066
rect 6018 87014 6070 87066
rect 6082 87014 6134 87066
rect 6146 87014 6198 87066
rect 6210 87014 6262 87066
rect 18722 87014 18774 87066
rect 18786 87014 18838 87066
rect 18850 87014 18902 87066
rect 18914 87014 18966 87066
rect 18978 87014 19030 87066
rect 37722 87014 37774 87066
rect 37786 87014 37838 87066
rect 37850 87014 37902 87066
rect 37914 87014 37966 87066
rect 37978 87014 38030 87066
rect 56722 87014 56774 87066
rect 56786 87014 56838 87066
rect 56850 87014 56902 87066
rect 56914 87014 56966 87066
rect 56978 87014 57030 87066
rect 75722 87014 75774 87066
rect 75786 87014 75838 87066
rect 75850 87014 75902 87066
rect 75914 87014 75966 87066
rect 75978 87014 76030 87066
rect 87098 87014 87150 87066
rect 87162 87014 87214 87066
rect 87226 87014 87278 87066
rect 87290 87014 87342 87066
rect 87354 87014 87406 87066
rect 7600 86676 7652 86728
rect 47988 86676 48040 86728
rect 50012 86748 50064 86757
rect 50012 86714 50021 86748
rect 50021 86714 50055 86748
rect 50055 86714 50064 86748
rect 50012 86705 50064 86714
rect 84052 86676 84104 86728
rect 31704 86651 31756 86660
rect 31704 86617 31713 86651
rect 31713 86617 31747 86651
rect 31747 86617 31756 86651
rect 31704 86608 31756 86617
rect 6690 86470 6742 86522
rect 6754 86470 6806 86522
rect 6818 86470 6870 86522
rect 6882 86470 6934 86522
rect 6946 86470 6998 86522
rect 19382 86470 19434 86522
rect 19446 86470 19498 86522
rect 19510 86470 19562 86522
rect 19574 86470 19626 86522
rect 19638 86470 19690 86522
rect 38382 86470 38434 86522
rect 38446 86470 38498 86522
rect 38510 86470 38562 86522
rect 38574 86470 38626 86522
rect 38638 86470 38690 86522
rect 57382 86470 57434 86522
rect 57446 86470 57498 86522
rect 57510 86470 57562 86522
rect 57574 86470 57626 86522
rect 57638 86470 57690 86522
rect 76382 86470 76434 86522
rect 76446 86470 76498 86522
rect 76510 86470 76562 86522
rect 76574 86470 76626 86522
rect 76638 86470 76690 86522
rect 87834 86470 87886 86522
rect 87898 86470 87950 86522
rect 87962 86470 88014 86522
rect 88026 86470 88078 86522
rect 88090 86470 88142 86522
rect 5954 85926 6006 85978
rect 6018 85926 6070 85978
rect 6082 85926 6134 85978
rect 6146 85926 6198 85978
rect 6210 85926 6262 85978
rect 87098 85926 87150 85978
rect 87162 85926 87214 85978
rect 87226 85926 87278 85978
rect 87290 85926 87342 85978
rect 87354 85926 87406 85978
rect 6690 85382 6742 85434
rect 6754 85382 6806 85434
rect 6818 85382 6870 85434
rect 6882 85382 6934 85434
rect 6946 85382 6998 85434
rect 87834 85382 87886 85434
rect 87898 85382 87950 85434
rect 87962 85382 88014 85434
rect 88026 85382 88078 85434
rect 88090 85382 88142 85434
rect 5954 84838 6006 84890
rect 6018 84838 6070 84890
rect 6082 84838 6134 84890
rect 6146 84838 6198 84890
rect 6210 84838 6262 84890
rect 87098 84838 87150 84890
rect 87162 84838 87214 84890
rect 87226 84838 87278 84890
rect 87290 84838 87342 84890
rect 87354 84838 87406 84890
rect 6690 84294 6742 84346
rect 6754 84294 6806 84346
rect 6818 84294 6870 84346
rect 6882 84294 6934 84346
rect 6946 84294 6998 84346
rect 87834 84294 87886 84346
rect 87898 84294 87950 84346
rect 87962 84294 88014 84346
rect 88026 84294 88078 84346
rect 88090 84294 88142 84346
rect 13672 84228 13724 84280
rect 50012 84228 50064 84280
rect 12568 84160 12620 84212
rect 48908 84160 48960 84212
rect 11280 84092 11332 84144
rect 31704 84092 31756 84144
rect 47804 84092 47856 84144
rect 5954 83750 6006 83802
rect 6018 83750 6070 83802
rect 6082 83750 6134 83802
rect 6146 83750 6198 83802
rect 6210 83750 6262 83802
rect 87098 83750 87150 83802
rect 87162 83750 87214 83802
rect 87226 83750 87278 83802
rect 87290 83750 87342 83802
rect 87354 83750 87406 83802
rect 6690 83206 6742 83258
rect 6754 83206 6806 83258
rect 6818 83206 6870 83258
rect 6882 83206 6934 83258
rect 6946 83206 6998 83258
rect 87834 83206 87886 83258
rect 87898 83206 87950 83258
rect 87962 83206 88014 83258
rect 88026 83206 88078 83258
rect 88090 83206 88142 83258
rect 5954 82662 6006 82714
rect 6018 82662 6070 82714
rect 6082 82662 6134 82714
rect 6146 82662 6198 82714
rect 6210 82662 6262 82714
rect 87098 82662 87150 82714
rect 87162 82662 87214 82714
rect 87226 82662 87278 82714
rect 87290 82662 87342 82714
rect 87354 82662 87406 82714
rect 6690 82118 6742 82170
rect 6754 82118 6806 82170
rect 6818 82118 6870 82170
rect 6882 82118 6934 82170
rect 6946 82118 6998 82170
rect 87834 82118 87886 82170
rect 87898 82118 87950 82170
rect 87962 82118 88014 82170
rect 88026 82118 88078 82170
rect 88090 82118 88142 82170
rect 5954 81574 6006 81626
rect 6018 81574 6070 81626
rect 6082 81574 6134 81626
rect 6146 81574 6198 81626
rect 6210 81574 6262 81626
rect 87098 81574 87150 81626
rect 87162 81574 87214 81626
rect 87226 81574 87278 81626
rect 87290 81574 87342 81626
rect 87354 81574 87406 81626
rect 6690 81030 6742 81082
rect 6754 81030 6806 81082
rect 6818 81030 6870 81082
rect 6882 81030 6934 81082
rect 6946 81030 6998 81082
rect 87834 81030 87886 81082
rect 87898 81030 87950 81082
rect 87962 81030 88014 81082
rect 88026 81030 88078 81082
rect 88090 81030 88142 81082
rect 7140 80760 7192 80812
rect 88652 80803 88704 80812
rect 88652 80769 88671 80803
rect 88671 80769 88704 80803
rect 88652 80760 88704 80769
rect 2908 80624 2960 80676
rect 84328 80624 84380 80676
rect 5954 80486 6006 80538
rect 6018 80486 6070 80538
rect 6082 80486 6134 80538
rect 6146 80486 6198 80538
rect 6210 80486 6262 80538
rect 87098 80486 87150 80538
rect 87162 80486 87214 80538
rect 87226 80486 87278 80538
rect 87290 80486 87342 80538
rect 87354 80486 87406 80538
rect 6690 79942 6742 79994
rect 6754 79942 6806 79994
rect 6818 79942 6870 79994
rect 6882 79942 6934 79994
rect 6946 79942 6998 79994
rect 87834 79942 87886 79994
rect 87898 79942 87950 79994
rect 87962 79942 88014 79994
rect 88026 79942 88078 79994
rect 88090 79942 88142 79994
rect 88652 79749 88704 79758
rect 7140 79672 7192 79724
rect 88652 79715 88671 79749
rect 88671 79715 88704 79749
rect 88652 79706 88704 79715
rect 2724 79536 2776 79588
rect 84328 79536 84380 79588
rect 5954 79398 6006 79450
rect 6018 79398 6070 79450
rect 6082 79398 6134 79450
rect 6146 79398 6198 79450
rect 6210 79398 6262 79450
rect 87098 79398 87150 79450
rect 87162 79398 87214 79450
rect 87226 79398 87278 79450
rect 87290 79398 87342 79450
rect 87354 79398 87406 79450
rect 6690 78854 6742 78906
rect 6754 78854 6806 78906
rect 6818 78854 6870 78906
rect 6882 78854 6934 78906
rect 6946 78854 6998 78906
rect 87834 78854 87886 78906
rect 87898 78854 87950 78906
rect 87962 78854 88014 78906
rect 88026 78854 88078 78906
rect 88090 78854 88142 78906
rect 88652 78661 88704 78670
rect 7140 78584 7192 78636
rect 88652 78627 88671 78661
rect 88671 78627 88704 78661
rect 88652 78618 88704 78627
rect 2908 78448 2960 78500
rect 84328 78448 84380 78500
rect 5954 78310 6006 78362
rect 6018 78310 6070 78362
rect 6082 78310 6134 78362
rect 6146 78310 6198 78362
rect 6210 78310 6262 78362
rect 87098 78310 87150 78362
rect 87162 78310 87214 78362
rect 87226 78310 87278 78362
rect 87290 78310 87342 78362
rect 87354 78310 87406 78362
rect 6690 77766 6742 77818
rect 6754 77766 6806 77818
rect 6818 77766 6870 77818
rect 6882 77766 6934 77818
rect 6946 77766 6998 77818
rect 87834 77766 87886 77818
rect 87898 77766 87950 77818
rect 87962 77766 88014 77818
rect 88026 77766 88078 77818
rect 88090 77766 88142 77818
rect 4380 77632 4432 77684
rect 5668 77530 5720 77582
rect 90032 77564 90084 77616
rect 84328 77428 84380 77480
rect 5954 77222 6006 77274
rect 6018 77222 6070 77274
rect 6082 77222 6134 77274
rect 6146 77222 6198 77274
rect 6210 77222 6262 77274
rect 87098 77222 87150 77274
rect 87162 77222 87214 77274
rect 87226 77222 87278 77274
rect 87290 77222 87342 77274
rect 87354 77222 87406 77274
rect 6690 76678 6742 76730
rect 6754 76678 6806 76730
rect 6818 76678 6870 76730
rect 6882 76678 6934 76730
rect 6946 76678 6998 76730
rect 87834 76678 87886 76730
rect 87898 76678 87950 76730
rect 87962 76678 88014 76730
rect 88026 76678 88078 76730
rect 88090 76678 88142 76730
rect 5954 76134 6006 76186
rect 6018 76134 6070 76186
rect 6082 76134 6134 76186
rect 6146 76134 6198 76186
rect 6210 76134 6262 76186
rect 87098 76134 87150 76186
rect 87162 76134 87214 76186
rect 87226 76134 87278 76186
rect 87290 76134 87342 76186
rect 87354 76134 87406 76186
rect 84328 75932 84380 75984
rect 7140 75864 7192 75916
rect 88744 75796 88796 75848
rect 2908 75728 2960 75780
rect 6690 75590 6742 75642
rect 6754 75590 6806 75642
rect 6818 75590 6870 75642
rect 6882 75590 6934 75642
rect 6946 75590 6998 75642
rect 87834 75590 87886 75642
rect 87898 75590 87950 75642
rect 87962 75590 88014 75642
rect 88026 75590 88078 75642
rect 88090 75590 88142 75642
rect 88560 75431 88612 75440
rect 88560 75397 88569 75431
rect 88569 75397 88603 75431
rect 88603 75397 88612 75431
rect 88560 75388 88612 75397
rect 7140 75320 7192 75372
rect 84328 75252 84380 75304
rect 2908 75184 2960 75236
rect 5954 75046 6006 75098
rect 6018 75046 6070 75098
rect 6082 75046 6134 75098
rect 6146 75046 6198 75098
rect 6210 75046 6262 75098
rect 87098 75046 87150 75098
rect 87162 75046 87214 75098
rect 87226 75046 87278 75098
rect 87290 75046 87342 75098
rect 87354 75046 87406 75098
rect 6690 74502 6742 74554
rect 6754 74502 6806 74554
rect 6818 74502 6870 74554
rect 6882 74502 6934 74554
rect 6946 74502 6998 74554
rect 87834 74502 87886 74554
rect 87898 74502 87950 74554
rect 87962 74502 88014 74554
rect 88026 74502 88078 74554
rect 88090 74502 88142 74554
rect 88560 74343 88612 74352
rect 88560 74309 88569 74343
rect 88569 74309 88603 74343
rect 88603 74309 88612 74343
rect 88560 74300 88612 74309
rect 7140 74232 7192 74284
rect 84328 74164 84380 74216
rect 2908 74096 2960 74148
rect 5954 73958 6006 74010
rect 6018 73958 6070 74010
rect 6082 73958 6134 74010
rect 6146 73958 6198 74010
rect 6210 73958 6262 74010
rect 87098 73958 87150 74010
rect 87162 73958 87214 74010
rect 87226 73958 87278 74010
rect 87290 73958 87342 74010
rect 87354 73958 87406 74010
rect 6690 73414 6742 73466
rect 6754 73414 6806 73466
rect 6818 73414 6870 73466
rect 6882 73414 6934 73466
rect 6946 73414 6998 73466
rect 87834 73414 87886 73466
rect 87898 73414 87950 73466
rect 87962 73414 88014 73466
rect 88026 73414 88078 73466
rect 88090 73414 88142 73466
rect 88652 73221 88704 73230
rect 7140 73144 7192 73196
rect 88652 73187 88667 73221
rect 88667 73187 88704 73221
rect 88652 73178 88704 73187
rect 2908 73008 2960 73060
rect 84328 73008 84380 73060
rect 5954 72870 6006 72922
rect 6018 72870 6070 72922
rect 6082 72870 6134 72922
rect 6146 72870 6198 72922
rect 6210 72870 6262 72922
rect 87098 72870 87150 72922
rect 87162 72870 87214 72922
rect 87226 72870 87278 72922
rect 87290 72870 87342 72922
rect 87354 72870 87406 72922
rect 6690 72326 6742 72378
rect 6754 72326 6806 72378
rect 6818 72326 6870 72378
rect 6882 72326 6934 72378
rect 6946 72326 6998 72378
rect 87834 72326 87886 72378
rect 87898 72326 87950 72378
rect 87962 72326 88014 72378
rect 88026 72326 88078 72378
rect 88090 72326 88142 72378
rect 5668 72090 5720 72142
rect 90124 72056 90176 72108
rect 4380 71988 4432 72040
rect 87180 71988 87232 72040
rect 5954 71782 6006 71834
rect 6018 71782 6070 71834
rect 6082 71782 6134 71834
rect 6146 71782 6198 71834
rect 6210 71782 6262 71834
rect 87098 71782 87150 71834
rect 87162 71782 87214 71834
rect 87226 71782 87278 71834
rect 87290 71782 87342 71834
rect 87354 71782 87406 71834
rect 6690 71238 6742 71290
rect 6754 71238 6806 71290
rect 6818 71238 6870 71290
rect 6882 71238 6934 71290
rect 6946 71238 6998 71290
rect 87834 71238 87886 71290
rect 87898 71238 87950 71290
rect 87962 71238 88014 71290
rect 88026 71238 88078 71290
rect 88090 71238 88142 71290
rect 5954 70694 6006 70746
rect 6018 70694 6070 70746
rect 6082 70694 6134 70746
rect 6146 70694 6198 70746
rect 6210 70694 6262 70746
rect 87098 70694 87150 70746
rect 87162 70694 87214 70746
rect 87226 70694 87278 70746
rect 87290 70694 87342 70746
rect 87354 70694 87406 70746
rect 84328 70492 84380 70544
rect 5668 70390 5720 70442
rect 89940 70356 89992 70408
rect 2908 70288 2960 70340
rect 6690 70150 6742 70202
rect 6754 70150 6806 70202
rect 6818 70150 6870 70202
rect 6882 70150 6934 70202
rect 6946 70150 6998 70202
rect 87834 70150 87886 70202
rect 87898 70150 87950 70202
rect 87962 70150 88014 70202
rect 88026 70150 88078 70202
rect 88090 70150 88142 70202
rect 88560 69991 88612 70000
rect 88560 69957 88569 69991
rect 88569 69957 88603 69991
rect 88603 69957 88612 69991
rect 88560 69948 88612 69957
rect 7140 69880 7192 69932
rect 84328 69812 84380 69864
rect 2908 69744 2960 69796
rect 5954 69606 6006 69658
rect 6018 69606 6070 69658
rect 6082 69606 6134 69658
rect 6146 69606 6198 69658
rect 6210 69606 6262 69658
rect 87098 69606 87150 69658
rect 87162 69606 87214 69658
rect 87226 69606 87278 69658
rect 87290 69606 87342 69658
rect 87354 69606 87406 69658
rect 89940 69268 89992 69320
rect 6690 69062 6742 69114
rect 6754 69062 6806 69114
rect 6818 69062 6870 69114
rect 6882 69062 6934 69114
rect 6946 69062 6998 69114
rect 87834 69062 87886 69114
rect 87898 69062 87950 69114
rect 87962 69062 88014 69114
rect 88026 69062 88078 69114
rect 88090 69062 88142 69114
rect 88652 68869 88704 68878
rect 7140 68792 7192 68844
rect 88652 68835 88667 68869
rect 88667 68835 88704 68869
rect 88652 68826 88704 68835
rect 2908 68656 2960 68708
rect 84328 68656 84380 68708
rect 5954 68518 6006 68570
rect 6018 68518 6070 68570
rect 6082 68518 6134 68570
rect 6146 68518 6198 68570
rect 6210 68518 6262 68570
rect 87098 68518 87150 68570
rect 87162 68518 87214 68570
rect 87226 68518 87278 68570
rect 87290 68518 87342 68570
rect 87354 68518 87406 68570
rect 6690 67974 6742 68026
rect 6754 67974 6806 68026
rect 6818 67974 6870 68026
rect 6882 67974 6934 68026
rect 6946 67974 6998 68026
rect 87834 67974 87886 68026
rect 87898 67974 87950 68026
rect 87962 67974 88014 68026
rect 88026 67974 88078 68026
rect 88090 67974 88142 68026
rect 88652 67781 88704 67790
rect 7140 67704 7192 67756
rect 88652 67747 88667 67781
rect 88667 67747 88704 67781
rect 88652 67738 88704 67747
rect 2908 67568 2960 67620
rect 84328 67568 84380 67620
rect 5954 67430 6006 67482
rect 6018 67430 6070 67482
rect 6082 67430 6134 67482
rect 6146 67430 6198 67482
rect 6210 67430 6262 67482
rect 87098 67430 87150 67482
rect 87162 67430 87214 67482
rect 87226 67430 87278 67482
rect 87290 67430 87342 67482
rect 87354 67430 87406 67482
rect 6690 66886 6742 66938
rect 6754 66886 6806 66938
rect 6818 66886 6870 66938
rect 6882 66886 6934 66938
rect 6946 66886 6998 66938
rect 87834 66886 87886 66938
rect 87898 66886 87950 66938
rect 87962 66886 88014 66938
rect 88026 66886 88078 66938
rect 88090 66886 88142 66938
rect 5484 66693 5536 66702
rect 5484 66659 5503 66693
rect 5503 66659 5536 66693
rect 5484 66650 5536 66659
rect 90124 66616 90176 66668
rect 4380 66480 4432 66532
rect 87456 66480 87508 66532
rect 5954 66342 6006 66394
rect 6018 66342 6070 66394
rect 6082 66342 6134 66394
rect 6146 66342 6198 66394
rect 6210 66342 6262 66394
rect 87098 66342 87150 66394
rect 87162 66342 87214 66394
rect 87226 66342 87278 66394
rect 87290 66342 87342 66394
rect 87354 66342 87406 66394
rect 6690 65798 6742 65850
rect 6754 65798 6806 65850
rect 6818 65798 6870 65850
rect 6882 65798 6934 65850
rect 6946 65798 6998 65850
rect 87834 65798 87886 65850
rect 87898 65798 87950 65850
rect 87962 65798 88014 65850
rect 88026 65798 88078 65850
rect 88090 65798 88142 65850
rect 5954 65254 6006 65306
rect 6018 65254 6070 65306
rect 6082 65254 6134 65306
rect 6146 65254 6198 65306
rect 6210 65254 6262 65306
rect 87098 65254 87150 65306
rect 87162 65254 87214 65306
rect 87226 65254 87278 65306
rect 87290 65254 87342 65306
rect 87354 65254 87406 65306
rect 5392 65095 5444 65104
rect 5392 65061 5410 65095
rect 5410 65061 5444 65095
rect 5392 65052 5444 65061
rect 2908 64916 2960 64968
rect 84328 64984 84380 65036
rect 89940 64848 89992 64900
rect 6690 64710 6742 64762
rect 6754 64710 6806 64762
rect 6818 64710 6870 64762
rect 6882 64710 6934 64762
rect 6946 64710 6998 64762
rect 87834 64710 87886 64762
rect 87898 64710 87950 64762
rect 87962 64710 88014 64762
rect 88026 64710 88078 64762
rect 88090 64710 88142 64762
rect 2908 64440 2960 64492
rect 84328 64440 84380 64492
rect 7232 64304 7284 64356
rect 88560 64347 88612 64356
rect 88560 64313 88583 64347
rect 88583 64313 88612 64347
rect 88560 64304 88612 64313
rect 5954 64166 6006 64218
rect 6018 64166 6070 64218
rect 6082 64166 6134 64218
rect 6146 64166 6198 64218
rect 6210 64166 6262 64218
rect 87098 64166 87150 64218
rect 87162 64166 87214 64218
rect 87226 64166 87278 64218
rect 87290 64166 87342 64218
rect 87354 64166 87406 64218
rect 6690 63622 6742 63674
rect 6754 63622 6806 63674
rect 6818 63622 6870 63674
rect 6882 63622 6934 63674
rect 6946 63622 6998 63674
rect 87834 63622 87886 63674
rect 87898 63622 87950 63674
rect 87962 63622 88014 63674
rect 88026 63622 88078 63674
rect 88090 63622 88142 63674
rect 2908 63352 2960 63404
rect 84328 63352 84380 63404
rect 7232 63216 7284 63268
rect 88560 63259 88612 63268
rect 88560 63225 88583 63259
rect 88583 63225 88612 63259
rect 88560 63216 88612 63225
rect 5954 63078 6006 63130
rect 6018 63078 6070 63130
rect 6082 63078 6134 63130
rect 6146 63078 6198 63130
rect 6210 63078 6262 63130
rect 87098 63078 87150 63130
rect 87162 63078 87214 63130
rect 87226 63078 87278 63130
rect 87290 63078 87342 63130
rect 87354 63078 87406 63130
rect 6690 62534 6742 62586
rect 6754 62534 6806 62586
rect 6818 62534 6870 62586
rect 6882 62534 6934 62586
rect 6946 62534 6998 62586
rect 87834 62534 87886 62586
rect 87898 62534 87950 62586
rect 87962 62534 88014 62586
rect 88026 62534 88078 62586
rect 88090 62534 88142 62586
rect 5208 62341 5260 62350
rect 5208 62307 5217 62341
rect 5217 62307 5251 62341
rect 5251 62307 5260 62341
rect 5208 62298 5260 62307
rect 9624 62332 9676 62384
rect 88376 62341 88428 62350
rect 88376 62307 88385 62341
rect 88385 62307 88419 62341
rect 88419 62307 88428 62341
rect 88376 62298 88428 62307
rect 89940 62332 89992 62384
rect 5954 61990 6006 62042
rect 6018 61990 6070 62042
rect 6082 61990 6134 62042
rect 6146 61990 6198 62042
rect 6210 61990 6262 62042
rect 87098 61990 87150 62042
rect 87162 61990 87214 62042
rect 87226 61990 87278 62042
rect 87290 61990 87342 62042
rect 87354 61990 87406 62042
rect 6690 61446 6742 61498
rect 6754 61446 6806 61498
rect 6818 61446 6870 61498
rect 6882 61446 6934 61498
rect 6946 61446 6998 61498
rect 87834 61446 87886 61498
rect 87898 61446 87950 61498
rect 87962 61446 88014 61498
rect 88026 61446 88078 61498
rect 88090 61446 88142 61498
rect 5208 61253 5260 61262
rect 5208 61219 5217 61253
rect 5217 61219 5251 61253
rect 5251 61219 5260 61253
rect 5208 61210 5260 61219
rect 88376 61253 88428 61262
rect 88376 61219 88385 61253
rect 88385 61219 88419 61253
rect 88419 61219 88428 61253
rect 88376 61210 88428 61219
rect 9624 61040 9676 61092
rect 89940 61040 89992 61092
rect 5954 60902 6006 60954
rect 6018 60902 6070 60954
rect 6082 60902 6134 60954
rect 6146 60902 6198 60954
rect 6210 60902 6262 60954
rect 87098 60902 87150 60954
rect 87162 60902 87214 60954
rect 87226 60902 87278 60954
rect 87290 60902 87342 60954
rect 87354 60902 87406 60954
rect 6690 60358 6742 60410
rect 6754 60358 6806 60410
rect 6818 60358 6870 60410
rect 6882 60358 6934 60410
rect 6946 60358 6998 60410
rect 87834 60358 87886 60410
rect 87898 60358 87950 60410
rect 87962 60358 88014 60410
rect 88026 60358 88078 60410
rect 88090 60358 88142 60410
rect 5954 59814 6006 59866
rect 6018 59814 6070 59866
rect 6082 59814 6134 59866
rect 6146 59814 6198 59866
rect 6210 59814 6262 59866
rect 87098 59814 87150 59866
rect 87162 59814 87214 59866
rect 87226 59814 87278 59866
rect 87290 59814 87342 59866
rect 87354 59814 87406 59866
rect 2908 59476 2960 59528
rect 5668 59476 5720 59528
rect 84328 59476 84380 59528
rect 89940 59408 89992 59460
rect 6690 59270 6742 59322
rect 6754 59270 6806 59322
rect 6818 59270 6870 59322
rect 6882 59270 6934 59322
rect 6946 59270 6998 59322
rect 87834 59270 87886 59322
rect 87898 59270 87950 59322
rect 87962 59270 88014 59322
rect 88026 59270 88078 59322
rect 88090 59270 88142 59322
rect 2908 59000 2960 59052
rect 84328 59000 84380 59052
rect 7232 58864 7284 58916
rect 88560 58907 88612 58916
rect 88560 58873 88583 58907
rect 88583 58873 88612 58907
rect 88560 58864 88612 58873
rect 5954 58726 6006 58778
rect 6018 58726 6070 58778
rect 6082 58726 6134 58778
rect 6146 58726 6198 58778
rect 6210 58726 6262 58778
rect 87098 58726 87150 58778
rect 87162 58726 87214 58778
rect 87226 58726 87278 58778
rect 87290 58726 87342 58778
rect 87354 58726 87406 58778
rect 6690 58182 6742 58234
rect 6754 58182 6806 58234
rect 6818 58182 6870 58234
rect 6882 58182 6934 58234
rect 6946 58182 6998 58234
rect 87834 58182 87886 58234
rect 87898 58182 87950 58234
rect 87962 58182 88014 58234
rect 88026 58182 88078 58234
rect 88090 58182 88142 58234
rect 2908 57912 2960 57964
rect 84328 57912 84380 57964
rect 7232 57776 7284 57828
rect 88560 57819 88612 57828
rect 88560 57785 88583 57819
rect 88583 57785 88612 57819
rect 88560 57776 88612 57785
rect 5954 57638 6006 57690
rect 6018 57638 6070 57690
rect 6082 57638 6134 57690
rect 6146 57638 6198 57690
rect 6210 57638 6262 57690
rect 87098 57638 87150 57690
rect 87162 57638 87214 57690
rect 87226 57638 87278 57690
rect 87290 57638 87342 57690
rect 87354 57638 87406 57690
rect 6690 57094 6742 57146
rect 6754 57094 6806 57146
rect 6818 57094 6870 57146
rect 6882 57094 6934 57146
rect 6946 57094 6998 57146
rect 87834 57094 87886 57146
rect 87898 57094 87950 57146
rect 87962 57094 88014 57146
rect 88026 57094 88078 57146
rect 88090 57094 88142 57146
rect 4932 56858 4984 56910
rect 5392 56867 5444 56876
rect 5392 56833 5410 56867
rect 5410 56833 5444 56867
rect 5392 56824 5444 56833
rect 88284 56858 88336 56910
rect 89940 56824 89992 56876
rect 5954 56550 6006 56602
rect 6018 56550 6070 56602
rect 6082 56550 6134 56602
rect 6146 56550 6198 56602
rect 6210 56550 6262 56602
rect 87098 56550 87150 56602
rect 87162 56550 87214 56602
rect 87226 56550 87278 56602
rect 87290 56550 87342 56602
rect 87354 56550 87406 56602
rect 6690 56006 6742 56058
rect 6754 56006 6806 56058
rect 6818 56006 6870 56058
rect 6882 56006 6934 56058
rect 6946 56006 6998 56058
rect 87834 56006 87886 56058
rect 87898 56006 87950 56058
rect 87962 56006 88014 56058
rect 88026 56006 88078 56058
rect 88090 56006 88142 56058
rect 5024 55770 5076 55822
rect 88376 55813 88428 55822
rect 88376 55779 88385 55813
rect 88385 55779 88419 55813
rect 88419 55779 88428 55813
rect 88376 55770 88428 55779
rect 5668 55600 5720 55652
rect 89940 55600 89992 55652
rect 5954 55462 6006 55514
rect 6018 55462 6070 55514
rect 6082 55462 6134 55514
rect 6146 55462 6198 55514
rect 6210 55462 6262 55514
rect 87098 55462 87150 55514
rect 87162 55462 87214 55514
rect 87226 55462 87278 55514
rect 87290 55462 87342 55514
rect 87354 55462 87406 55514
rect 2540 55124 2592 55176
rect 6690 54918 6742 54970
rect 6754 54918 6806 54970
rect 6818 54918 6870 54970
rect 6882 54918 6934 54970
rect 6946 54918 6998 54970
rect 87834 54918 87886 54970
rect 87898 54918 87950 54970
rect 87962 54918 88014 54970
rect 88026 54918 88078 54970
rect 88090 54918 88142 54970
rect 7600 54759 7652 54768
rect 7600 54725 7619 54759
rect 7619 54725 7652 54759
rect 7600 54716 7652 54725
rect 7048 54512 7100 54564
rect 5954 54374 6006 54426
rect 6018 54374 6070 54426
rect 6082 54374 6134 54426
rect 6146 54374 6198 54426
rect 6210 54374 6262 54426
rect 87098 54374 87150 54426
rect 87162 54374 87214 54426
rect 87226 54374 87278 54426
rect 87290 54374 87342 54426
rect 87354 54374 87406 54426
rect 84328 54104 84380 54156
rect 5208 54079 5260 54088
rect 5208 54045 5217 54079
rect 5217 54045 5251 54079
rect 5251 54045 5260 54079
rect 5208 54036 5260 54045
rect 89940 54036 89992 54088
rect 6690 53830 6742 53882
rect 6754 53830 6806 53882
rect 6818 53830 6870 53882
rect 6882 53830 6934 53882
rect 6946 53830 6998 53882
rect 87834 53830 87886 53882
rect 87898 53830 87950 53882
rect 87962 53830 88014 53882
rect 88026 53830 88078 53882
rect 88090 53830 88142 53882
rect 5668 53696 5720 53748
rect 2908 53560 2960 53612
rect 84328 53560 84380 53612
rect 88560 53467 88612 53476
rect 88560 53433 88583 53467
rect 88583 53433 88612 53467
rect 88560 53424 88612 53433
rect 5954 53286 6006 53338
rect 6018 53286 6070 53338
rect 6082 53286 6134 53338
rect 6146 53286 6198 53338
rect 6210 53286 6262 53338
rect 87098 53286 87150 53338
rect 87162 53286 87214 53338
rect 87226 53286 87278 53338
rect 87290 53286 87342 53338
rect 87354 53286 87406 53338
rect 7140 53152 7192 53204
rect 2908 52948 2960 53000
rect 89940 52948 89992 53000
rect 6690 52742 6742 52794
rect 6754 52742 6806 52794
rect 6818 52742 6870 52794
rect 6882 52742 6934 52794
rect 6946 52742 6998 52794
rect 87834 52742 87886 52794
rect 87898 52742 87950 52794
rect 87962 52742 88014 52794
rect 88026 52742 88078 52794
rect 88090 52742 88142 52794
rect 2908 52472 2960 52524
rect 84328 52472 84380 52524
rect 7140 52336 7192 52388
rect 88560 52379 88612 52388
rect 88560 52345 88583 52379
rect 88583 52345 88612 52379
rect 88560 52336 88612 52345
rect 5954 52198 6006 52250
rect 6018 52198 6070 52250
rect 6082 52198 6134 52250
rect 6146 52198 6198 52250
rect 6210 52198 6262 52250
rect 87098 52198 87150 52250
rect 87162 52198 87214 52250
rect 87226 52198 87278 52250
rect 87290 52198 87342 52250
rect 87354 52198 87406 52250
rect 6690 51654 6742 51706
rect 6754 51654 6806 51706
rect 6818 51654 6870 51706
rect 6882 51654 6934 51706
rect 6946 51654 6998 51706
rect 87834 51654 87886 51706
rect 87898 51654 87950 51706
rect 87962 51654 88014 51706
rect 88026 51654 88078 51706
rect 88090 51654 88142 51706
rect 2908 51384 2960 51436
rect 88376 51461 88428 51470
rect 88376 51427 88385 51461
rect 88385 51427 88419 51461
rect 88419 51427 88428 51461
rect 88376 51418 88428 51427
rect 5668 51316 5720 51368
rect 88560 51359 88612 51368
rect 88560 51325 88583 51359
rect 88583 51325 88612 51359
rect 88560 51316 88612 51325
rect 5954 51110 6006 51162
rect 6018 51110 6070 51162
rect 6082 51110 6134 51162
rect 6146 51110 6198 51162
rect 6210 51110 6262 51162
rect 87098 51110 87150 51162
rect 87162 51110 87214 51162
rect 87226 51110 87278 51162
rect 87290 51110 87342 51162
rect 87354 51110 87406 51162
rect 6690 50566 6742 50618
rect 6754 50566 6806 50618
rect 6818 50566 6870 50618
rect 6882 50566 6934 50618
rect 6946 50566 6998 50618
rect 87834 50566 87886 50618
rect 87898 50566 87950 50618
rect 87962 50566 88014 50618
rect 88026 50566 88078 50618
rect 88090 50566 88142 50618
rect 5954 50022 6006 50074
rect 6018 50022 6070 50074
rect 6082 50022 6134 50074
rect 6146 50022 6198 50074
rect 6210 50022 6262 50074
rect 87098 50022 87150 50074
rect 87162 50022 87214 50074
rect 87226 50022 87278 50074
rect 87290 50022 87342 50074
rect 87354 50022 87406 50074
rect 2908 49684 2960 49736
rect 89940 49684 89992 49736
rect 6690 49478 6742 49530
rect 6754 49478 6806 49530
rect 6818 49478 6870 49530
rect 6882 49478 6934 49530
rect 6946 49478 6998 49530
rect 87834 49478 87886 49530
rect 87898 49478 87950 49530
rect 87962 49478 88014 49530
rect 88026 49478 88078 49530
rect 88090 49478 88142 49530
rect 5954 48934 6006 48986
rect 6018 48934 6070 48986
rect 6082 48934 6134 48986
rect 6146 48934 6198 48986
rect 6210 48934 6262 48986
rect 87098 48934 87150 48986
rect 87162 48934 87214 48986
rect 87226 48934 87278 48986
rect 87290 48934 87342 48986
rect 87354 48934 87406 48986
rect 89940 48596 89992 48648
rect 6690 48390 6742 48442
rect 6754 48390 6806 48442
rect 6818 48390 6870 48442
rect 6882 48390 6934 48442
rect 6946 48390 6998 48442
rect 87834 48390 87886 48442
rect 87898 48390 87950 48442
rect 87962 48390 88014 48442
rect 88026 48390 88078 48442
rect 88090 48390 88142 48442
rect 5954 47846 6006 47898
rect 6018 47846 6070 47898
rect 6082 47846 6134 47898
rect 6146 47846 6198 47898
rect 6210 47846 6262 47898
rect 6690 47302 6742 47354
rect 6754 47302 6806 47354
rect 6818 47302 6870 47354
rect 6882 47302 6934 47354
rect 6946 47302 6998 47354
rect 12228 47304 12280 47356
rect 49230 47304 49282 47356
rect 51438 47304 51490 47356
rect 84420 47304 84472 47356
rect 8152 47236 8204 47288
rect 14436 47236 14488 47288
rect 7876 47168 7928 47220
rect 12200 47168 12252 47220
rect 48172 47168 48224 47220
rect 88560 48027 88612 48036
rect 88560 47993 88583 48027
rect 88583 47993 88612 48027
rect 88560 47984 88612 47993
rect 87098 47846 87150 47898
rect 87162 47846 87214 47898
rect 87226 47846 87278 47898
rect 87290 47846 87342 47898
rect 87354 47846 87406 47898
rect 87834 47302 87886 47354
rect 87898 47302 87950 47354
rect 87962 47302 88014 47354
rect 88026 47302 88078 47354
rect 88090 47302 88142 47354
rect 2908 47100 2960 47152
rect 7048 47100 7100 47152
rect 11004 47100 11056 47152
rect 14132 46896 14184 46948
rect 88560 46939 88612 46948
rect 88560 46905 88569 46939
rect 88569 46905 88603 46939
rect 88603 46905 88612 46939
rect 88560 46896 88612 46905
rect 13580 46828 13632 46880
rect 50196 46828 50248 46880
rect 5954 46758 6006 46810
rect 6018 46758 6070 46810
rect 6082 46758 6134 46810
rect 6146 46758 6198 46810
rect 6210 46758 6262 46810
rect 12476 46760 12528 46812
rect 49092 46760 49144 46812
rect 50656 46760 50708 46812
rect 84052 46760 84104 46812
rect 87098 46758 87150 46810
rect 87162 46758 87214 46810
rect 87226 46758 87278 46810
rect 87290 46758 87342 46810
rect 87354 46758 87406 46810
rect 11004 46692 11056 46744
rect 47804 46692 47856 46744
rect 49552 46692 49604 46744
rect 83684 46692 83736 46744
rect 6690 46214 6742 46266
rect 6754 46214 6806 46266
rect 6818 46214 6870 46266
rect 6882 46214 6934 46266
rect 6946 46214 6998 46266
rect 87834 46214 87886 46266
rect 87898 46214 87950 46266
rect 87962 46214 88014 46266
rect 88026 46214 88078 46266
rect 88090 46214 88142 46266
rect 2908 45808 2960 45860
rect 5954 45670 6006 45722
rect 6018 45670 6070 45722
rect 6082 45670 6134 45722
rect 6146 45670 6198 45722
rect 6210 45670 6262 45722
rect 87098 45670 87150 45722
rect 87162 45670 87214 45722
rect 87226 45670 87278 45722
rect 87290 45670 87342 45722
rect 87354 45670 87406 45722
rect 6690 45126 6742 45178
rect 6754 45126 6806 45178
rect 6818 45126 6870 45178
rect 6882 45126 6934 45178
rect 6946 45126 6998 45178
rect 87834 45126 87886 45178
rect 87898 45126 87950 45178
rect 87962 45126 88014 45178
rect 88026 45126 88078 45178
rect 88090 45126 88142 45178
rect 2540 44720 2592 44772
rect 5954 44582 6006 44634
rect 6018 44582 6070 44634
rect 6082 44582 6134 44634
rect 6146 44582 6198 44634
rect 6210 44582 6262 44634
rect 87098 44582 87150 44634
rect 87162 44582 87214 44634
rect 87226 44582 87278 44634
rect 87290 44582 87342 44634
rect 87354 44582 87406 44634
rect 5208 44423 5260 44432
rect 5208 44389 5217 44423
rect 5217 44389 5251 44423
rect 5251 44389 5260 44423
rect 5208 44380 5260 44389
rect 6690 44038 6742 44090
rect 6754 44038 6806 44090
rect 6818 44038 6870 44090
rect 6882 44038 6934 44090
rect 6946 44038 6998 44090
rect 87834 44038 87886 44090
rect 87898 44038 87950 44090
rect 87962 44038 88014 44090
rect 88026 44038 88078 44090
rect 88090 44038 88142 44090
rect 5954 43494 6006 43546
rect 6018 43494 6070 43546
rect 6082 43494 6134 43546
rect 6146 43494 6198 43546
rect 6210 43494 6262 43546
rect 87098 43494 87150 43546
rect 87162 43494 87214 43546
rect 87226 43494 87278 43546
rect 87290 43494 87342 43546
rect 87354 43494 87406 43546
rect 89940 43224 89992 43276
rect 7140 43156 7192 43208
rect 2908 43088 2960 43140
rect 84328 43088 84380 43140
rect 6690 42950 6742 43002
rect 6754 42950 6806 43002
rect 6818 42950 6870 43002
rect 6882 42950 6934 43002
rect 6946 42950 6998 43002
rect 87834 42950 87886 43002
rect 87898 42950 87950 43002
rect 87962 42950 88014 43002
rect 88026 42950 88078 43002
rect 88090 42950 88142 43002
rect 2908 42544 2960 42596
rect 5954 42406 6006 42458
rect 6018 42406 6070 42458
rect 6082 42406 6134 42458
rect 6146 42406 6198 42458
rect 6210 42406 6262 42458
rect 87098 42406 87150 42458
rect 87162 42406 87214 42458
rect 87226 42406 87278 42458
rect 87290 42406 87342 42458
rect 87354 42406 87406 42458
rect 88560 42145 88612 42154
rect 7140 42068 7192 42120
rect 88560 42111 88579 42145
rect 88579 42111 88612 42145
rect 88560 42102 88612 42111
rect 2908 42000 2960 42052
rect 84328 42000 84380 42052
rect 6690 41862 6742 41914
rect 6754 41862 6806 41914
rect 6818 41862 6870 41914
rect 6882 41862 6934 41914
rect 6946 41862 6998 41914
rect 87834 41862 87886 41914
rect 87898 41862 87950 41914
rect 87962 41862 88014 41914
rect 88026 41862 88078 41914
rect 88090 41862 88142 41914
rect 4380 41728 4432 41780
rect 87456 41728 87508 41780
rect 5668 41626 5720 41678
rect 89940 41660 89992 41712
rect 5954 41318 6006 41370
rect 6018 41318 6070 41370
rect 6082 41318 6134 41370
rect 6146 41318 6198 41370
rect 6210 41318 6262 41370
rect 87098 41318 87150 41370
rect 87162 41318 87214 41370
rect 87226 41318 87278 41370
rect 87290 41318 87342 41370
rect 87354 41318 87406 41370
rect 6690 40774 6742 40826
rect 6754 40774 6806 40826
rect 6818 40774 6870 40826
rect 6882 40774 6934 40826
rect 6946 40774 6998 40826
rect 87834 40774 87886 40826
rect 87898 40774 87950 40826
rect 87962 40774 88014 40826
rect 88026 40774 88078 40826
rect 88090 40774 88142 40826
rect 5954 40230 6006 40282
rect 6018 40230 6070 40282
rect 6082 40230 6134 40282
rect 6146 40230 6198 40282
rect 6210 40230 6262 40282
rect 87098 40230 87150 40282
rect 87162 40230 87214 40282
rect 87226 40230 87278 40282
rect 87290 40230 87342 40282
rect 87354 40230 87406 40282
rect 7140 39892 7192 39944
rect 84328 39892 84380 39944
rect 89940 39892 89992 39944
rect 2908 39824 2960 39876
rect 6690 39686 6742 39738
rect 6754 39686 6806 39738
rect 6818 39686 6870 39738
rect 6882 39686 6934 39738
rect 6946 39686 6998 39738
rect 87834 39686 87886 39738
rect 87898 39686 87950 39738
rect 87962 39686 88014 39738
rect 88026 39686 88078 39738
rect 88090 39686 88142 39738
rect 5954 39142 6006 39194
rect 6018 39142 6070 39194
rect 6082 39142 6134 39194
rect 6146 39142 6198 39194
rect 6210 39142 6262 39194
rect 87098 39142 87150 39194
rect 87162 39142 87214 39194
rect 87226 39142 87278 39194
rect 87290 39142 87342 39194
rect 87354 39142 87406 39194
rect 4380 38940 4432 38992
rect 87180 38940 87232 38992
rect 7416 38804 7468 38856
rect 89296 38804 89348 38856
rect 6690 38598 6742 38650
rect 6754 38598 6806 38650
rect 6818 38598 6870 38650
rect 6882 38598 6934 38650
rect 6946 38598 6998 38650
rect 87834 38598 87886 38650
rect 87898 38598 87950 38650
rect 87962 38598 88014 38650
rect 88026 38598 88078 38650
rect 88090 38598 88142 38650
rect 5954 38054 6006 38106
rect 6018 38054 6070 38106
rect 6082 38054 6134 38106
rect 6146 38054 6198 38106
rect 6210 38054 6262 38106
rect 87098 38054 87150 38106
rect 87162 38054 87214 38106
rect 87226 38054 87278 38106
rect 87290 38054 87342 38106
rect 87354 38054 87406 38106
rect 7140 37716 7192 37768
rect 84328 37716 84380 37768
rect 89940 37716 89992 37768
rect 2908 37648 2960 37700
rect 6690 37510 6742 37562
rect 6754 37510 6806 37562
rect 6818 37510 6870 37562
rect 6882 37510 6934 37562
rect 6946 37510 6998 37562
rect 87834 37510 87886 37562
rect 87898 37510 87950 37562
rect 87962 37510 88014 37562
rect 88026 37510 88078 37562
rect 88090 37510 88142 37562
rect 5954 36966 6006 37018
rect 6018 36966 6070 37018
rect 6082 36966 6134 37018
rect 6146 36966 6198 37018
rect 6210 36966 6262 37018
rect 87098 36966 87150 37018
rect 87162 36966 87214 37018
rect 87226 36966 87278 37018
rect 87290 36966 87342 37018
rect 87354 36966 87406 37018
rect 7140 36628 7192 36680
rect 84328 36628 84380 36680
rect 89940 36628 89992 36680
rect 2908 36560 2960 36612
rect 6690 36422 6742 36474
rect 6754 36422 6806 36474
rect 6818 36422 6870 36474
rect 6882 36422 6934 36474
rect 6946 36422 6998 36474
rect 87834 36422 87886 36474
rect 87898 36422 87950 36474
rect 87962 36422 88014 36474
rect 88026 36422 88078 36474
rect 88090 36422 88142 36474
rect 5668 36186 5720 36238
rect 90124 36152 90176 36204
rect 4380 36084 4432 36136
rect 87456 36084 87508 36136
rect 5954 35878 6006 35930
rect 6018 35878 6070 35930
rect 6082 35878 6134 35930
rect 6146 35878 6198 35930
rect 6210 35878 6262 35930
rect 87098 35878 87150 35930
rect 87162 35878 87214 35930
rect 87226 35878 87278 35930
rect 87290 35878 87342 35930
rect 87354 35878 87406 35930
rect 6690 35334 6742 35386
rect 6754 35334 6806 35386
rect 6818 35334 6870 35386
rect 6882 35334 6934 35386
rect 6946 35334 6998 35386
rect 87834 35334 87886 35386
rect 87898 35334 87950 35386
rect 87962 35334 88014 35386
rect 88026 35334 88078 35386
rect 88090 35334 88142 35386
rect 5954 34790 6006 34842
rect 6018 34790 6070 34842
rect 6082 34790 6134 34842
rect 6146 34790 6198 34842
rect 6210 34790 6262 34842
rect 87098 34790 87150 34842
rect 87162 34790 87214 34842
rect 87226 34790 87278 34842
rect 87290 34790 87342 34842
rect 87354 34790 87406 34842
rect 88560 34523 88612 34532
rect 7140 34452 7192 34504
rect 88560 34489 88575 34523
rect 88575 34489 88612 34523
rect 88560 34480 88612 34489
rect 2908 34384 2960 34436
rect 84328 34384 84380 34436
rect 6690 34246 6742 34298
rect 6754 34246 6806 34298
rect 6818 34246 6870 34298
rect 6882 34246 6934 34298
rect 6946 34246 6998 34298
rect 87834 34246 87886 34298
rect 87898 34246 87950 34298
rect 87962 34246 88014 34298
rect 88026 34246 88078 34298
rect 88090 34246 88142 34298
rect 2908 33840 2960 33892
rect 5954 33702 6006 33754
rect 6018 33702 6070 33754
rect 6082 33702 6134 33754
rect 6146 33702 6198 33754
rect 6210 33702 6262 33754
rect 87098 33702 87150 33754
rect 87162 33702 87214 33754
rect 87226 33702 87278 33754
rect 87290 33702 87342 33754
rect 87354 33702 87406 33754
rect 4380 33500 4432 33552
rect 5668 33398 5720 33450
rect 87180 33364 87232 33416
rect 89940 33364 89992 33416
rect 6690 33158 6742 33210
rect 6754 33158 6806 33210
rect 6818 33158 6870 33210
rect 6882 33158 6934 33210
rect 6946 33158 6998 33210
rect 87834 33158 87886 33210
rect 87898 33158 87950 33210
rect 87962 33158 88014 33210
rect 88026 33158 88078 33210
rect 88090 33158 88142 33210
rect 5954 32614 6006 32666
rect 6018 32614 6070 32666
rect 6082 32614 6134 32666
rect 6146 32614 6198 32666
rect 6210 32614 6262 32666
rect 87098 32614 87150 32666
rect 87162 32614 87214 32666
rect 87226 32614 87278 32666
rect 87290 32614 87342 32666
rect 87354 32614 87406 32666
rect 7140 32276 7192 32328
rect 84328 32276 84380 32328
rect 89940 32276 89992 32328
rect 2908 32208 2960 32260
rect 6690 32070 6742 32122
rect 6754 32070 6806 32122
rect 6818 32070 6870 32122
rect 6882 32070 6934 32122
rect 6946 32070 6998 32122
rect 87834 32070 87886 32122
rect 87898 32070 87950 32122
rect 87962 32070 88014 32122
rect 88026 32070 88078 32122
rect 88090 32070 88142 32122
rect 5954 31526 6006 31578
rect 6018 31526 6070 31578
rect 6082 31526 6134 31578
rect 6146 31526 6198 31578
rect 6210 31526 6262 31578
rect 87098 31526 87150 31578
rect 87162 31526 87214 31578
rect 87226 31526 87278 31578
rect 87290 31526 87342 31578
rect 87354 31526 87406 31578
rect 88560 31259 88612 31268
rect 7140 31188 7192 31240
rect 88560 31225 88575 31259
rect 88575 31225 88612 31259
rect 88560 31216 88612 31225
rect 2908 31120 2960 31172
rect 84328 31120 84380 31172
rect 6690 30982 6742 31034
rect 6754 30982 6806 31034
rect 6818 30982 6870 31034
rect 6882 30982 6934 31034
rect 6946 30982 6998 31034
rect 87834 30982 87886 31034
rect 87898 30982 87950 31034
rect 87962 30982 88014 31034
rect 88026 30982 88078 31034
rect 88090 30982 88142 31034
rect 5668 30746 5720 30798
rect 89940 30712 89992 30764
rect 4380 30576 4432 30628
rect 87456 30576 87508 30628
rect 5954 30438 6006 30490
rect 6018 30438 6070 30490
rect 6082 30438 6134 30490
rect 6146 30438 6198 30490
rect 6210 30438 6262 30490
rect 87098 30438 87150 30490
rect 87162 30438 87214 30490
rect 87226 30438 87278 30490
rect 87290 30438 87342 30490
rect 87354 30438 87406 30490
rect 6690 29894 6742 29946
rect 6754 29894 6806 29946
rect 6818 29894 6870 29946
rect 6882 29894 6934 29946
rect 6946 29894 6998 29946
rect 87834 29894 87886 29946
rect 87898 29894 87950 29946
rect 87962 29894 88014 29946
rect 88026 29894 88078 29946
rect 88090 29894 88142 29946
rect 5954 29350 6006 29402
rect 6018 29350 6070 29402
rect 6082 29350 6134 29402
rect 6146 29350 6198 29402
rect 6210 29350 6262 29402
rect 87098 29350 87150 29402
rect 87162 29350 87214 29402
rect 87226 29350 87278 29402
rect 87290 29350 87342 29402
rect 87354 29350 87406 29402
rect 88560 29083 88612 29092
rect 7140 29012 7192 29064
rect 88560 29049 88575 29083
rect 88575 29049 88612 29083
rect 88560 29040 88612 29049
rect 2908 28944 2960 28996
rect 84328 28944 84380 28996
rect 6690 28806 6742 28858
rect 6754 28806 6806 28858
rect 6818 28806 6870 28858
rect 6882 28806 6934 28858
rect 6946 28806 6998 28858
rect 87834 28806 87886 28858
rect 87898 28806 87950 28858
rect 87962 28806 88014 28858
rect 88026 28806 88078 28858
rect 88090 28806 88142 28858
rect 5954 28262 6006 28314
rect 6018 28262 6070 28314
rect 6082 28262 6134 28314
rect 6146 28262 6198 28314
rect 6210 28262 6262 28314
rect 87098 28262 87150 28314
rect 87162 28262 87214 28314
rect 87226 28262 87278 28314
rect 87290 28262 87342 28314
rect 87354 28262 87406 28314
rect 5116 27958 5168 28010
rect 87548 27924 87600 27976
rect 5392 27899 5444 27908
rect 5392 27865 5410 27899
rect 5410 27865 5444 27899
rect 5392 27856 5444 27865
rect 89940 27856 89992 27908
rect 6690 27718 6742 27770
rect 6754 27718 6806 27770
rect 6818 27718 6870 27770
rect 6882 27718 6934 27770
rect 6946 27718 6998 27770
rect 87834 27718 87886 27770
rect 87898 27718 87950 27770
rect 87962 27718 88014 27770
rect 88026 27718 88078 27770
rect 88090 27718 88142 27770
rect 5954 27174 6006 27226
rect 6018 27174 6070 27226
rect 6082 27174 6134 27226
rect 6146 27174 6198 27226
rect 6210 27174 6262 27226
rect 87098 27174 87150 27226
rect 87162 27174 87214 27226
rect 87226 27174 87278 27226
rect 87290 27174 87342 27226
rect 87354 27174 87406 27226
rect 2908 26836 2960 26888
rect 84328 26836 84380 26888
rect 7140 26768 7192 26820
rect 89940 26768 89992 26820
rect 6690 26630 6742 26682
rect 6754 26630 6806 26682
rect 6818 26630 6870 26682
rect 6882 26630 6934 26682
rect 6946 26630 6998 26682
rect 87834 26630 87886 26682
rect 87898 26630 87950 26682
rect 87962 26630 88014 26682
rect 88026 26630 88078 26682
rect 88090 26630 88142 26682
rect 5954 26086 6006 26138
rect 6018 26086 6070 26138
rect 6082 26086 6134 26138
rect 6146 26086 6198 26138
rect 6210 26086 6262 26138
rect 87098 26086 87150 26138
rect 87162 26086 87214 26138
rect 87226 26086 87278 26138
rect 87290 26086 87342 26138
rect 87354 26086 87406 26138
rect 2908 25748 2960 25800
rect 84328 25748 84380 25800
rect 7140 25680 7192 25732
rect 89940 25680 89992 25732
rect 6690 25542 6742 25594
rect 6754 25542 6806 25594
rect 6818 25542 6870 25594
rect 6882 25542 6934 25594
rect 6946 25542 6998 25594
rect 87834 25542 87886 25594
rect 87898 25542 87950 25594
rect 87962 25542 88014 25594
rect 88026 25542 88078 25594
rect 88090 25542 88142 25594
rect 4932 25306 4984 25358
rect 88376 25349 88428 25358
rect 88376 25315 88385 25349
rect 88385 25315 88419 25349
rect 88419 25315 88428 25349
rect 88376 25306 88428 25315
rect 5668 25136 5720 25188
rect 89940 25136 89992 25188
rect 5954 24998 6006 25050
rect 6018 24998 6070 25050
rect 6082 24998 6134 25050
rect 6146 24998 6198 25050
rect 6210 24998 6262 25050
rect 87098 24998 87150 25050
rect 87162 24998 87214 25050
rect 87226 24998 87278 25050
rect 87290 24998 87342 25050
rect 87354 24998 87406 25050
rect 6690 24454 6742 24506
rect 6754 24454 6806 24506
rect 6818 24454 6870 24506
rect 6882 24454 6934 24506
rect 6946 24454 6998 24506
rect 87834 24454 87886 24506
rect 87898 24454 87950 24506
rect 87962 24454 88014 24506
rect 88026 24454 88078 24506
rect 88090 24454 88142 24506
rect 5954 23910 6006 23962
rect 6018 23910 6070 23962
rect 6082 23910 6134 23962
rect 6146 23910 6198 23962
rect 6210 23910 6262 23962
rect 87098 23910 87150 23962
rect 87162 23910 87214 23962
rect 87226 23910 87278 23962
rect 87290 23910 87342 23962
rect 87354 23910 87406 23962
rect 2908 23572 2960 23624
rect 84328 23572 84380 23624
rect 7140 23504 7192 23556
rect 89940 23504 89992 23556
rect 6690 23366 6742 23418
rect 6754 23366 6806 23418
rect 6818 23366 6870 23418
rect 6882 23366 6934 23418
rect 6946 23366 6998 23418
rect 87834 23366 87886 23418
rect 87898 23366 87950 23418
rect 87962 23366 88014 23418
rect 88026 23366 88078 23418
rect 88090 23366 88142 23418
rect 5954 22822 6006 22874
rect 6018 22822 6070 22874
rect 6082 22822 6134 22874
rect 6146 22822 6198 22874
rect 6210 22822 6262 22874
rect 87098 22822 87150 22874
rect 87162 22822 87214 22874
rect 87226 22822 87278 22874
rect 87290 22822 87342 22874
rect 87354 22822 87406 22874
rect 5208 22561 5260 22570
rect 5208 22527 5217 22561
rect 5217 22527 5251 22561
rect 5251 22527 5260 22561
rect 5208 22518 5260 22527
rect 84328 22484 84380 22536
rect 7140 22416 7192 22468
rect 89940 22416 89992 22468
rect 6690 22278 6742 22330
rect 6754 22278 6806 22330
rect 6818 22278 6870 22330
rect 6882 22278 6934 22330
rect 6946 22278 6998 22330
rect 87834 22278 87886 22330
rect 87898 22278 87950 22330
rect 87962 22278 88014 22330
rect 88026 22278 88078 22330
rect 88090 22278 88142 22330
rect 5954 21734 6006 21786
rect 6018 21734 6070 21786
rect 6082 21734 6134 21786
rect 6146 21734 6198 21786
rect 6210 21734 6262 21786
rect 87098 21734 87150 21786
rect 87162 21734 87214 21786
rect 87226 21734 87278 21786
rect 87290 21734 87342 21786
rect 87354 21734 87406 21786
rect 2908 21396 2960 21448
rect 84328 21396 84380 21448
rect 7140 21328 7192 21380
rect 89940 21328 89992 21380
rect 6690 21190 6742 21242
rect 6754 21190 6806 21242
rect 6818 21190 6870 21242
rect 6882 21190 6934 21242
rect 6946 21190 6998 21242
rect 87834 21190 87886 21242
rect 87898 21190 87950 21242
rect 87962 21190 88014 21242
rect 88026 21190 88078 21242
rect 88090 21190 88142 21242
rect 5954 20646 6006 20698
rect 6018 20646 6070 20698
rect 6082 20646 6134 20698
rect 6146 20646 6198 20698
rect 6210 20646 6262 20698
rect 87098 20646 87150 20698
rect 87162 20646 87214 20698
rect 87226 20646 87278 20698
rect 87290 20646 87342 20698
rect 87354 20646 87406 20698
rect 2908 20308 2960 20360
rect 84328 20308 84380 20360
rect 7140 20240 7192 20292
rect 89940 20240 89992 20292
rect 6690 20102 6742 20154
rect 6754 20102 6806 20154
rect 6818 20102 6870 20154
rect 6882 20102 6934 20154
rect 6946 20102 6998 20154
rect 87834 20102 87886 20154
rect 87898 20102 87950 20154
rect 87962 20102 88014 20154
rect 88026 20102 88078 20154
rect 88090 20102 88142 20154
rect 4932 19866 4984 19918
rect 88376 19909 88428 19918
rect 88376 19875 88385 19909
rect 88385 19875 88419 19909
rect 88419 19875 88428 19909
rect 88376 19866 88428 19875
rect 9624 19696 9676 19748
rect 90032 19696 90084 19748
rect 5954 19558 6006 19610
rect 6018 19558 6070 19610
rect 6082 19558 6134 19610
rect 6146 19558 6198 19610
rect 6210 19558 6262 19610
rect 87098 19558 87150 19610
rect 87162 19558 87214 19610
rect 87226 19558 87278 19610
rect 87290 19558 87342 19610
rect 87354 19558 87406 19610
rect 6690 19014 6742 19066
rect 6754 19014 6806 19066
rect 6818 19014 6870 19066
rect 6882 19014 6934 19066
rect 6946 19014 6998 19066
rect 87834 19014 87886 19066
rect 87898 19014 87950 19066
rect 87962 19014 88014 19066
rect 88026 19014 88078 19066
rect 88090 19014 88142 19066
rect 5954 18470 6006 18522
rect 6018 18470 6070 18522
rect 6082 18470 6134 18522
rect 6146 18470 6198 18522
rect 6210 18470 6262 18522
rect 87098 18470 87150 18522
rect 87162 18470 87214 18522
rect 87226 18470 87278 18522
rect 87290 18470 87342 18522
rect 87354 18470 87406 18522
rect 5116 18166 5168 18218
rect 9624 18200 9676 18252
rect 88192 18166 88244 18218
rect 89940 18200 89992 18252
rect 6690 17926 6742 17978
rect 6754 17926 6806 17978
rect 6818 17926 6870 17978
rect 6882 17926 6934 17978
rect 6946 17926 6998 17978
rect 87834 17926 87886 17978
rect 87898 17926 87950 17978
rect 87962 17926 88014 17978
rect 88026 17926 88078 17978
rect 88090 17926 88142 17978
rect 5954 17382 6006 17434
rect 6018 17382 6070 17434
rect 6082 17382 6134 17434
rect 6146 17382 6198 17434
rect 6210 17382 6262 17434
rect 87098 17382 87150 17434
rect 87162 17382 87214 17434
rect 87226 17382 87278 17434
rect 87290 17382 87342 17434
rect 87354 17382 87406 17434
rect 5208 17121 5260 17130
rect 5208 17087 5217 17121
rect 5217 17087 5251 17121
rect 5251 17087 5260 17121
rect 5208 17078 5260 17087
rect 84328 17044 84380 17096
rect 7140 16976 7192 17028
rect 89940 16976 89992 17028
rect 6690 16838 6742 16890
rect 6754 16838 6806 16890
rect 6818 16838 6870 16890
rect 6882 16838 6934 16890
rect 6946 16838 6998 16890
rect 87834 16838 87886 16890
rect 87898 16838 87950 16890
rect 87962 16838 88014 16890
rect 88026 16838 88078 16890
rect 88090 16838 88142 16890
rect 5954 16294 6006 16346
rect 6018 16294 6070 16346
rect 6082 16294 6134 16346
rect 6146 16294 6198 16346
rect 6210 16294 6262 16346
rect 87098 16294 87150 16346
rect 87162 16294 87214 16346
rect 87226 16294 87278 16346
rect 87290 16294 87342 16346
rect 87354 16294 87406 16346
rect 2908 15956 2960 16008
rect 84328 15956 84380 16008
rect 7600 15888 7652 15940
rect 89940 15888 89992 15940
rect 6690 15750 6742 15802
rect 6754 15750 6806 15802
rect 6818 15750 6870 15802
rect 6882 15750 6934 15802
rect 6946 15750 6998 15802
rect 87834 15750 87886 15802
rect 87898 15750 87950 15802
rect 87962 15750 88014 15802
rect 88026 15750 88078 15802
rect 88090 15750 88142 15802
rect 5954 15206 6006 15258
rect 6018 15206 6070 15258
rect 6082 15206 6134 15258
rect 6146 15206 6198 15258
rect 6210 15206 6262 15258
rect 87098 15206 87150 15258
rect 87162 15206 87214 15258
rect 87226 15206 87278 15258
rect 87290 15206 87342 15258
rect 87354 15206 87406 15258
rect 2908 14868 2960 14920
rect 84328 14868 84380 14920
rect 7600 14800 7652 14852
rect 89940 14800 89992 14852
rect 6690 14662 6742 14714
rect 6754 14662 6806 14714
rect 6818 14662 6870 14714
rect 6882 14662 6934 14714
rect 6946 14662 6998 14714
rect 87834 14662 87886 14714
rect 87898 14662 87950 14714
rect 87962 14662 88014 14714
rect 88026 14662 88078 14714
rect 88090 14662 88142 14714
rect 4932 14426 4984 14478
rect 88376 14469 88428 14478
rect 88376 14435 88385 14469
rect 88385 14435 88419 14469
rect 88419 14435 88428 14469
rect 88376 14426 88428 14435
rect 5668 14256 5720 14308
rect 89940 14256 89992 14308
rect 5954 14118 6006 14170
rect 6018 14118 6070 14170
rect 6082 14118 6134 14170
rect 6146 14118 6198 14170
rect 6210 14118 6262 14170
rect 87098 14118 87150 14170
rect 87162 14118 87214 14170
rect 87226 14118 87278 14170
rect 87290 14118 87342 14170
rect 87354 14118 87406 14170
rect 6690 13574 6742 13626
rect 6754 13574 6806 13626
rect 6818 13574 6870 13626
rect 6882 13574 6934 13626
rect 6946 13574 6998 13626
rect 87834 13574 87886 13626
rect 87898 13574 87950 13626
rect 87962 13574 88014 13626
rect 88026 13574 88078 13626
rect 88090 13574 88142 13626
rect 5954 13030 6006 13082
rect 6018 13030 6070 13082
rect 6082 13030 6134 13082
rect 6146 13030 6198 13082
rect 6210 13030 6262 13082
rect 87098 13030 87150 13082
rect 87162 13030 87214 13082
rect 87226 13030 87278 13082
rect 87290 13030 87342 13082
rect 87354 13030 87406 13082
rect 6690 12486 6742 12538
rect 6754 12486 6806 12538
rect 6818 12486 6870 12538
rect 6882 12486 6934 12538
rect 6946 12486 6998 12538
rect 87834 12486 87886 12538
rect 87898 12486 87950 12538
rect 87962 12486 88014 12538
rect 88026 12486 88078 12538
rect 88090 12486 88142 12538
rect 5954 11942 6006 11994
rect 6018 11942 6070 11994
rect 6082 11942 6134 11994
rect 6146 11942 6198 11994
rect 6210 11942 6262 11994
rect 87098 11942 87150 11994
rect 87162 11942 87214 11994
rect 87226 11942 87278 11994
rect 87290 11942 87342 11994
rect 87354 11942 87406 11994
rect 6690 11398 6742 11450
rect 6754 11398 6806 11450
rect 6818 11398 6870 11450
rect 6882 11398 6934 11450
rect 6946 11398 6998 11450
rect 87834 11398 87886 11450
rect 87898 11398 87950 11450
rect 87962 11398 88014 11450
rect 88026 11398 88078 11450
rect 88090 11398 88142 11450
rect 5954 10854 6006 10906
rect 6018 10854 6070 10906
rect 6082 10854 6134 10906
rect 6146 10854 6198 10906
rect 6210 10854 6262 10906
rect 87098 10854 87150 10906
rect 87162 10854 87214 10906
rect 87226 10854 87278 10906
rect 87290 10854 87342 10906
rect 87354 10854 87406 10906
rect 6690 10310 6742 10362
rect 6754 10310 6806 10362
rect 6818 10310 6870 10362
rect 6882 10310 6934 10362
rect 6946 10310 6998 10362
rect 87834 10310 87886 10362
rect 87898 10310 87950 10362
rect 87962 10310 88014 10362
rect 88026 10310 88078 10362
rect 88090 10310 88142 10362
rect 5954 9766 6006 9818
rect 6018 9766 6070 9818
rect 6082 9766 6134 9818
rect 6146 9766 6198 9818
rect 6210 9766 6262 9818
rect 87098 9766 87150 9818
rect 87162 9766 87214 9818
rect 87226 9766 87278 9818
rect 87290 9766 87342 9818
rect 87354 9766 87406 9818
rect 6690 9222 6742 9274
rect 6754 9222 6806 9274
rect 6818 9222 6870 9274
rect 6882 9222 6934 9274
rect 6946 9222 6998 9274
rect 87834 9222 87886 9274
rect 87898 9222 87950 9274
rect 87962 9222 88014 9274
rect 88026 9222 88078 9274
rect 88090 9222 88142 9274
rect 5954 8678 6006 8730
rect 6018 8678 6070 8730
rect 6082 8678 6134 8730
rect 6146 8678 6198 8730
rect 6210 8678 6262 8730
rect 87098 8678 87150 8730
rect 87162 8678 87214 8730
rect 87226 8678 87278 8730
rect 87290 8678 87342 8730
rect 87354 8678 87406 8730
rect 6690 8134 6742 8186
rect 6754 8134 6806 8186
rect 6818 8134 6870 8186
rect 6882 8134 6934 8186
rect 6946 8134 6998 8186
rect 87834 8134 87886 8186
rect 87898 8134 87950 8186
rect 87962 8134 88014 8186
rect 88026 8134 88078 8186
rect 88090 8134 88142 8186
rect 5954 7590 6006 7642
rect 6018 7590 6070 7642
rect 6082 7590 6134 7642
rect 6146 7590 6198 7642
rect 6210 7590 6262 7642
rect 18722 7590 18774 7642
rect 18786 7590 18838 7642
rect 18850 7590 18902 7642
rect 18914 7590 18966 7642
rect 18978 7590 19030 7642
rect 37722 7590 37774 7642
rect 37786 7590 37838 7642
rect 37850 7590 37902 7642
rect 37914 7590 37966 7642
rect 37978 7590 38030 7642
rect 56722 7590 56774 7642
rect 56786 7590 56838 7642
rect 56850 7590 56902 7642
rect 56914 7590 56966 7642
rect 56978 7590 57030 7642
rect 75722 7590 75774 7642
rect 75786 7590 75838 7642
rect 75850 7590 75902 7642
rect 75914 7590 75966 7642
rect 75978 7590 76030 7642
rect 87098 7590 87150 7642
rect 87162 7590 87214 7642
rect 87226 7590 87278 7642
rect 87290 7590 87342 7642
rect 87354 7590 87406 7642
rect 6690 7046 6742 7098
rect 6754 7046 6806 7098
rect 6818 7046 6870 7098
rect 6882 7046 6934 7098
rect 6946 7046 6998 7098
rect 19382 7046 19434 7098
rect 19446 7046 19498 7098
rect 19510 7046 19562 7098
rect 19574 7046 19626 7098
rect 19638 7046 19690 7098
rect 38382 7046 38434 7098
rect 38446 7046 38498 7098
rect 38510 7046 38562 7098
rect 38574 7046 38626 7098
rect 38638 7046 38690 7098
rect 57382 7046 57434 7098
rect 57446 7046 57498 7098
rect 57510 7046 57562 7098
rect 57574 7046 57626 7098
rect 57638 7046 57690 7098
rect 76382 7046 76434 7098
rect 76446 7046 76498 7098
rect 76510 7046 76562 7098
rect 76574 7046 76626 7098
rect 76638 7046 76690 7098
rect 87834 7046 87886 7098
rect 87898 7046 87950 7098
rect 87962 7046 88014 7098
rect 88026 7046 88078 7098
rect 88090 7046 88142 7098
rect 18722 6502 18774 6554
rect 18786 6502 18838 6554
rect 18850 6502 18902 6554
rect 18914 6502 18966 6554
rect 18978 6502 19030 6554
rect 37722 6502 37774 6554
rect 37786 6502 37838 6554
rect 37850 6502 37902 6554
rect 37914 6502 37966 6554
rect 37978 6502 38030 6554
rect 56722 6502 56774 6554
rect 56786 6502 56838 6554
rect 56850 6502 56902 6554
rect 56914 6502 56966 6554
rect 56978 6502 57030 6554
rect 75722 6502 75774 6554
rect 75786 6502 75838 6554
rect 75850 6502 75902 6554
rect 75914 6502 75966 6554
rect 75978 6502 76030 6554
rect 19382 5958 19434 6010
rect 19446 5958 19498 6010
rect 19510 5958 19562 6010
rect 19574 5958 19626 6010
rect 19638 5958 19690 6010
rect 38382 5958 38434 6010
rect 38446 5958 38498 6010
rect 38510 5958 38562 6010
rect 38574 5958 38626 6010
rect 38638 5958 38690 6010
rect 57382 5958 57434 6010
rect 57446 5958 57498 6010
rect 57510 5958 57562 6010
rect 57574 5958 57626 6010
rect 57638 5958 57690 6010
rect 76382 5958 76434 6010
rect 76446 5958 76498 6010
rect 76510 5958 76562 6010
rect 76574 5958 76626 6010
rect 76638 5958 76690 6010
rect 82120 5688 82172 5740
rect 82396 5620 82448 5672
rect 18722 5414 18774 5466
rect 18786 5414 18838 5466
rect 18850 5414 18902 5466
rect 18914 5414 18966 5466
rect 18978 5414 19030 5466
rect 37722 5414 37774 5466
rect 37786 5414 37838 5466
rect 37850 5414 37902 5466
rect 37914 5414 37966 5466
rect 37978 5414 38030 5466
rect 56722 5414 56774 5466
rect 56786 5414 56838 5466
rect 56850 5414 56902 5466
rect 56914 5414 56966 5466
rect 56978 5414 57030 5466
rect 75722 5414 75774 5466
rect 75786 5414 75838 5466
rect 75850 5414 75902 5466
rect 75914 5414 75966 5466
rect 75978 5414 76030 5466
rect 12660 5280 12712 5332
rect 14684 5323 14736 5332
rect 14684 5289 14693 5323
rect 14693 5289 14727 5323
rect 14727 5289 14736 5323
rect 14684 5280 14736 5289
rect 30968 5280 31020 5332
rect 33176 5280 33228 5332
rect 34280 5280 34332 5332
rect 35384 5323 35436 5332
rect 35384 5289 35402 5323
rect 35402 5289 35436 5323
rect 35384 5280 35436 5289
rect 36488 5280 36540 5332
rect 37592 5280 37644 5332
rect 38788 5280 38840 5332
rect 40904 5280 40956 5332
rect 44216 5280 44268 5332
rect 45320 5280 45372 5332
rect 68044 5280 68096 5332
rect 69332 5280 69384 5332
rect 70160 5323 70212 5332
rect 70160 5289 70178 5323
rect 70178 5289 70212 5323
rect 70160 5280 70212 5289
rect 72460 5280 72512 5332
rect 73564 5280 73616 5332
rect 74760 5323 74812 5332
rect 74760 5289 74778 5323
rect 74778 5289 74812 5323
rect 74760 5280 74812 5289
rect 75588 5280 75640 5332
rect 76876 5280 76928 5332
rect 77888 5323 77940 5332
rect 77888 5289 77906 5323
rect 77906 5289 77940 5323
rect 77888 5280 77940 5289
rect 81660 5280 81712 5332
rect 32072 5212 32124 5264
rect 39800 5212 39852 5264
rect 42008 5212 42060 5264
rect 43112 5212 43164 5264
rect 71356 5212 71408 5264
rect 79084 5212 79136 5264
rect 80280 5212 80332 5264
rect 12568 5076 12620 5128
rect 13856 5076 13908 5128
rect 14500 5076 14552 5128
rect 15512 5144 15564 5196
rect 15420 5076 15472 5128
rect 16616 5110 16668 5162
rect 17720 5110 17772 5162
rect 19100 5153 19152 5162
rect 19100 5119 19109 5153
rect 19109 5119 19143 5153
rect 19143 5119 19152 5153
rect 19100 5110 19152 5119
rect 19928 5153 19980 5162
rect 19928 5119 19968 5153
rect 19968 5119 19980 5153
rect 19928 5110 19980 5119
rect 21032 5153 21084 5162
rect 21032 5119 21041 5153
rect 21041 5119 21075 5153
rect 21075 5119 21084 5153
rect 21032 5110 21084 5119
rect 22136 5110 22188 5162
rect 23332 5110 23384 5162
rect 24344 5110 24396 5162
rect 25448 5110 25500 5162
rect 26552 5110 26604 5162
rect 27656 5153 27708 5162
rect 27656 5119 27696 5153
rect 27696 5119 27708 5153
rect 27656 5110 27708 5119
rect 28760 5153 28812 5162
rect 28760 5119 28769 5153
rect 28769 5119 28803 5153
rect 28803 5119 28812 5153
rect 28760 5110 28812 5119
rect 29864 5110 29916 5162
rect 31244 5104 31296 5156
rect 31888 5110 31940 5162
rect 33176 5076 33228 5128
rect 34464 5084 34516 5136
rect 35108 5110 35160 5162
rect 36396 5110 36448 5162
rect 37684 5104 37736 5156
rect 38972 5104 39024 5156
rect 39616 5110 39668 5162
rect 44124 5144 44176 5196
rect 45412 5144 45464 5196
rect 40904 5076 40956 5128
rect 42192 5076 42244 5128
rect 42836 5076 42888 5128
rect 52588 5153 52640 5162
rect 52588 5119 52597 5153
rect 52597 5119 52631 5153
rect 52631 5119 52640 5153
rect 52588 5110 52640 5119
rect 53692 5110 53744 5162
rect 54796 5153 54848 5162
rect 54796 5119 54815 5153
rect 54815 5119 54848 5153
rect 54796 5110 54848 5119
rect 55808 5153 55860 5162
rect 55808 5119 55817 5153
rect 55817 5119 55851 5153
rect 55851 5119 55860 5153
rect 55808 5110 55860 5119
rect 57096 5153 57148 5162
rect 57096 5119 57105 5153
rect 57105 5119 57139 5153
rect 57139 5119 57148 5153
rect 57096 5110 57148 5119
rect 58200 5110 58252 5162
rect 59120 5153 59172 5162
rect 59120 5119 59129 5153
rect 59129 5119 59163 5153
rect 59163 5119 59172 5153
rect 59120 5110 59172 5119
rect 60316 5153 60368 5162
rect 60316 5119 60325 5153
rect 60325 5119 60359 5153
rect 60359 5119 60368 5153
rect 60316 5110 60368 5119
rect 61420 5110 61472 5162
rect 62524 5153 62576 5162
rect 62524 5119 62543 5153
rect 62543 5119 62576 5153
rect 62524 5110 62576 5119
rect 63536 5153 63588 5162
rect 63536 5119 63545 5153
rect 63545 5119 63579 5153
rect 63579 5119 63588 5153
rect 63536 5110 63588 5119
rect 64732 5110 64784 5162
rect 65836 5110 65888 5162
rect 66848 5153 66900 5162
rect 66848 5119 66857 5153
rect 66857 5119 66891 5153
rect 66891 5119 66900 5153
rect 66848 5110 66900 5119
rect 67952 5084 68004 5136
rect 69240 5076 69292 5128
rect 69884 5110 69936 5162
rect 71172 5110 71224 5162
rect 72460 5104 72512 5156
rect 73748 5104 73800 5156
rect 74392 5110 74444 5162
rect 75680 5084 75732 5136
rect 76968 5076 77020 5128
rect 77612 5110 77664 5162
rect 81476 5144 81528 5196
rect 78900 5076 78952 5128
rect 80188 5076 80240 5128
rect 15788 5008 15840 5060
rect 16432 5008 16484 5060
rect 17720 5008 17772 5060
rect 19008 5008 19060 5060
rect 19744 5008 19796 5060
rect 20940 5008 20992 5060
rect 22228 5008 22280 5060
rect 23516 5008 23568 5060
rect 24160 5008 24212 5060
rect 25448 5008 25500 5060
rect 26736 5008 26788 5060
rect 27380 5008 27432 5060
rect 28668 5008 28720 5060
rect 29956 5008 30008 5060
rect 52496 5008 52548 5060
rect 53784 5008 53836 5060
rect 54428 5008 54480 5060
rect 55716 5008 55768 5060
rect 57004 5008 57056 5060
rect 58292 5008 58344 5060
rect 58936 5008 58988 5060
rect 60224 5008 60276 5060
rect 61512 5008 61564 5060
rect 62156 5008 62208 5060
rect 63444 5008 63496 5060
rect 64732 5008 64784 5060
rect 66020 5008 66072 5060
rect 66664 5008 66716 5060
rect 19382 4870 19434 4922
rect 19446 4870 19498 4922
rect 19510 4870 19562 4922
rect 19574 4870 19626 4922
rect 19638 4870 19690 4922
rect 38382 4870 38434 4922
rect 38446 4870 38498 4922
rect 38510 4870 38562 4922
rect 38574 4870 38626 4922
rect 38638 4870 38690 4922
rect 57382 4870 57434 4922
rect 57446 4870 57498 4922
rect 57510 4870 57562 4922
rect 57574 4870 57626 4922
rect 57638 4870 57690 4922
rect 76382 4870 76434 4922
rect 76446 4870 76498 4922
rect 76510 4870 76562 4922
rect 76574 4870 76626 4922
rect 76638 4870 76690 4922
<< metal2 >>
rect 15786 91800 15842 92600
rect 16430 91800 16486 92600
rect 17718 91800 17774 92600
rect 19006 91800 19062 92600
rect 19650 91800 19706 92600
rect 20938 91800 20994 92600
rect 22226 91800 22282 92600
rect 23514 91800 23570 92600
rect 24158 91800 24214 92600
rect 25446 91800 25502 92600
rect 26734 91800 26790 92600
rect 27378 91800 27434 92600
rect 28666 91800 28722 92600
rect 29954 91800 30010 92600
rect 31242 91800 31298 92600
rect 31886 91800 31942 92600
rect 33174 91800 33230 92600
rect 34462 91800 34518 92600
rect 35106 91800 35162 92600
rect 36394 91800 36450 92600
rect 37682 91800 37738 92600
rect 38970 91800 39026 92600
rect 39614 91800 39670 92600
rect 40902 91800 40958 92600
rect 42190 91800 42246 92600
rect 42834 91800 42890 92600
rect 44122 91800 44178 92600
rect 45410 91800 45466 92600
rect 46698 91800 46754 92600
rect 47986 91800 48042 92600
rect 48630 91800 48686 92600
rect 49918 91800 49974 92600
rect 52494 91800 52550 92600
rect 53782 91800 53838 92600
rect 54426 91800 54482 92600
rect 55714 91800 55770 92600
rect 56358 91800 56414 92600
rect 57002 91800 57058 92600
rect 57646 91800 57702 92600
rect 58290 91800 58346 92600
rect 58934 91800 58990 92600
rect 60222 91800 60278 92600
rect 61510 91800 61566 92600
rect 62154 91800 62210 92600
rect 63442 91800 63498 92600
rect 64730 91800 64786 92600
rect 66018 91800 66074 92600
rect 66662 91800 66718 92600
rect 67950 91800 68006 92600
rect 69238 91800 69294 92600
rect 69882 91800 69938 92600
rect 71170 91800 71226 92600
rect 72458 91800 72514 92600
rect 73746 91800 73802 92600
rect 74390 91800 74446 92600
rect 75678 91800 75734 92600
rect 76966 91800 77022 92600
rect 77610 91800 77666 92600
rect 78898 91800 78954 92600
rect 80186 91800 80242 92600
rect 81474 91800 81530 92600
rect 82118 91800 82174 92600
rect 15800 88944 15828 91800
rect 16444 88944 16472 91800
rect 15788 88938 15840 88944
rect 15788 88880 15840 88886
rect 16432 88938 16484 88944
rect 17732 88910 17760 91800
rect 19020 90354 19048 91800
rect 19020 90326 19140 90354
rect 18722 89244 19030 89253
rect 18722 89242 18728 89244
rect 18784 89242 18808 89244
rect 18864 89242 18888 89244
rect 18944 89242 18968 89244
rect 19024 89242 19030 89244
rect 18784 89190 18786 89242
rect 18966 89190 18968 89242
rect 18722 89188 18728 89190
rect 18784 89188 18808 89190
rect 18864 89188 18888 89190
rect 18944 89188 18968 89190
rect 19024 89188 19030 89190
rect 18722 89179 19030 89188
rect 19112 88944 19140 90326
rect 19664 88944 19692 91800
rect 19100 88938 19152 88944
rect 16432 88880 16484 88886
rect 17720 88904 17772 88910
rect 19100 88880 19152 88886
rect 19652 88938 19704 88944
rect 20952 88910 20980 91800
rect 22240 88944 22268 91800
rect 23528 88944 23556 91800
rect 24172 88944 24200 91800
rect 25460 88978 25488 91800
rect 25448 88972 25500 88978
rect 22228 88938 22280 88944
rect 19652 88880 19704 88886
rect 20940 88904 20992 88910
rect 17720 88846 17772 88852
rect 22228 88880 22280 88886
rect 23516 88938 23568 88944
rect 23516 88880 23568 88886
rect 24160 88938 24212 88944
rect 25448 88914 25500 88920
rect 26748 88910 26776 91800
rect 27392 88910 27420 91800
rect 28680 88944 28708 91800
rect 29968 88944 29996 91800
rect 31256 89114 31284 91800
rect 31900 89114 31928 91800
rect 33188 89114 33216 91800
rect 34476 89114 34504 91800
rect 35120 89114 35148 91800
rect 36408 89114 36436 91800
rect 37696 89402 37724 91800
rect 37604 89374 37724 89402
rect 37604 89114 37632 89374
rect 37722 89244 38030 89253
rect 37722 89242 37728 89244
rect 37784 89242 37808 89244
rect 37864 89242 37888 89244
rect 37944 89242 37968 89244
rect 38024 89242 38030 89244
rect 37784 89190 37786 89242
rect 37966 89190 37968 89242
rect 37722 89188 37728 89190
rect 37784 89188 37808 89190
rect 37864 89188 37888 89190
rect 37944 89188 37968 89190
rect 38024 89188 38030 89190
rect 37722 89179 38030 89188
rect 38984 89114 39012 91800
rect 39628 89114 39656 91800
rect 40916 89114 40944 91800
rect 42204 89114 42232 91800
rect 42848 89114 42876 91800
rect 44136 89114 44164 91800
rect 45424 89114 45452 91800
rect 46712 89114 46740 91800
rect 31244 89108 31296 89114
rect 31244 89050 31296 89056
rect 31888 89108 31940 89114
rect 31888 89050 31940 89056
rect 33176 89108 33228 89114
rect 33176 89050 33228 89056
rect 34464 89108 34516 89114
rect 34464 89050 34516 89056
rect 35108 89108 35160 89114
rect 35108 89050 35160 89056
rect 36396 89108 36448 89114
rect 36396 89050 36448 89056
rect 37592 89108 37644 89114
rect 37592 89050 37644 89056
rect 38972 89108 39024 89114
rect 38972 89050 39024 89056
rect 39616 89108 39668 89114
rect 39616 89050 39668 89056
rect 40904 89108 40956 89114
rect 40904 89050 40956 89056
rect 42192 89108 42244 89114
rect 42192 89050 42244 89056
rect 42836 89108 42888 89114
rect 42836 89050 42888 89056
rect 44124 89108 44176 89114
rect 44124 89050 44176 89056
rect 45412 89108 45464 89114
rect 45412 89050 45464 89056
rect 46700 89108 46752 89114
rect 46700 89050 46752 89056
rect 28668 88938 28720 88944
rect 24160 88880 24212 88886
rect 24344 88904 24396 88910
rect 20940 88846 20992 88852
rect 24344 88846 24396 88852
rect 26736 88904 26788 88910
rect 26736 88846 26788 88852
rect 27380 88904 27432 88910
rect 28668 88880 28720 88886
rect 29956 88938 30008 88944
rect 32072 88938 32124 88944
rect 29956 88880 30008 88886
rect 30968 88904 31020 88910
rect 27380 88846 27432 88852
rect 32072 88880 32124 88886
rect 33176 88938 33228 88944
rect 33176 88880 33228 88886
rect 34280 88938 34332 88944
rect 34280 88880 34332 88886
rect 35384 88938 35436 88944
rect 35384 88880 35436 88886
rect 36488 88938 36540 88944
rect 36488 88880 36540 88886
rect 37592 88938 37644 88944
rect 37592 88880 37644 88886
rect 38788 88938 38840 88944
rect 38788 88880 38840 88886
rect 39800 88938 39852 88944
rect 39800 88880 39852 88886
rect 40904 88938 40956 88944
rect 40904 88880 40956 88886
rect 42008 88938 42060 88944
rect 42008 88880 42060 88886
rect 43112 88938 43164 88944
rect 43112 88880 43164 88886
rect 44216 88938 44268 88944
rect 44216 88880 44268 88886
rect 45320 88938 45372 88944
rect 45320 88880 45372 88886
rect 30968 88846 31020 88852
rect 15512 88836 15564 88842
rect 15512 88778 15564 88784
rect 16708 88836 16760 88842
rect 16708 88778 16760 88784
rect 17812 88836 17864 88842
rect 17812 88778 17864 88784
rect 18640 88836 18692 88842
rect 18640 88778 18692 88784
rect 19928 88836 19980 88842
rect 19928 88778 19980 88784
rect 21032 88836 21084 88842
rect 21032 88778 21084 88784
rect 22136 88836 22188 88842
rect 22136 88778 22188 88784
rect 23240 88836 23292 88842
rect 23240 88778 23292 88784
rect 5954 87068 6262 87077
rect 5954 87066 5960 87068
rect 6016 87066 6040 87068
rect 6096 87066 6120 87068
rect 6176 87066 6200 87068
rect 6256 87066 6262 87068
rect 6016 87014 6018 87066
rect 6198 87014 6200 87066
rect 5954 87012 5960 87014
rect 6016 87012 6040 87014
rect 6096 87012 6120 87014
rect 6176 87012 6200 87014
rect 6256 87012 6262 87014
rect 5954 87003 6262 87012
rect 7600 86728 7652 86734
rect 7600 86670 7652 86676
rect 6690 86524 6998 86533
rect 6690 86522 6696 86524
rect 6752 86522 6776 86524
rect 6832 86522 6856 86524
rect 6912 86522 6936 86524
rect 6992 86522 6998 86524
rect 6752 86470 6754 86522
rect 6934 86470 6936 86522
rect 6690 86468 6696 86470
rect 6752 86468 6776 86470
rect 6832 86468 6856 86470
rect 6912 86468 6936 86470
rect 6992 86468 6998 86470
rect 6690 86459 6998 86468
rect 5954 85980 6262 85989
rect 5954 85978 5960 85980
rect 6016 85978 6040 85980
rect 6096 85978 6120 85980
rect 6176 85978 6200 85980
rect 6256 85978 6262 85980
rect 6016 85926 6018 85978
rect 6198 85926 6200 85978
rect 5954 85924 5960 85926
rect 6016 85924 6040 85926
rect 6096 85924 6120 85926
rect 6176 85924 6200 85926
rect 6256 85924 6262 85926
rect 5954 85915 6262 85924
rect 6690 85436 6998 85445
rect 6690 85434 6696 85436
rect 6752 85434 6776 85436
rect 6832 85434 6856 85436
rect 6912 85434 6936 85436
rect 6992 85434 6998 85436
rect 6752 85382 6754 85434
rect 6934 85382 6936 85434
rect 6690 85380 6696 85382
rect 6752 85380 6776 85382
rect 6832 85380 6856 85382
rect 6912 85380 6936 85382
rect 6992 85380 6998 85382
rect 6690 85371 6998 85380
rect 5954 84892 6262 84901
rect 5954 84890 5960 84892
rect 6016 84890 6040 84892
rect 6096 84890 6120 84892
rect 6176 84890 6200 84892
rect 6256 84890 6262 84892
rect 6016 84838 6018 84890
rect 6198 84838 6200 84890
rect 5954 84836 5960 84838
rect 6016 84836 6040 84838
rect 6096 84836 6120 84838
rect 6176 84836 6200 84838
rect 6256 84836 6262 84838
rect 5954 84827 6262 84836
rect 6690 84348 6998 84357
rect 6690 84346 6696 84348
rect 6752 84346 6776 84348
rect 6832 84346 6856 84348
rect 6912 84346 6936 84348
rect 6992 84346 6998 84348
rect 6752 84294 6754 84346
rect 6934 84294 6936 84346
rect 6690 84292 6696 84294
rect 6752 84292 6776 84294
rect 6832 84292 6856 84294
rect 6912 84292 6936 84294
rect 6992 84292 6998 84294
rect 6690 84283 6998 84292
rect 5954 83804 6262 83813
rect 5954 83802 5960 83804
rect 6016 83802 6040 83804
rect 6096 83802 6120 83804
rect 6176 83802 6200 83804
rect 6256 83802 6262 83804
rect 6016 83750 6018 83802
rect 6198 83750 6200 83802
rect 5954 83748 5960 83750
rect 6016 83748 6040 83750
rect 6096 83748 6120 83750
rect 6176 83748 6200 83750
rect 6256 83748 6262 83750
rect 5954 83739 6262 83748
rect 6690 83260 6998 83269
rect 6690 83258 6696 83260
rect 6752 83258 6776 83260
rect 6832 83258 6856 83260
rect 6912 83258 6936 83260
rect 6992 83258 6998 83260
rect 6752 83206 6754 83258
rect 6934 83206 6936 83258
rect 6690 83204 6696 83206
rect 6752 83204 6776 83206
rect 6832 83204 6856 83206
rect 6912 83204 6936 83206
rect 6992 83204 6998 83206
rect 6690 83195 6998 83204
rect 5954 82716 6262 82725
rect 5954 82714 5960 82716
rect 6016 82714 6040 82716
rect 6096 82714 6120 82716
rect 6176 82714 6200 82716
rect 6256 82714 6262 82716
rect 6016 82662 6018 82714
rect 6198 82662 6200 82714
rect 5954 82660 5960 82662
rect 6016 82660 6040 82662
rect 6096 82660 6120 82662
rect 6176 82660 6200 82662
rect 6256 82660 6262 82662
rect 5954 82651 6262 82660
rect 6690 82172 6998 82181
rect 6690 82170 6696 82172
rect 6752 82170 6776 82172
rect 6832 82170 6856 82172
rect 6912 82170 6936 82172
rect 6992 82170 6998 82172
rect 6752 82118 6754 82170
rect 6934 82118 6936 82170
rect 6690 82116 6696 82118
rect 6752 82116 6776 82118
rect 6832 82116 6856 82118
rect 6912 82116 6936 82118
rect 6992 82116 6998 82118
rect 6690 82107 6998 82116
rect 5954 81628 6262 81637
rect 5954 81626 5960 81628
rect 6016 81626 6040 81628
rect 6096 81626 6120 81628
rect 6176 81626 6200 81628
rect 6256 81626 6262 81628
rect 6016 81574 6018 81626
rect 6198 81574 6200 81626
rect 5954 81572 5960 81574
rect 6016 81572 6040 81574
rect 6096 81572 6120 81574
rect 6176 81572 6200 81574
rect 6256 81572 6262 81574
rect 5954 81563 6262 81572
rect 6690 81084 6998 81093
rect 6690 81082 6696 81084
rect 6752 81082 6776 81084
rect 6832 81082 6856 81084
rect 6912 81082 6936 81084
rect 6992 81082 6998 81084
rect 6752 81030 6754 81082
rect 6934 81030 6936 81082
rect 6690 81028 6696 81030
rect 6752 81028 6776 81030
rect 6832 81028 6856 81030
rect 6912 81028 6936 81030
rect 6992 81028 6998 81030
rect 6690 81019 6998 81028
rect 7140 80812 7192 80818
rect 7140 80754 7192 80760
rect 2908 80676 2960 80682
rect 2908 80618 2960 80624
rect 2920 80585 2948 80618
rect 2906 80576 2962 80585
rect 2906 80511 2962 80520
rect 5954 80540 6262 80549
rect 5954 80538 5960 80540
rect 6016 80538 6040 80540
rect 6096 80538 6120 80540
rect 6176 80538 6200 80540
rect 6256 80538 6262 80540
rect 6016 80486 6018 80538
rect 6198 80486 6200 80538
rect 5954 80484 5960 80486
rect 6016 80484 6040 80486
rect 6096 80484 6120 80486
rect 6176 80484 6200 80486
rect 6256 80484 6262 80486
rect 5954 80475 6262 80484
rect 7152 80449 7180 80754
rect 7138 80440 7194 80449
rect 7138 80375 7194 80384
rect 6690 79996 6998 80005
rect 6690 79994 6696 79996
rect 6752 79994 6776 79996
rect 6832 79994 6856 79996
rect 6912 79994 6936 79996
rect 6992 79994 6998 79996
rect 6752 79942 6754 79994
rect 6934 79942 6936 79994
rect 6690 79940 6696 79942
rect 6752 79940 6776 79942
rect 6832 79940 6856 79942
rect 6912 79940 6936 79942
rect 6992 79940 6998 79942
rect 6690 79931 6998 79940
rect 7140 79724 7192 79730
rect 7140 79666 7192 79672
rect 2724 79588 2776 79594
rect 2724 79530 2776 79536
rect 2736 79225 2764 79530
rect 5954 79452 6262 79461
rect 5954 79450 5960 79452
rect 6016 79450 6040 79452
rect 6096 79450 6120 79452
rect 6176 79450 6200 79452
rect 6256 79450 6262 79452
rect 6016 79398 6018 79450
rect 6198 79398 6200 79450
rect 5954 79396 5960 79398
rect 6016 79396 6040 79398
rect 6096 79396 6120 79398
rect 6176 79396 6200 79398
rect 6256 79396 6262 79398
rect 5954 79387 6262 79396
rect 7152 79361 7180 79666
rect 7138 79352 7194 79361
rect 7138 79287 7194 79296
rect 2722 79216 2778 79225
rect 2722 79151 2778 79160
rect 6690 78908 6998 78917
rect 6690 78906 6696 78908
rect 6752 78906 6776 78908
rect 6832 78906 6856 78908
rect 6912 78906 6936 78908
rect 6992 78906 6998 78908
rect 6752 78854 6754 78906
rect 6934 78854 6936 78906
rect 6690 78852 6696 78854
rect 6752 78852 6776 78854
rect 6832 78852 6856 78854
rect 6912 78852 6936 78854
rect 6992 78852 6998 78854
rect 6690 78843 6998 78852
rect 7140 78636 7192 78642
rect 7140 78578 7192 78584
rect 2906 78536 2962 78545
rect 2906 78471 2908 78480
rect 2960 78471 2962 78480
rect 2908 78442 2960 78448
rect 5954 78364 6262 78373
rect 5954 78362 5960 78364
rect 6016 78362 6040 78364
rect 6096 78362 6120 78364
rect 6176 78362 6200 78364
rect 6256 78362 6262 78364
rect 6016 78310 6018 78362
rect 6198 78310 6200 78362
rect 5954 78308 5960 78310
rect 6016 78308 6040 78310
rect 6096 78308 6120 78310
rect 6176 78308 6200 78310
rect 6256 78308 6262 78310
rect 5954 78299 6262 78308
rect 7152 78273 7180 78578
rect 7138 78264 7194 78273
rect 7138 78199 7194 78208
rect 6690 77820 6998 77829
rect 6690 77818 6696 77820
rect 6752 77818 6776 77820
rect 6832 77818 6856 77820
rect 6912 77818 6936 77820
rect 6992 77818 6998 77820
rect 6752 77766 6754 77818
rect 6934 77766 6936 77818
rect 6690 77764 6696 77766
rect 6752 77764 6776 77766
rect 6832 77764 6856 77766
rect 6912 77764 6936 77766
rect 6992 77764 6998 77766
rect 6690 77755 6998 77764
rect 4380 77684 4432 77690
rect 4380 77626 4432 77632
rect 4392 77185 4420 77626
rect 5668 77582 5720 77588
rect 5668 77524 5720 77530
rect 4378 77176 4434 77185
rect 4378 77111 4434 77120
rect 5680 77049 5708 77524
rect 5954 77276 6262 77285
rect 5954 77274 5960 77276
rect 6016 77274 6040 77276
rect 6096 77274 6120 77276
rect 6176 77274 6200 77276
rect 6256 77274 6262 77276
rect 6016 77222 6018 77274
rect 6198 77222 6200 77274
rect 5954 77220 5960 77222
rect 6016 77220 6040 77222
rect 6096 77220 6120 77222
rect 6176 77220 6200 77222
rect 6256 77220 6262 77222
rect 5954 77211 6262 77220
rect 5666 77040 5722 77049
rect 5666 76975 5722 76984
rect 6690 76732 6998 76741
rect 6690 76730 6696 76732
rect 6752 76730 6776 76732
rect 6832 76730 6856 76732
rect 6912 76730 6936 76732
rect 6992 76730 6998 76732
rect 6752 76678 6754 76730
rect 6934 76678 6936 76730
rect 6690 76676 6696 76678
rect 6752 76676 6776 76678
rect 6832 76676 6856 76678
rect 6912 76676 6936 76678
rect 6992 76676 6998 76678
rect 6690 76667 6998 76676
rect 5954 76188 6262 76197
rect 5954 76186 5960 76188
rect 6016 76186 6040 76188
rect 6096 76186 6120 76188
rect 6176 76186 6200 76188
rect 6256 76186 6262 76188
rect 6016 76134 6018 76186
rect 6198 76134 6200 76186
rect 5954 76132 5960 76134
rect 6016 76132 6040 76134
rect 6096 76132 6120 76134
rect 6176 76132 6200 76134
rect 6256 76132 6262 76134
rect 5954 76123 6262 76132
rect 7138 76088 7194 76097
rect 7138 76023 7194 76032
rect 7152 75922 7180 76023
rect 7140 75916 7192 75922
rect 7140 75858 7192 75864
rect 2906 75816 2962 75825
rect 2906 75751 2908 75760
rect 2960 75751 2962 75760
rect 2908 75722 2960 75728
rect 6690 75644 6998 75653
rect 6690 75642 6696 75644
rect 6752 75642 6776 75644
rect 6832 75642 6856 75644
rect 6912 75642 6936 75644
rect 6992 75642 6998 75644
rect 6752 75590 6754 75642
rect 6934 75590 6936 75642
rect 6690 75588 6696 75590
rect 6752 75588 6776 75590
rect 6832 75588 6856 75590
rect 6912 75588 6936 75590
rect 6992 75588 6998 75590
rect 6690 75579 6998 75588
rect 7140 75372 7192 75378
rect 7140 75314 7192 75320
rect 2908 75236 2960 75242
rect 2908 75178 2960 75184
rect 2920 75145 2948 75178
rect 2906 75136 2962 75145
rect 2906 75071 2962 75080
rect 5954 75100 6262 75109
rect 5954 75098 5960 75100
rect 6016 75098 6040 75100
rect 6096 75098 6120 75100
rect 6176 75098 6200 75100
rect 6256 75098 6262 75100
rect 6016 75046 6018 75098
rect 6198 75046 6200 75098
rect 5954 75044 5960 75046
rect 6016 75044 6040 75046
rect 6096 75044 6120 75046
rect 6176 75044 6200 75046
rect 6256 75044 6262 75046
rect 5954 75035 6262 75044
rect 7152 75009 7180 75314
rect 7138 75000 7194 75009
rect 7138 74935 7194 74944
rect 6690 74556 6998 74565
rect 6690 74554 6696 74556
rect 6752 74554 6776 74556
rect 6832 74554 6856 74556
rect 6912 74554 6936 74556
rect 6992 74554 6998 74556
rect 6752 74502 6754 74554
rect 6934 74502 6936 74554
rect 6690 74500 6696 74502
rect 6752 74500 6776 74502
rect 6832 74500 6856 74502
rect 6912 74500 6936 74502
rect 6992 74500 6998 74502
rect 6690 74491 6998 74500
rect 7140 74284 7192 74290
rect 7140 74226 7192 74232
rect 2908 74148 2960 74154
rect 2908 74090 2960 74096
rect 2920 73785 2948 74090
rect 5954 74012 6262 74021
rect 5954 74010 5960 74012
rect 6016 74010 6040 74012
rect 6096 74010 6120 74012
rect 6176 74010 6200 74012
rect 6256 74010 6262 74012
rect 6016 73958 6018 74010
rect 6198 73958 6200 74010
rect 5954 73956 5960 73958
rect 6016 73956 6040 73958
rect 6096 73956 6120 73958
rect 6176 73956 6200 73958
rect 6256 73956 6262 73958
rect 5954 73947 6262 73956
rect 7152 73921 7180 74226
rect 7138 73912 7194 73921
rect 7138 73847 7194 73856
rect 2906 73776 2962 73785
rect 2906 73711 2962 73720
rect 6690 73468 6998 73477
rect 6690 73466 6696 73468
rect 6752 73466 6776 73468
rect 6832 73466 6856 73468
rect 6912 73466 6936 73468
rect 6992 73466 6998 73468
rect 6752 73414 6754 73466
rect 6934 73414 6936 73466
rect 6690 73412 6696 73414
rect 6752 73412 6776 73414
rect 6832 73412 6856 73414
rect 6912 73412 6936 73414
rect 6992 73412 6998 73414
rect 6690 73403 6998 73412
rect 7140 73196 7192 73202
rect 7140 73138 7192 73144
rect 2906 73096 2962 73105
rect 2906 73031 2908 73040
rect 2960 73031 2962 73040
rect 2908 73002 2960 73008
rect 5954 72924 6262 72933
rect 5954 72922 5960 72924
rect 6016 72922 6040 72924
rect 6096 72922 6120 72924
rect 6176 72922 6200 72924
rect 6256 72922 6262 72924
rect 6016 72870 6018 72922
rect 6198 72870 6200 72922
rect 5954 72868 5960 72870
rect 6016 72868 6040 72870
rect 6096 72868 6120 72870
rect 6176 72868 6200 72870
rect 6256 72868 6262 72870
rect 5954 72859 6262 72868
rect 7152 72833 7180 73138
rect 7138 72824 7194 72833
rect 7138 72759 7194 72768
rect 6690 72380 6998 72389
rect 6690 72378 6696 72380
rect 6752 72378 6776 72380
rect 6832 72378 6856 72380
rect 6912 72378 6936 72380
rect 6992 72378 6998 72380
rect 6752 72326 6754 72378
rect 6934 72326 6936 72378
rect 6690 72324 6696 72326
rect 6752 72324 6776 72326
rect 6832 72324 6856 72326
rect 6912 72324 6936 72326
rect 6992 72324 6998 72326
rect 6690 72315 6998 72324
rect 5668 72142 5720 72148
rect 5668 72084 5720 72090
rect 4380 72040 4432 72046
rect 4380 71982 4432 71988
rect 4392 71745 4420 71982
rect 4378 71736 4434 71745
rect 4378 71671 4434 71680
rect 5680 71609 5708 72084
rect 5954 71836 6262 71845
rect 5954 71834 5960 71836
rect 6016 71834 6040 71836
rect 6096 71834 6120 71836
rect 6176 71834 6200 71836
rect 6256 71834 6262 71836
rect 6016 71782 6018 71834
rect 6198 71782 6200 71834
rect 5954 71780 5960 71782
rect 6016 71780 6040 71782
rect 6096 71780 6120 71782
rect 6176 71780 6200 71782
rect 6256 71780 6262 71782
rect 5954 71771 6262 71780
rect 5666 71600 5722 71609
rect 5666 71535 5722 71544
rect 6690 71292 6998 71301
rect 6690 71290 6696 71292
rect 6752 71290 6776 71292
rect 6832 71290 6856 71292
rect 6912 71290 6936 71292
rect 6992 71290 6998 71292
rect 6752 71238 6754 71290
rect 6934 71238 6936 71290
rect 6690 71236 6696 71238
rect 6752 71236 6776 71238
rect 6832 71236 6856 71238
rect 6912 71236 6936 71238
rect 6992 71236 6998 71238
rect 6690 71227 6998 71236
rect 5666 70920 5722 70929
rect 5666 70855 5722 70864
rect 5680 70448 5708 70855
rect 5954 70748 6262 70757
rect 5954 70746 5960 70748
rect 6016 70746 6040 70748
rect 6096 70746 6120 70748
rect 6176 70746 6200 70748
rect 6256 70746 6262 70748
rect 6016 70694 6018 70746
rect 6198 70694 6200 70746
rect 5954 70692 5960 70694
rect 6016 70692 6040 70694
rect 6096 70692 6120 70694
rect 6176 70692 6200 70694
rect 6256 70692 6262 70694
rect 5954 70683 6262 70692
rect 5668 70442 5720 70448
rect 2906 70376 2962 70385
rect 5668 70384 5720 70390
rect 2906 70311 2908 70320
rect 2960 70311 2962 70320
rect 2908 70282 2960 70288
rect 6690 70204 6998 70213
rect 6690 70202 6696 70204
rect 6752 70202 6776 70204
rect 6832 70202 6856 70204
rect 6912 70202 6936 70204
rect 6992 70202 6998 70204
rect 6752 70150 6754 70202
rect 6934 70150 6936 70202
rect 6690 70148 6696 70150
rect 6752 70148 6776 70150
rect 6832 70148 6856 70150
rect 6912 70148 6936 70150
rect 6992 70148 6998 70150
rect 6690 70139 6998 70148
rect 7140 69932 7192 69938
rect 7140 69874 7192 69880
rect 2908 69796 2960 69802
rect 2908 69738 2960 69744
rect 2920 69705 2948 69738
rect 2906 69696 2962 69705
rect 2906 69631 2962 69640
rect 5954 69660 6262 69669
rect 5954 69658 5960 69660
rect 6016 69658 6040 69660
rect 6096 69658 6120 69660
rect 6176 69658 6200 69660
rect 6256 69658 6262 69660
rect 6016 69606 6018 69658
rect 6198 69606 6200 69658
rect 5954 69604 5960 69606
rect 6016 69604 6040 69606
rect 6096 69604 6120 69606
rect 6176 69604 6200 69606
rect 6256 69604 6262 69606
rect 5954 69595 6262 69604
rect 7152 69569 7180 69874
rect 7138 69560 7194 69569
rect 7138 69495 7194 69504
rect 6690 69116 6998 69125
rect 6690 69114 6696 69116
rect 6752 69114 6776 69116
rect 6832 69114 6856 69116
rect 6912 69114 6936 69116
rect 6992 69114 6998 69116
rect 6752 69062 6754 69114
rect 6934 69062 6936 69114
rect 6690 69060 6696 69062
rect 6752 69060 6776 69062
rect 6832 69060 6856 69062
rect 6912 69060 6936 69062
rect 6992 69060 6998 69062
rect 6690 69051 6998 69060
rect 7140 68844 7192 68850
rect 7140 68786 7192 68792
rect 2908 68708 2960 68714
rect 2908 68650 2960 68656
rect 2920 68345 2948 68650
rect 5954 68572 6262 68581
rect 5954 68570 5960 68572
rect 6016 68570 6040 68572
rect 6096 68570 6120 68572
rect 6176 68570 6200 68572
rect 6256 68570 6262 68572
rect 6016 68518 6018 68570
rect 6198 68518 6200 68570
rect 5954 68516 5960 68518
rect 6016 68516 6040 68518
rect 6096 68516 6120 68518
rect 6176 68516 6200 68518
rect 6256 68516 6262 68518
rect 5954 68507 6262 68516
rect 7152 68481 7180 68786
rect 7138 68472 7194 68481
rect 7138 68407 7194 68416
rect 2906 68336 2962 68345
rect 2906 68271 2962 68280
rect 6690 68028 6998 68037
rect 6690 68026 6696 68028
rect 6752 68026 6776 68028
rect 6832 68026 6856 68028
rect 6912 68026 6936 68028
rect 6992 68026 6998 68028
rect 6752 67974 6754 68026
rect 6934 67974 6936 68026
rect 6690 67972 6696 67974
rect 6752 67972 6776 67974
rect 6832 67972 6856 67974
rect 6912 67972 6936 67974
rect 6992 67972 6998 67974
rect 6690 67963 6998 67972
rect 7140 67756 7192 67762
rect 7140 67698 7192 67704
rect 2906 67656 2962 67665
rect 2906 67591 2908 67600
rect 2960 67591 2962 67600
rect 2908 67562 2960 67568
rect 5954 67484 6262 67493
rect 5954 67482 5960 67484
rect 6016 67482 6040 67484
rect 6096 67482 6120 67484
rect 6176 67482 6200 67484
rect 6256 67482 6262 67484
rect 6016 67430 6018 67482
rect 6198 67430 6200 67482
rect 5954 67428 5960 67430
rect 6016 67428 6040 67430
rect 6096 67428 6120 67430
rect 6176 67428 6200 67430
rect 6256 67428 6262 67430
rect 5954 67419 6262 67428
rect 7152 67393 7180 67698
rect 7138 67384 7194 67393
rect 7138 67319 7194 67328
rect 6690 66940 6998 66949
rect 6690 66938 6696 66940
rect 6752 66938 6776 66940
rect 6832 66938 6856 66940
rect 6912 66938 6936 66940
rect 6992 66938 6998 66940
rect 6752 66886 6754 66938
rect 6934 66886 6936 66938
rect 6690 66884 6696 66886
rect 6752 66884 6776 66886
rect 6832 66884 6856 66886
rect 6912 66884 6936 66886
rect 6992 66884 6998 66886
rect 6690 66875 6998 66884
rect 5484 66702 5536 66708
rect 5484 66644 5536 66650
rect 4380 66532 4432 66538
rect 4380 66474 4432 66480
rect 4392 66305 4420 66474
rect 4378 66296 4434 66305
rect 4378 66231 4434 66240
rect 5496 66169 5524 66644
rect 5954 66396 6262 66405
rect 5954 66394 5960 66396
rect 6016 66394 6040 66396
rect 6096 66394 6120 66396
rect 6176 66394 6200 66396
rect 6256 66394 6262 66396
rect 6016 66342 6018 66394
rect 6198 66342 6200 66394
rect 5954 66340 5960 66342
rect 6016 66340 6040 66342
rect 6096 66340 6120 66342
rect 6176 66340 6200 66342
rect 6256 66340 6262 66342
rect 5954 66331 6262 66340
rect 5482 66160 5538 66169
rect 5482 66095 5538 66104
rect 6690 65852 6998 65861
rect 6690 65850 6696 65852
rect 6752 65850 6776 65852
rect 6832 65850 6856 65852
rect 6912 65850 6936 65852
rect 6992 65850 6998 65852
rect 6752 65798 6754 65850
rect 6934 65798 6936 65850
rect 6690 65796 6696 65798
rect 6752 65796 6776 65798
rect 6832 65796 6856 65798
rect 6912 65796 6936 65798
rect 6992 65796 6998 65798
rect 6690 65787 6998 65796
rect 5390 65480 5446 65489
rect 5390 65415 5446 65424
rect 5404 65110 5432 65415
rect 5954 65308 6262 65317
rect 5954 65306 5960 65308
rect 6016 65306 6040 65308
rect 6096 65306 6120 65308
rect 6176 65306 6200 65308
rect 6256 65306 6262 65308
rect 6016 65254 6018 65306
rect 6198 65254 6200 65306
rect 5954 65252 5960 65254
rect 6016 65252 6040 65254
rect 6096 65252 6120 65254
rect 6176 65252 6200 65254
rect 6256 65252 6262 65254
rect 5954 65243 6262 65252
rect 5392 65104 5444 65110
rect 5392 65046 5444 65052
rect 2908 64968 2960 64974
rect 2906 64936 2908 64945
rect 2960 64936 2962 64945
rect 2906 64871 2962 64880
rect 6690 64764 6998 64773
rect 6690 64762 6696 64764
rect 6752 64762 6776 64764
rect 6832 64762 6856 64764
rect 6912 64762 6936 64764
rect 6992 64762 6998 64764
rect 6752 64710 6754 64762
rect 6934 64710 6936 64762
rect 6690 64708 6696 64710
rect 6752 64708 6776 64710
rect 6832 64708 6856 64710
rect 6912 64708 6936 64710
rect 6992 64708 6998 64710
rect 6690 64699 6998 64708
rect 2908 64492 2960 64498
rect 2908 64434 2960 64440
rect 2920 64265 2948 64434
rect 7232 64356 7284 64362
rect 7232 64298 7284 64304
rect 2906 64256 2962 64265
rect 2906 64191 2962 64200
rect 5954 64220 6262 64229
rect 5954 64218 5960 64220
rect 6016 64218 6040 64220
rect 6096 64218 6120 64220
rect 6176 64218 6200 64220
rect 6256 64218 6262 64220
rect 6016 64166 6018 64218
rect 6198 64166 6200 64218
rect 5954 64164 5960 64166
rect 6016 64164 6040 64166
rect 6096 64164 6120 64166
rect 6176 64164 6200 64166
rect 6256 64164 6262 64166
rect 5954 64155 6262 64164
rect 7244 64129 7272 64298
rect 7230 64120 7286 64129
rect 7230 64055 7286 64064
rect 6690 63676 6998 63685
rect 6690 63674 6696 63676
rect 6752 63674 6776 63676
rect 6832 63674 6856 63676
rect 6912 63674 6936 63676
rect 6992 63674 6998 63676
rect 6752 63622 6754 63674
rect 6934 63622 6936 63674
rect 6690 63620 6696 63622
rect 6752 63620 6776 63622
rect 6832 63620 6856 63622
rect 6912 63620 6936 63622
rect 6992 63620 6998 63622
rect 6690 63611 6998 63620
rect 2908 63404 2960 63410
rect 2908 63346 2960 63352
rect 2920 62905 2948 63346
rect 7232 63268 7284 63274
rect 7232 63210 7284 63216
rect 5954 63132 6262 63141
rect 5954 63130 5960 63132
rect 6016 63130 6040 63132
rect 6096 63130 6120 63132
rect 6176 63130 6200 63132
rect 6256 63130 6262 63132
rect 6016 63078 6018 63130
rect 6198 63078 6200 63130
rect 5954 63076 5960 63078
rect 6016 63076 6040 63078
rect 6096 63076 6120 63078
rect 6176 63076 6200 63078
rect 6256 63076 6262 63078
rect 5954 63067 6262 63076
rect 7244 63041 7272 63210
rect 7230 63032 7286 63041
rect 7230 62967 7286 62976
rect 2906 62896 2962 62905
rect 2906 62831 2962 62840
rect 6690 62588 6998 62597
rect 6690 62586 6696 62588
rect 6752 62586 6776 62588
rect 6832 62586 6856 62588
rect 6912 62586 6936 62588
rect 6992 62586 6998 62588
rect 6752 62534 6754 62586
rect 6934 62534 6936 62586
rect 6690 62532 6696 62534
rect 6752 62532 6776 62534
rect 6832 62532 6856 62534
rect 6912 62532 6936 62534
rect 6992 62532 6998 62534
rect 6690 62523 6998 62532
rect 5208 62350 5260 62356
rect 5208 62292 5260 62298
rect 5220 62225 5248 62292
rect 5206 62216 5262 62225
rect 5206 62151 5262 62160
rect 5954 62044 6262 62053
rect 5954 62042 5960 62044
rect 6016 62042 6040 62044
rect 6096 62042 6120 62044
rect 6176 62042 6200 62044
rect 6256 62042 6262 62044
rect 6016 61990 6018 62042
rect 6198 61990 6200 62042
rect 5954 61988 5960 61990
rect 6016 61988 6040 61990
rect 6096 61988 6120 61990
rect 6176 61988 6200 61990
rect 6256 61988 6262 61990
rect 5954 61979 6262 61988
rect 6690 61500 6998 61509
rect 6690 61498 6696 61500
rect 6752 61498 6776 61500
rect 6832 61498 6856 61500
rect 6912 61498 6936 61500
rect 6992 61498 6998 61500
rect 6752 61446 6754 61498
rect 6934 61446 6936 61498
rect 6690 61444 6696 61446
rect 6752 61444 6776 61446
rect 6832 61444 6856 61446
rect 6912 61444 6936 61446
rect 6992 61444 6998 61446
rect 6690 61435 6998 61444
rect 5208 61262 5260 61268
rect 5208 61204 5260 61210
rect 5220 60865 5248 61204
rect 5954 60956 6262 60965
rect 5954 60954 5960 60956
rect 6016 60954 6040 60956
rect 6096 60954 6120 60956
rect 6176 60954 6200 60956
rect 6256 60954 6262 60956
rect 6016 60902 6018 60954
rect 6198 60902 6200 60954
rect 5954 60900 5960 60902
rect 6016 60900 6040 60902
rect 6096 60900 6120 60902
rect 6176 60900 6200 60902
rect 6256 60900 6262 60902
rect 5954 60891 6262 60900
rect 5206 60856 5262 60865
rect 5206 60791 5262 60800
rect 6690 60412 6998 60421
rect 6690 60410 6696 60412
rect 6752 60410 6776 60412
rect 6832 60410 6856 60412
rect 6912 60410 6936 60412
rect 6992 60410 6998 60412
rect 6752 60358 6754 60410
rect 6934 60358 6936 60410
rect 6690 60356 6696 60358
rect 6752 60356 6776 60358
rect 6832 60356 6856 60358
rect 6912 60356 6936 60358
rect 6992 60356 6998 60358
rect 6690 60347 6998 60356
rect 5954 59868 6262 59877
rect 5954 59866 5960 59868
rect 6016 59866 6040 59868
rect 6096 59866 6120 59868
rect 6176 59866 6200 59868
rect 6256 59866 6262 59868
rect 6016 59814 6018 59866
rect 6198 59814 6200 59866
rect 5954 59812 5960 59814
rect 6016 59812 6040 59814
rect 6096 59812 6120 59814
rect 6176 59812 6200 59814
rect 6256 59812 6262 59814
rect 5954 59803 6262 59812
rect 5666 59632 5722 59641
rect 5666 59567 5722 59576
rect 5680 59534 5708 59567
rect 2908 59528 2960 59534
rect 2906 59496 2908 59505
rect 5668 59528 5720 59534
rect 2960 59496 2962 59505
rect 5668 59470 5720 59476
rect 2906 59431 2962 59440
rect 6690 59324 6998 59333
rect 6690 59322 6696 59324
rect 6752 59322 6776 59324
rect 6832 59322 6856 59324
rect 6912 59322 6936 59324
rect 6992 59322 6998 59324
rect 6752 59270 6754 59322
rect 6934 59270 6936 59322
rect 6690 59268 6696 59270
rect 6752 59268 6776 59270
rect 6832 59268 6856 59270
rect 6912 59268 6936 59270
rect 6992 59268 6998 59270
rect 6690 59259 6998 59268
rect 2908 59052 2960 59058
rect 2908 58994 2960 59000
rect 2920 58825 2948 58994
rect 7232 58916 7284 58922
rect 7232 58858 7284 58864
rect 2906 58816 2962 58825
rect 2906 58751 2962 58760
rect 5954 58780 6262 58789
rect 5954 58778 5960 58780
rect 6016 58778 6040 58780
rect 6096 58778 6120 58780
rect 6176 58778 6200 58780
rect 6256 58778 6262 58780
rect 6016 58726 6018 58778
rect 6198 58726 6200 58778
rect 5954 58724 5960 58726
rect 6016 58724 6040 58726
rect 6096 58724 6120 58726
rect 6176 58724 6200 58726
rect 6256 58724 6262 58726
rect 5954 58715 6262 58724
rect 7244 58689 7272 58858
rect 7230 58680 7286 58689
rect 7230 58615 7286 58624
rect 6690 58236 6998 58245
rect 6690 58234 6696 58236
rect 6752 58234 6776 58236
rect 6832 58234 6856 58236
rect 6912 58234 6936 58236
rect 6992 58234 6998 58236
rect 6752 58182 6754 58234
rect 6934 58182 6936 58234
rect 6690 58180 6696 58182
rect 6752 58180 6776 58182
rect 6832 58180 6856 58182
rect 6912 58180 6936 58182
rect 6992 58180 6998 58182
rect 6690 58171 6998 58180
rect 2908 57964 2960 57970
rect 2908 57906 2960 57912
rect 2920 57465 2948 57906
rect 7232 57828 7284 57834
rect 7232 57770 7284 57776
rect 5954 57692 6262 57701
rect 5954 57690 5960 57692
rect 6016 57690 6040 57692
rect 6096 57690 6120 57692
rect 6176 57690 6200 57692
rect 6256 57690 6262 57692
rect 6016 57638 6018 57690
rect 6198 57638 6200 57690
rect 5954 57636 5960 57638
rect 6016 57636 6040 57638
rect 6096 57636 6120 57638
rect 6176 57636 6200 57638
rect 6256 57636 6262 57638
rect 5954 57627 6262 57636
rect 7244 57601 7272 57770
rect 7230 57592 7286 57601
rect 7230 57527 7286 57536
rect 2906 57456 2962 57465
rect 2906 57391 2962 57400
rect 6690 57148 6998 57157
rect 6690 57146 6696 57148
rect 6752 57146 6776 57148
rect 6832 57146 6856 57148
rect 6912 57146 6936 57148
rect 6992 57146 6998 57148
rect 6752 57094 6754 57146
rect 6934 57094 6936 57146
rect 6690 57092 6696 57094
rect 6752 57092 6776 57094
rect 6832 57092 6856 57094
rect 6912 57092 6936 57094
rect 6992 57092 6998 57094
rect 6690 57083 6998 57092
rect 4932 56910 4984 56916
rect 4932 56852 4984 56858
rect 5392 56876 5444 56882
rect 4944 56785 4972 56852
rect 5392 56818 5444 56824
rect 4930 56776 4986 56785
rect 4930 56711 4986 56720
rect 5404 56377 5432 56818
rect 5954 56604 6262 56613
rect 5954 56602 5960 56604
rect 6016 56602 6040 56604
rect 6096 56602 6120 56604
rect 6176 56602 6200 56604
rect 6256 56602 6262 56604
rect 6016 56550 6018 56602
rect 6198 56550 6200 56602
rect 5954 56548 5960 56550
rect 6016 56548 6040 56550
rect 6096 56548 6120 56550
rect 6176 56548 6200 56550
rect 6256 56548 6262 56550
rect 5954 56539 6262 56548
rect 5390 56368 5446 56377
rect 5390 56303 5446 56312
rect 6690 56060 6998 56069
rect 6690 56058 6696 56060
rect 6752 56058 6776 56060
rect 6832 56058 6856 56060
rect 6912 56058 6936 56060
rect 6992 56058 6998 56060
rect 6752 56006 6754 56058
rect 6934 56006 6936 56058
rect 6690 56004 6696 56006
rect 6752 56004 6776 56006
rect 6832 56004 6856 56006
rect 6912 56004 6936 56006
rect 6992 56004 6998 56006
rect 6690 55995 6998 56004
rect 5024 55822 5076 55828
rect 5024 55764 5076 55770
rect 5036 55425 5064 55764
rect 5668 55652 5720 55658
rect 5668 55594 5720 55600
rect 5022 55416 5078 55425
rect 5022 55351 5078 55360
rect 5680 55289 5708 55594
rect 5954 55516 6262 55525
rect 5954 55514 5960 55516
rect 6016 55514 6040 55516
rect 6096 55514 6120 55516
rect 6176 55514 6200 55516
rect 6256 55514 6262 55516
rect 6016 55462 6018 55514
rect 6198 55462 6200 55514
rect 5954 55460 5960 55462
rect 6016 55460 6040 55462
rect 6096 55460 6120 55462
rect 6176 55460 6200 55462
rect 6256 55460 6262 55462
rect 5954 55451 6262 55460
rect 5666 55280 5722 55289
rect 5666 55215 5722 55224
rect 2540 55176 2592 55182
rect 2540 55118 2592 55124
rect 2552 54745 2580 55118
rect 6690 54972 6998 54981
rect 6690 54970 6696 54972
rect 6752 54970 6776 54972
rect 6832 54970 6856 54972
rect 6912 54970 6936 54972
rect 6992 54970 6998 54972
rect 6752 54918 6754 54970
rect 6934 54918 6936 54970
rect 6690 54916 6696 54918
rect 6752 54916 6776 54918
rect 6832 54916 6856 54918
rect 6912 54916 6936 54918
rect 6992 54916 6998 54918
rect 6690 54907 6998 54916
rect 7612 54774 7640 86670
rect 8426 84384 8482 84393
rect 8426 84319 8482 84328
rect 14406 84384 14462 84393
rect 15524 84356 15552 88778
rect 16720 85794 16748 88778
rect 17824 85794 17852 88778
rect 16628 85766 16748 85794
rect 17732 85766 17852 85794
rect 16628 84356 16656 85766
rect 17732 84356 17760 85766
rect 18652 84370 18680 88778
rect 19382 88700 19690 88709
rect 19382 88698 19388 88700
rect 19444 88698 19468 88700
rect 19524 88698 19548 88700
rect 19604 88698 19628 88700
rect 19684 88698 19690 88700
rect 19444 88646 19446 88698
rect 19626 88646 19628 88698
rect 19382 88644 19388 88646
rect 19444 88644 19468 88646
rect 19524 88644 19548 88646
rect 19604 88644 19628 88646
rect 19684 88644 19690 88646
rect 19382 88635 19690 88644
rect 18722 88156 19030 88165
rect 18722 88154 18728 88156
rect 18784 88154 18808 88156
rect 18864 88154 18888 88156
rect 18944 88154 18968 88156
rect 19024 88154 19030 88156
rect 18784 88102 18786 88154
rect 18966 88102 18968 88154
rect 18722 88100 18728 88102
rect 18784 88100 18808 88102
rect 18864 88100 18888 88102
rect 18944 88100 18968 88102
rect 19024 88100 19030 88102
rect 18722 88091 19030 88100
rect 19382 87612 19690 87621
rect 19382 87610 19388 87612
rect 19444 87610 19468 87612
rect 19524 87610 19548 87612
rect 19604 87610 19628 87612
rect 19684 87610 19690 87612
rect 19444 87558 19446 87610
rect 19626 87558 19628 87610
rect 19382 87556 19388 87558
rect 19444 87556 19468 87558
rect 19524 87556 19548 87558
rect 19604 87556 19628 87558
rect 19684 87556 19690 87558
rect 19382 87547 19690 87556
rect 18722 87068 19030 87077
rect 18722 87066 18728 87068
rect 18784 87066 18808 87068
rect 18864 87066 18888 87068
rect 18944 87066 18968 87068
rect 19024 87066 19030 87068
rect 18784 87014 18786 87066
rect 18966 87014 18968 87066
rect 18722 87012 18728 87014
rect 18784 87012 18808 87014
rect 18864 87012 18888 87014
rect 18944 87012 18968 87014
rect 19024 87012 19030 87014
rect 18722 87003 19030 87012
rect 19382 86524 19690 86533
rect 19382 86522 19388 86524
rect 19444 86522 19468 86524
rect 19524 86522 19548 86524
rect 19604 86522 19628 86524
rect 19684 86522 19690 86524
rect 19444 86470 19446 86522
rect 19626 86470 19628 86522
rect 19382 86468 19388 86470
rect 19444 86468 19468 86470
rect 19524 86468 19548 86470
rect 19604 86468 19628 86470
rect 19684 86468 19690 86470
rect 19382 86459 19690 86468
rect 18652 84342 18850 84370
rect 19940 84356 19968 88778
rect 21044 84356 21072 88778
rect 22148 84356 22176 88778
rect 23252 84356 23280 88778
rect 24356 84356 24384 88846
rect 25448 88836 25500 88842
rect 25448 88778 25500 88784
rect 26552 88836 26604 88842
rect 26552 88778 26604 88784
rect 27656 88836 27708 88842
rect 27656 88778 27708 88784
rect 28760 88836 28812 88842
rect 28760 88778 28812 88784
rect 29864 88836 29916 88842
rect 29864 88778 29916 88784
rect 25460 84356 25488 88778
rect 26564 84356 26592 88778
rect 27668 84356 27696 88778
rect 28772 84356 28800 88778
rect 29876 84356 29904 88778
rect 30980 84356 31008 88846
rect 31704 86660 31756 86666
rect 31704 86602 31756 86608
rect 14406 84319 14462 84328
rect 7600 54768 7652 54774
rect 2538 54736 2594 54745
rect 7600 54710 7652 54716
rect 2538 54671 2594 54680
rect 7048 54564 7100 54570
rect 7048 54506 7100 54512
rect 5954 54428 6262 54437
rect 5954 54426 5960 54428
rect 6016 54426 6040 54428
rect 6096 54426 6120 54428
rect 6176 54426 6200 54428
rect 6256 54426 6262 54428
rect 6016 54374 6018 54426
rect 6198 54374 6200 54426
rect 5954 54372 5960 54374
rect 6016 54372 6040 54374
rect 6096 54372 6120 54374
rect 6176 54372 6200 54374
rect 6256 54372 6262 54374
rect 5954 54363 6262 54372
rect 5666 54192 5722 54201
rect 5666 54127 5722 54136
rect 5208 54088 5260 54094
rect 5206 54056 5208 54065
rect 5260 54056 5262 54065
rect 5206 53991 5262 54000
rect 5680 53754 5708 54127
rect 6690 53884 6998 53893
rect 6690 53882 6696 53884
rect 6752 53882 6776 53884
rect 6832 53882 6856 53884
rect 6912 53882 6936 53884
rect 6992 53882 6998 53884
rect 6752 53830 6754 53882
rect 6934 53830 6936 53882
rect 6690 53828 6696 53830
rect 6752 53828 6776 53830
rect 6832 53828 6856 53830
rect 6912 53828 6936 53830
rect 6992 53828 6998 53830
rect 6690 53819 6998 53828
rect 5668 53748 5720 53754
rect 5668 53690 5720 53696
rect 2908 53612 2960 53618
rect 2908 53554 2960 53560
rect 2920 53385 2948 53554
rect 2906 53376 2962 53385
rect 2906 53311 2962 53320
rect 5954 53340 6262 53349
rect 5954 53338 5960 53340
rect 6016 53338 6040 53340
rect 6096 53338 6120 53340
rect 6176 53338 6200 53340
rect 6256 53338 6262 53340
rect 6016 53286 6018 53338
rect 6198 53286 6200 53338
rect 5954 53284 5960 53286
rect 6016 53284 6040 53286
rect 6096 53284 6120 53286
rect 6176 53284 6200 53286
rect 6256 53284 6262 53286
rect 5954 53275 6262 53284
rect 2908 53000 2960 53006
rect 2908 52942 2960 52948
rect 2920 52705 2948 52942
rect 6690 52796 6998 52805
rect 6690 52794 6696 52796
rect 6752 52794 6776 52796
rect 6832 52794 6856 52796
rect 6912 52794 6936 52796
rect 6992 52794 6998 52796
rect 6752 52742 6754 52794
rect 6934 52742 6936 52794
rect 6690 52740 6696 52742
rect 6752 52740 6776 52742
rect 6832 52740 6856 52742
rect 6912 52740 6936 52742
rect 6992 52740 6998 52742
rect 6690 52731 6998 52740
rect 2906 52696 2962 52705
rect 2906 52631 2962 52640
rect 2908 52524 2960 52530
rect 2908 52466 2960 52472
rect 2920 52025 2948 52466
rect 5954 52252 6262 52261
rect 5954 52250 5960 52252
rect 6016 52250 6040 52252
rect 6096 52250 6120 52252
rect 6176 52250 6200 52252
rect 6256 52250 6262 52252
rect 6016 52198 6018 52250
rect 6198 52198 6200 52250
rect 5954 52196 5960 52198
rect 6016 52196 6040 52198
rect 6096 52196 6120 52198
rect 6176 52196 6200 52198
rect 6256 52196 6262 52198
rect 5954 52187 6262 52196
rect 2906 52016 2962 52025
rect 2906 51951 2962 51960
rect 6690 51708 6998 51717
rect 6690 51706 6696 51708
rect 6752 51706 6776 51708
rect 6832 51706 6856 51708
rect 6912 51706 6936 51708
rect 6992 51706 6998 51708
rect 6752 51654 6754 51706
rect 6934 51654 6936 51706
rect 6690 51652 6696 51654
rect 6752 51652 6776 51654
rect 6832 51652 6856 51654
rect 6912 51652 6936 51654
rect 6992 51652 6998 51654
rect 6690 51643 6998 51652
rect 2908 51436 2960 51442
rect 2908 51378 2960 51384
rect 2920 51345 2948 51378
rect 5668 51368 5720 51374
rect 2906 51336 2962 51345
rect 5668 51310 5720 51316
rect 2906 51271 2962 51280
rect 5680 50937 5708 51310
rect 5954 51164 6262 51173
rect 5954 51162 5960 51164
rect 6016 51162 6040 51164
rect 6096 51162 6120 51164
rect 6176 51162 6200 51164
rect 6256 51162 6262 51164
rect 6016 51110 6018 51162
rect 6198 51110 6200 51162
rect 5954 51108 5960 51110
rect 6016 51108 6040 51110
rect 6096 51108 6120 51110
rect 6176 51108 6200 51110
rect 6256 51108 6262 51110
rect 5954 51099 6262 51108
rect 5666 50928 5722 50937
rect 5666 50863 5722 50872
rect 6690 50620 6998 50629
rect 6690 50618 6696 50620
rect 6752 50618 6776 50620
rect 6832 50618 6856 50620
rect 6912 50618 6936 50620
rect 6992 50618 6998 50620
rect 6752 50566 6754 50618
rect 6934 50566 6936 50618
rect 6690 50564 6696 50566
rect 6752 50564 6776 50566
rect 6832 50564 6856 50566
rect 6912 50564 6936 50566
rect 6992 50564 6998 50566
rect 6690 50555 6998 50564
rect 5954 50076 6262 50085
rect 5954 50074 5960 50076
rect 6016 50074 6040 50076
rect 6096 50074 6120 50076
rect 6176 50074 6200 50076
rect 6256 50074 6262 50076
rect 6016 50022 6018 50074
rect 6198 50022 6200 50074
rect 5954 50020 5960 50022
rect 6016 50020 6040 50022
rect 6096 50020 6120 50022
rect 6176 50020 6200 50022
rect 6256 50020 6262 50022
rect 5954 50011 6262 50020
rect 2908 49736 2960 49742
rect 2908 49678 2960 49684
rect 2920 49305 2948 49678
rect 6690 49532 6998 49541
rect 6690 49530 6696 49532
rect 6752 49530 6776 49532
rect 6832 49530 6856 49532
rect 6912 49530 6936 49532
rect 6992 49530 6998 49532
rect 6752 49478 6754 49530
rect 6934 49478 6936 49530
rect 6690 49476 6696 49478
rect 6752 49476 6776 49478
rect 6832 49476 6856 49478
rect 6912 49476 6936 49478
rect 6992 49476 6998 49478
rect 6690 49467 6998 49476
rect 2906 49296 2962 49305
rect 2906 49231 2962 49240
rect 5954 48988 6262 48997
rect 5954 48986 5960 48988
rect 6016 48986 6040 48988
rect 6096 48986 6120 48988
rect 6176 48986 6200 48988
rect 6256 48986 6262 48988
rect 6016 48934 6018 48986
rect 6198 48934 6200 48986
rect 5954 48932 5960 48934
rect 6016 48932 6040 48934
rect 6096 48932 6120 48934
rect 6176 48932 6200 48934
rect 6256 48932 6262 48934
rect 5954 48923 6262 48932
rect 6690 48444 6998 48453
rect 6690 48442 6696 48444
rect 6752 48442 6776 48444
rect 6832 48442 6856 48444
rect 6912 48442 6936 48444
rect 6992 48442 6998 48444
rect 6752 48390 6754 48442
rect 6934 48390 6936 48442
rect 6690 48388 6696 48390
rect 6752 48388 6776 48390
rect 6832 48388 6856 48390
rect 6912 48388 6936 48390
rect 6992 48388 6998 48390
rect 6690 48379 6998 48388
rect 5954 47900 6262 47909
rect 5954 47898 5960 47900
rect 6016 47898 6040 47900
rect 6096 47898 6120 47900
rect 6176 47898 6200 47900
rect 6256 47898 6262 47900
rect 6016 47846 6018 47898
rect 6198 47846 6200 47898
rect 5954 47844 5960 47846
rect 6016 47844 6040 47846
rect 6096 47844 6120 47846
rect 6176 47844 6200 47846
rect 6256 47844 6262 47846
rect 5954 47835 6262 47844
rect 6690 47356 6998 47365
rect 6690 47354 6696 47356
rect 6752 47354 6776 47356
rect 6832 47354 6856 47356
rect 6912 47354 6936 47356
rect 6992 47354 6998 47356
rect 6752 47302 6754 47354
rect 6934 47302 6936 47354
rect 6690 47300 6696 47302
rect 6752 47300 6776 47302
rect 6832 47300 6856 47302
rect 6912 47300 6936 47302
rect 6992 47300 6998 47302
rect 6690 47291 6998 47300
rect 7060 47158 7088 54506
rect 7138 53240 7194 53249
rect 7138 53175 7140 53184
rect 7192 53175 7194 53184
rect 7140 53146 7192 53152
rect 7140 52388 7192 52394
rect 7140 52330 7192 52336
rect 7152 52161 7180 52330
rect 7138 52152 7194 52161
rect 7138 52087 7194 52096
rect 8152 47288 8204 47294
rect 8152 47230 8204 47236
rect 8334 47256 8390 47265
rect 7876 47220 7928 47226
rect 7876 47162 7928 47168
rect 2908 47152 2960 47158
rect 2908 47094 2960 47100
rect 7048 47152 7100 47158
rect 7048 47094 7100 47100
rect 2920 46585 2948 47094
rect 5954 46812 6262 46821
rect 5954 46810 5960 46812
rect 6016 46810 6040 46812
rect 6096 46810 6120 46812
rect 6176 46810 6200 46812
rect 6256 46810 6262 46812
rect 6016 46758 6018 46810
rect 6198 46758 6200 46810
rect 5954 46756 5960 46758
rect 6016 46756 6040 46758
rect 6096 46756 6120 46758
rect 6176 46756 6200 46758
rect 6256 46756 6262 46758
rect 5954 46747 6262 46756
rect 2906 46576 2962 46585
rect 2906 46511 2962 46520
rect 6690 46268 6998 46277
rect 6690 46266 6696 46268
rect 6752 46266 6776 46268
rect 6832 46266 6856 46268
rect 6912 46266 6936 46268
rect 6992 46266 6998 46268
rect 6752 46214 6754 46266
rect 6934 46214 6936 46266
rect 6690 46212 6696 46214
rect 6752 46212 6776 46214
rect 6832 46212 6856 46214
rect 6912 46212 6936 46214
rect 6992 46212 6998 46214
rect 6690 46203 6998 46212
rect 2906 45896 2962 45905
rect 2906 45831 2908 45840
rect 2960 45831 2962 45840
rect 2908 45802 2960 45808
rect 5954 45724 6262 45733
rect 5954 45722 5960 45724
rect 6016 45722 6040 45724
rect 6096 45722 6120 45724
rect 6176 45722 6200 45724
rect 6256 45722 6262 45724
rect 6016 45670 6018 45722
rect 6198 45670 6200 45722
rect 5954 45668 5960 45670
rect 6016 45668 6040 45670
rect 6096 45668 6120 45670
rect 6176 45668 6200 45670
rect 6256 45668 6262 45670
rect 5954 45659 6262 45668
rect 6690 45180 6998 45189
rect 6690 45178 6696 45180
rect 6752 45178 6776 45180
rect 6832 45178 6856 45180
rect 6912 45178 6936 45180
rect 6992 45178 6998 45180
rect 6752 45126 6754 45178
rect 6934 45126 6936 45178
rect 6690 45124 6696 45126
rect 6752 45124 6776 45126
rect 6832 45124 6856 45126
rect 6912 45124 6936 45126
rect 6992 45124 6998 45126
rect 6690 45115 6998 45124
rect 2540 44772 2592 44778
rect 2540 44714 2592 44720
rect 2552 44545 2580 44714
rect 5954 44636 6262 44645
rect 5954 44634 5960 44636
rect 6016 44634 6040 44636
rect 6096 44634 6120 44636
rect 6176 44634 6200 44636
rect 6256 44634 6262 44636
rect 6016 44582 6018 44634
rect 6198 44582 6200 44634
rect 5954 44580 5960 44582
rect 6016 44580 6040 44582
rect 6096 44580 6120 44582
rect 6176 44580 6200 44582
rect 6256 44580 6262 44582
rect 5954 44571 6262 44580
rect 2538 44536 2594 44545
rect 2538 44471 2594 44480
rect 5208 44432 5260 44438
rect 5208 44374 5260 44380
rect 5220 43865 5248 44374
rect 6690 44092 6998 44101
rect 6690 44090 6696 44092
rect 6752 44090 6776 44092
rect 6832 44090 6856 44092
rect 6912 44090 6936 44092
rect 6992 44090 6998 44092
rect 6752 44038 6754 44090
rect 6934 44038 6936 44090
rect 6690 44036 6696 44038
rect 6752 44036 6776 44038
rect 6832 44036 6856 44038
rect 6912 44036 6936 44038
rect 6992 44036 6998 44038
rect 6690 44027 6998 44036
rect 5206 43856 5262 43865
rect 5206 43791 5262 43800
rect 5954 43548 6262 43557
rect 5954 43546 5960 43548
rect 6016 43546 6040 43548
rect 6096 43546 6120 43548
rect 6176 43546 6200 43548
rect 6256 43546 6262 43548
rect 6016 43494 6018 43546
rect 6198 43494 6200 43546
rect 5954 43492 5960 43494
rect 6016 43492 6040 43494
rect 6096 43492 6120 43494
rect 6176 43492 6200 43494
rect 6256 43492 6262 43494
rect 5954 43483 6262 43492
rect 7140 43208 7192 43214
rect 2906 43176 2962 43185
rect 7140 43150 7192 43156
rect 2906 43111 2908 43120
rect 2960 43111 2962 43120
rect 2908 43082 2960 43088
rect 7152 43049 7180 43150
rect 7138 43040 7194 43049
rect 6690 43004 6998 43013
rect 6690 43002 6696 43004
rect 6752 43002 6776 43004
rect 6832 43002 6856 43004
rect 6912 43002 6936 43004
rect 6992 43002 6998 43004
rect 6752 42950 6754 43002
rect 6934 42950 6936 43002
rect 7138 42975 7194 42984
rect 6690 42948 6696 42950
rect 6752 42948 6776 42950
rect 6832 42948 6856 42950
rect 6912 42948 6936 42950
rect 6992 42948 6998 42950
rect 6690 42939 6998 42948
rect 2908 42596 2960 42602
rect 2908 42538 2960 42544
rect 2920 42505 2948 42538
rect 2906 42496 2962 42505
rect 2906 42431 2962 42440
rect 5954 42460 6262 42469
rect 5954 42458 5960 42460
rect 6016 42458 6040 42460
rect 6096 42458 6120 42460
rect 6176 42458 6200 42460
rect 6256 42458 6262 42460
rect 6016 42406 6018 42458
rect 6198 42406 6200 42458
rect 5954 42404 5960 42406
rect 6016 42404 6040 42406
rect 6096 42404 6120 42406
rect 6176 42404 6200 42406
rect 6256 42404 6262 42406
rect 5954 42395 6262 42404
rect 7140 42120 7192 42126
rect 7140 42062 7192 42068
rect 2908 42052 2960 42058
rect 2908 41994 2960 42000
rect 2920 41825 2948 41994
rect 7152 41961 7180 42062
rect 7138 41952 7194 41961
rect 6690 41916 6998 41925
rect 6690 41914 6696 41916
rect 6752 41914 6776 41916
rect 6832 41914 6856 41916
rect 6912 41914 6936 41916
rect 6992 41914 6998 41916
rect 6752 41862 6754 41914
rect 6934 41862 6936 41914
rect 7138 41887 7194 41896
rect 6690 41860 6696 41862
rect 6752 41860 6776 41862
rect 6832 41860 6856 41862
rect 6912 41860 6936 41862
rect 6992 41860 6998 41862
rect 6690 41851 6998 41860
rect 2906 41816 2962 41825
rect 2906 41751 2962 41760
rect 4380 41780 4432 41786
rect 4380 41722 4432 41728
rect 4392 41145 4420 41722
rect 5668 41678 5720 41684
rect 5668 41620 5720 41626
rect 4378 41136 4434 41145
rect 4378 41071 4434 41080
rect 5680 41009 5708 41620
rect 5954 41372 6262 41381
rect 5954 41370 5960 41372
rect 6016 41370 6040 41372
rect 6096 41370 6120 41372
rect 6176 41370 6200 41372
rect 6256 41370 6262 41372
rect 6016 41318 6018 41370
rect 6198 41318 6200 41370
rect 5954 41316 5960 41318
rect 6016 41316 6040 41318
rect 6096 41316 6120 41318
rect 6176 41316 6200 41318
rect 6256 41316 6262 41318
rect 5954 41307 6262 41316
rect 5666 41000 5722 41009
rect 5666 40935 5722 40944
rect 6690 40828 6998 40837
rect 6690 40826 6696 40828
rect 6752 40826 6776 40828
rect 6832 40826 6856 40828
rect 6912 40826 6936 40828
rect 6992 40826 6998 40828
rect 6752 40774 6754 40826
rect 6934 40774 6936 40826
rect 6690 40772 6696 40774
rect 6752 40772 6776 40774
rect 6832 40772 6856 40774
rect 6912 40772 6936 40774
rect 6992 40772 6998 40774
rect 6690 40763 6998 40772
rect 5954 40284 6262 40293
rect 5954 40282 5960 40284
rect 6016 40282 6040 40284
rect 6096 40282 6120 40284
rect 6176 40282 6200 40284
rect 6256 40282 6262 40284
rect 6016 40230 6018 40282
rect 6198 40230 6200 40282
rect 5954 40228 5960 40230
rect 6016 40228 6040 40230
rect 6096 40228 6120 40230
rect 6176 40228 6200 40230
rect 6256 40228 6262 40230
rect 5954 40219 6262 40228
rect 7140 39944 7192 39950
rect 7140 39886 7192 39892
rect 2908 39876 2960 39882
rect 2908 39818 2960 39824
rect 2920 39785 2948 39818
rect 7152 39785 7180 39886
rect 2906 39776 2962 39785
rect 7138 39776 7194 39785
rect 2906 39711 2962 39720
rect 6690 39740 6998 39749
rect 6690 39738 6696 39740
rect 6752 39738 6776 39740
rect 6832 39738 6856 39740
rect 6912 39738 6936 39740
rect 6992 39738 6998 39740
rect 6752 39686 6754 39738
rect 6934 39686 6936 39738
rect 7138 39711 7194 39720
rect 6690 39684 6696 39686
rect 6752 39684 6776 39686
rect 6832 39684 6856 39686
rect 6912 39684 6936 39686
rect 6992 39684 6998 39686
rect 6690 39675 6998 39684
rect 5954 39196 6262 39205
rect 5954 39194 5960 39196
rect 6016 39194 6040 39196
rect 6096 39194 6120 39196
rect 6176 39194 6200 39196
rect 6256 39194 6262 39196
rect 6016 39142 6018 39194
rect 6198 39142 6200 39194
rect 5954 39140 5960 39142
rect 6016 39140 6040 39142
rect 6096 39140 6120 39142
rect 6176 39140 6200 39142
rect 6256 39140 6262 39142
rect 5954 39131 6262 39140
rect 4380 38992 4432 38998
rect 4380 38934 4432 38940
rect 4392 38425 4420 38934
rect 7416 38856 7468 38862
rect 7416 38798 7468 38804
rect 7428 38697 7456 38798
rect 7414 38688 7470 38697
rect 6690 38652 6998 38661
rect 6690 38650 6696 38652
rect 6752 38650 6776 38652
rect 6832 38650 6856 38652
rect 6912 38650 6936 38652
rect 6992 38650 6998 38652
rect 6752 38598 6754 38650
rect 6934 38598 6936 38650
rect 7414 38623 7470 38632
rect 6690 38596 6696 38598
rect 6752 38596 6776 38598
rect 6832 38596 6856 38598
rect 6912 38596 6936 38598
rect 6992 38596 6998 38598
rect 6690 38587 6998 38596
rect 4378 38416 4434 38425
rect 4378 38351 4434 38360
rect 5954 38108 6262 38117
rect 5954 38106 5960 38108
rect 6016 38106 6040 38108
rect 6096 38106 6120 38108
rect 6176 38106 6200 38108
rect 6256 38106 6262 38108
rect 6016 38054 6018 38106
rect 6198 38054 6200 38106
rect 5954 38052 5960 38054
rect 6016 38052 6040 38054
rect 6096 38052 6120 38054
rect 6176 38052 6200 38054
rect 6256 38052 6262 38054
rect 5954 38043 6262 38052
rect 7140 37768 7192 37774
rect 2906 37736 2962 37745
rect 7140 37710 7192 37716
rect 2906 37671 2908 37680
rect 2960 37671 2962 37680
rect 2908 37642 2960 37648
rect 7152 37609 7180 37710
rect 7138 37600 7194 37609
rect 6690 37564 6998 37573
rect 6690 37562 6696 37564
rect 6752 37562 6776 37564
rect 6832 37562 6856 37564
rect 6912 37562 6936 37564
rect 6992 37562 6998 37564
rect 6752 37510 6754 37562
rect 6934 37510 6936 37562
rect 7138 37535 7194 37544
rect 6690 37508 6696 37510
rect 6752 37508 6776 37510
rect 6832 37508 6856 37510
rect 6912 37508 6936 37510
rect 6992 37508 6998 37510
rect 6690 37499 6998 37508
rect 5954 37020 6262 37029
rect 5954 37018 5960 37020
rect 6016 37018 6040 37020
rect 6096 37018 6120 37020
rect 6176 37018 6200 37020
rect 6256 37018 6262 37020
rect 6016 36966 6018 37018
rect 6198 36966 6200 37018
rect 5954 36964 5960 36966
rect 6016 36964 6040 36966
rect 6096 36964 6120 36966
rect 6176 36964 6200 36966
rect 6256 36964 6262 36966
rect 5954 36955 6262 36964
rect 7140 36680 7192 36686
rect 7140 36622 7192 36628
rect 2908 36612 2960 36618
rect 2908 36554 2960 36560
rect 2920 36385 2948 36554
rect 7152 36521 7180 36622
rect 7138 36512 7194 36521
rect 6690 36476 6998 36485
rect 6690 36474 6696 36476
rect 6752 36474 6776 36476
rect 6832 36474 6856 36476
rect 6912 36474 6936 36476
rect 6992 36474 6998 36476
rect 6752 36422 6754 36474
rect 6934 36422 6936 36474
rect 7138 36447 7194 36456
rect 6690 36420 6696 36422
rect 6752 36420 6776 36422
rect 6832 36420 6856 36422
rect 6912 36420 6936 36422
rect 6992 36420 6998 36422
rect 6690 36411 6998 36420
rect 2906 36376 2962 36385
rect 2906 36311 2962 36320
rect 5668 36238 5720 36244
rect 5668 36180 5720 36186
rect 4380 36136 4432 36142
rect 4380 36078 4432 36084
rect 4392 35705 4420 36078
rect 4378 35696 4434 35705
rect 4378 35631 4434 35640
rect 5680 35569 5708 36180
rect 5954 35932 6262 35941
rect 5954 35930 5960 35932
rect 6016 35930 6040 35932
rect 6096 35930 6120 35932
rect 6176 35930 6200 35932
rect 6256 35930 6262 35932
rect 6016 35878 6018 35930
rect 6198 35878 6200 35930
rect 5954 35876 5960 35878
rect 6016 35876 6040 35878
rect 6096 35876 6120 35878
rect 6176 35876 6200 35878
rect 6256 35876 6262 35878
rect 5954 35867 6262 35876
rect 5666 35560 5722 35569
rect 5666 35495 5722 35504
rect 6690 35388 6998 35397
rect 6690 35386 6696 35388
rect 6752 35386 6776 35388
rect 6832 35386 6856 35388
rect 6912 35386 6936 35388
rect 6992 35386 6998 35388
rect 6752 35334 6754 35386
rect 6934 35334 6936 35386
rect 6690 35332 6696 35334
rect 6752 35332 6776 35334
rect 6832 35332 6856 35334
rect 6912 35332 6936 35334
rect 6992 35332 6998 35334
rect 6690 35323 6998 35332
rect 5954 34844 6262 34853
rect 5954 34842 5960 34844
rect 6016 34842 6040 34844
rect 6096 34842 6120 34844
rect 6176 34842 6200 34844
rect 6256 34842 6262 34844
rect 6016 34790 6018 34842
rect 6198 34790 6200 34842
rect 5954 34788 5960 34790
rect 6016 34788 6040 34790
rect 6096 34788 6120 34790
rect 6176 34788 6200 34790
rect 6256 34788 6262 34790
rect 5954 34779 6262 34788
rect 7140 34504 7192 34510
rect 7140 34446 7192 34452
rect 2908 34436 2960 34442
rect 2908 34378 2960 34384
rect 2920 34345 2948 34378
rect 7152 34345 7180 34446
rect 2906 34336 2962 34345
rect 7138 34336 7194 34345
rect 2906 34271 2962 34280
rect 6690 34300 6998 34309
rect 6690 34298 6696 34300
rect 6752 34298 6776 34300
rect 6832 34298 6856 34300
rect 6912 34298 6936 34300
rect 6992 34298 6998 34300
rect 6752 34246 6754 34298
rect 6934 34246 6936 34298
rect 7138 34271 7194 34280
rect 6690 34244 6696 34246
rect 6752 34244 6776 34246
rect 6832 34244 6856 34246
rect 6912 34244 6936 34246
rect 6992 34244 6998 34246
rect 6690 34235 6998 34244
rect 2908 33892 2960 33898
rect 2908 33834 2960 33840
rect 2920 33665 2948 33834
rect 5954 33756 6262 33765
rect 5954 33754 5960 33756
rect 6016 33754 6040 33756
rect 6096 33754 6120 33756
rect 6176 33754 6200 33756
rect 6256 33754 6262 33756
rect 6016 33702 6018 33754
rect 6198 33702 6200 33754
rect 5954 33700 5960 33702
rect 6016 33700 6040 33702
rect 6096 33700 6120 33702
rect 6176 33700 6200 33702
rect 6256 33700 6262 33702
rect 5954 33691 6262 33700
rect 2906 33656 2962 33665
rect 2906 33591 2962 33600
rect 4380 33552 4432 33558
rect 4380 33494 4432 33500
rect 4392 32985 4420 33494
rect 5668 33450 5720 33456
rect 5668 33392 5720 33398
rect 5680 32985 5708 33392
rect 6690 33212 6998 33221
rect 6690 33210 6696 33212
rect 6752 33210 6776 33212
rect 6832 33210 6856 33212
rect 6912 33210 6936 33212
rect 6992 33210 6998 33212
rect 6752 33158 6754 33210
rect 6934 33158 6936 33210
rect 6690 33156 6696 33158
rect 6752 33156 6776 33158
rect 6832 33156 6856 33158
rect 6912 33156 6936 33158
rect 6992 33156 6998 33158
rect 6690 33147 6998 33156
rect 4378 32976 4434 32985
rect 4378 32911 4434 32920
rect 5666 32976 5722 32985
rect 5666 32911 5722 32920
rect 5954 32668 6262 32677
rect 5954 32666 5960 32668
rect 6016 32666 6040 32668
rect 6096 32666 6120 32668
rect 6176 32666 6200 32668
rect 6256 32666 6262 32668
rect 6016 32614 6018 32666
rect 6198 32614 6200 32666
rect 5954 32612 5960 32614
rect 6016 32612 6040 32614
rect 6096 32612 6120 32614
rect 6176 32612 6200 32614
rect 6256 32612 6262 32614
rect 5954 32603 6262 32612
rect 7140 32328 7192 32334
rect 2906 32296 2962 32305
rect 7140 32270 7192 32276
rect 2906 32231 2908 32240
rect 2960 32231 2962 32240
rect 2908 32202 2960 32208
rect 7152 32169 7180 32270
rect 7138 32160 7194 32169
rect 6690 32124 6998 32133
rect 6690 32122 6696 32124
rect 6752 32122 6776 32124
rect 6832 32122 6856 32124
rect 6912 32122 6936 32124
rect 6992 32122 6998 32124
rect 6752 32070 6754 32122
rect 6934 32070 6936 32122
rect 7138 32095 7194 32104
rect 6690 32068 6696 32070
rect 6752 32068 6776 32070
rect 6832 32068 6856 32070
rect 6912 32068 6936 32070
rect 6992 32068 6998 32070
rect 6690 32059 6998 32068
rect 5954 31580 6262 31589
rect 5954 31578 5960 31580
rect 6016 31578 6040 31580
rect 6096 31578 6120 31580
rect 6176 31578 6200 31580
rect 6256 31578 6262 31580
rect 6016 31526 6018 31578
rect 6198 31526 6200 31578
rect 5954 31524 5960 31526
rect 6016 31524 6040 31526
rect 6096 31524 6120 31526
rect 6176 31524 6200 31526
rect 6256 31524 6262 31526
rect 5954 31515 6262 31524
rect 7140 31240 7192 31246
rect 7140 31182 7192 31188
rect 2908 31172 2960 31178
rect 2908 31114 2960 31120
rect 2920 30945 2948 31114
rect 7152 31081 7180 31182
rect 7138 31072 7194 31081
rect 6690 31036 6998 31045
rect 6690 31034 6696 31036
rect 6752 31034 6776 31036
rect 6832 31034 6856 31036
rect 6912 31034 6936 31036
rect 6992 31034 6998 31036
rect 6752 30982 6754 31034
rect 6934 30982 6936 31034
rect 7138 31007 7194 31016
rect 6690 30980 6696 30982
rect 6752 30980 6776 30982
rect 6832 30980 6856 30982
rect 6912 30980 6936 30982
rect 6992 30980 6998 30982
rect 6690 30971 6998 30980
rect 2906 30936 2962 30945
rect 2906 30871 2962 30880
rect 5668 30798 5720 30804
rect 5668 30740 5720 30746
rect 4380 30628 4432 30634
rect 4380 30570 4432 30576
rect 4392 30265 4420 30570
rect 4378 30256 4434 30265
rect 4378 30191 4434 30200
rect 5680 30129 5708 30740
rect 5954 30492 6262 30501
rect 5954 30490 5960 30492
rect 6016 30490 6040 30492
rect 6096 30490 6120 30492
rect 6176 30490 6200 30492
rect 6256 30490 6262 30492
rect 6016 30438 6018 30490
rect 6198 30438 6200 30490
rect 5954 30436 5960 30438
rect 6016 30436 6040 30438
rect 6096 30436 6120 30438
rect 6176 30436 6200 30438
rect 6256 30436 6262 30438
rect 5954 30427 6262 30436
rect 5666 30120 5722 30129
rect 5666 30055 5722 30064
rect 6690 29948 6998 29957
rect 6690 29946 6696 29948
rect 6752 29946 6776 29948
rect 6832 29946 6856 29948
rect 6912 29946 6936 29948
rect 6992 29946 6998 29948
rect 6752 29894 6754 29946
rect 6934 29894 6936 29946
rect 6690 29892 6696 29894
rect 6752 29892 6776 29894
rect 6832 29892 6856 29894
rect 6912 29892 6936 29894
rect 6992 29892 6998 29894
rect 6690 29883 6998 29892
rect 5954 29404 6262 29413
rect 5954 29402 5960 29404
rect 6016 29402 6040 29404
rect 6096 29402 6120 29404
rect 6176 29402 6200 29404
rect 6256 29402 6262 29404
rect 6016 29350 6018 29402
rect 6198 29350 6200 29402
rect 5954 29348 5960 29350
rect 6016 29348 6040 29350
rect 6096 29348 6120 29350
rect 6176 29348 6200 29350
rect 6256 29348 6262 29350
rect 5954 29339 6262 29348
rect 7140 29064 7192 29070
rect 7140 29006 7192 29012
rect 2908 28996 2960 29002
rect 2908 28938 2960 28944
rect 2920 28905 2948 28938
rect 7152 28905 7180 29006
rect 2906 28896 2962 28905
rect 7138 28896 7194 28905
rect 2906 28831 2962 28840
rect 6690 28860 6998 28869
rect 6690 28858 6696 28860
rect 6752 28858 6776 28860
rect 6832 28858 6856 28860
rect 6912 28858 6936 28860
rect 6992 28858 6998 28860
rect 6752 28806 6754 28858
rect 6934 28806 6936 28858
rect 7138 28831 7194 28840
rect 6690 28804 6696 28806
rect 6752 28804 6776 28806
rect 6832 28804 6856 28806
rect 6912 28804 6936 28806
rect 6992 28804 6998 28806
rect 6690 28795 6998 28804
rect 5954 28316 6262 28325
rect 5954 28314 5960 28316
rect 6016 28314 6040 28316
rect 6096 28314 6120 28316
rect 6176 28314 6200 28316
rect 6256 28314 6262 28316
rect 6016 28262 6018 28314
rect 6198 28262 6200 28314
rect 5954 28260 5960 28262
rect 6016 28260 6040 28262
rect 6096 28260 6120 28262
rect 6176 28260 6200 28262
rect 6256 28260 6262 28262
rect 5954 28251 6262 28260
rect 5116 28010 5168 28016
rect 5116 27952 5168 27958
rect 5128 27545 5156 27952
rect 5392 27908 5444 27914
rect 5392 27850 5444 27856
rect 5404 27545 5432 27850
rect 6690 27772 6998 27781
rect 6690 27770 6696 27772
rect 6752 27770 6776 27772
rect 6832 27770 6856 27772
rect 6912 27770 6936 27772
rect 6992 27770 6998 27772
rect 6752 27718 6754 27770
rect 6934 27718 6936 27770
rect 6690 27716 6696 27718
rect 6752 27716 6776 27718
rect 6832 27716 6856 27718
rect 6912 27716 6936 27718
rect 6992 27716 6998 27718
rect 6690 27707 6998 27716
rect 5114 27536 5170 27545
rect 5114 27471 5170 27480
rect 5390 27536 5446 27545
rect 5390 27471 5446 27480
rect 5954 27228 6262 27237
rect 5954 27226 5960 27228
rect 6016 27226 6040 27228
rect 6096 27226 6120 27228
rect 6176 27226 6200 27228
rect 6256 27226 6262 27228
rect 6016 27174 6018 27226
rect 6198 27174 6200 27226
rect 5954 27172 5960 27174
rect 6016 27172 6040 27174
rect 6096 27172 6120 27174
rect 6176 27172 6200 27174
rect 6256 27172 6262 27174
rect 5954 27163 6262 27172
rect 2908 26888 2960 26894
rect 2906 26856 2908 26865
rect 2960 26856 2962 26865
rect 2906 26791 2962 26800
rect 7140 26820 7192 26826
rect 7140 26762 7192 26768
rect 7152 26729 7180 26762
rect 7138 26720 7194 26729
rect 6690 26684 6998 26693
rect 6690 26682 6696 26684
rect 6752 26682 6776 26684
rect 6832 26682 6856 26684
rect 6912 26682 6936 26684
rect 6992 26682 6998 26684
rect 6752 26630 6754 26682
rect 6934 26630 6936 26682
rect 7138 26655 7194 26664
rect 6690 26628 6696 26630
rect 6752 26628 6776 26630
rect 6832 26628 6856 26630
rect 6912 26628 6936 26630
rect 6992 26628 6998 26630
rect 6690 26619 6998 26628
rect 5954 26140 6262 26149
rect 5954 26138 5960 26140
rect 6016 26138 6040 26140
rect 6096 26138 6120 26140
rect 6176 26138 6200 26140
rect 6256 26138 6262 26140
rect 6016 26086 6018 26138
rect 6198 26086 6200 26138
rect 5954 26084 5960 26086
rect 6016 26084 6040 26086
rect 6096 26084 6120 26086
rect 6176 26084 6200 26086
rect 6256 26084 6262 26086
rect 5954 26075 6262 26084
rect 2908 25800 2960 25806
rect 2908 25742 2960 25748
rect 2920 25505 2948 25742
rect 7140 25732 7192 25738
rect 7140 25674 7192 25680
rect 7152 25641 7180 25674
rect 7138 25632 7194 25641
rect 6690 25596 6998 25605
rect 6690 25594 6696 25596
rect 6752 25594 6776 25596
rect 6832 25594 6856 25596
rect 6912 25594 6936 25596
rect 6992 25594 6998 25596
rect 6752 25542 6754 25594
rect 6934 25542 6936 25594
rect 7138 25567 7194 25576
rect 6690 25540 6696 25542
rect 6752 25540 6776 25542
rect 6832 25540 6856 25542
rect 6912 25540 6936 25542
rect 6992 25540 6998 25542
rect 6690 25531 6998 25540
rect 2906 25496 2962 25505
rect 2906 25431 2962 25440
rect 4932 25358 4984 25364
rect 4932 25300 4984 25306
rect 4944 24825 4972 25300
rect 5668 25188 5720 25194
rect 5668 25130 5720 25136
rect 4930 24816 4986 24825
rect 4930 24751 4986 24760
rect 5680 24689 5708 25130
rect 5954 25052 6262 25061
rect 5954 25050 5960 25052
rect 6016 25050 6040 25052
rect 6096 25050 6120 25052
rect 6176 25050 6200 25052
rect 6256 25050 6262 25052
rect 6016 24998 6018 25050
rect 6198 24998 6200 25050
rect 5954 24996 5960 24998
rect 6016 24996 6040 24998
rect 6096 24996 6120 24998
rect 6176 24996 6200 24998
rect 6256 24996 6262 24998
rect 5954 24987 6262 24996
rect 5666 24680 5722 24689
rect 5666 24615 5722 24624
rect 6690 24508 6998 24517
rect 6690 24506 6696 24508
rect 6752 24506 6776 24508
rect 6832 24506 6856 24508
rect 6912 24506 6936 24508
rect 6992 24506 6998 24508
rect 6752 24454 6754 24506
rect 6934 24454 6936 24506
rect 6690 24452 6696 24454
rect 6752 24452 6776 24454
rect 6832 24452 6856 24454
rect 6912 24452 6936 24454
rect 6992 24452 6998 24454
rect 6690 24443 6998 24452
rect 5954 23964 6262 23973
rect 5954 23962 5960 23964
rect 6016 23962 6040 23964
rect 6096 23962 6120 23964
rect 6176 23962 6200 23964
rect 6256 23962 6262 23964
rect 6016 23910 6018 23962
rect 6198 23910 6200 23962
rect 5954 23908 5960 23910
rect 6016 23908 6040 23910
rect 6096 23908 6120 23910
rect 6176 23908 6200 23910
rect 6256 23908 6262 23910
rect 5954 23899 6262 23908
rect 2908 23624 2960 23630
rect 2908 23566 2960 23572
rect 2920 23465 2948 23566
rect 7140 23556 7192 23562
rect 7140 23498 7192 23504
rect 7152 23465 7180 23498
rect 2906 23456 2962 23465
rect 7138 23456 7194 23465
rect 2906 23391 2962 23400
rect 6690 23420 6998 23429
rect 6690 23418 6696 23420
rect 6752 23418 6776 23420
rect 6832 23418 6856 23420
rect 6912 23418 6936 23420
rect 6992 23418 6998 23420
rect 6752 23366 6754 23418
rect 6934 23366 6936 23418
rect 7138 23391 7194 23400
rect 6690 23364 6696 23366
rect 6752 23364 6776 23366
rect 6832 23364 6856 23366
rect 6912 23364 6936 23366
rect 6992 23364 6998 23366
rect 6690 23355 6998 23364
rect 5954 22876 6262 22885
rect 5954 22874 5960 22876
rect 6016 22874 6040 22876
rect 6096 22874 6120 22876
rect 6176 22874 6200 22876
rect 6256 22874 6262 22876
rect 6016 22822 6018 22874
rect 6198 22822 6200 22874
rect 5954 22820 5960 22822
rect 6016 22820 6040 22822
rect 6096 22820 6120 22822
rect 6176 22820 6200 22822
rect 6256 22820 6262 22822
rect 5954 22811 6262 22820
rect 5208 22570 5260 22576
rect 5208 22512 5260 22518
rect 5220 22105 5248 22512
rect 7140 22468 7192 22474
rect 7140 22410 7192 22416
rect 7152 22377 7180 22410
rect 7138 22368 7194 22377
rect 6690 22332 6998 22341
rect 6690 22330 6696 22332
rect 6752 22330 6776 22332
rect 6832 22330 6856 22332
rect 6912 22330 6936 22332
rect 6992 22330 6998 22332
rect 6752 22278 6754 22330
rect 6934 22278 6936 22330
rect 7138 22303 7194 22312
rect 6690 22276 6696 22278
rect 6752 22276 6776 22278
rect 6832 22276 6856 22278
rect 6912 22276 6936 22278
rect 6992 22276 6998 22278
rect 6690 22267 6998 22276
rect 5206 22096 5262 22105
rect 5206 22031 5262 22040
rect 5954 21788 6262 21797
rect 5954 21786 5960 21788
rect 6016 21786 6040 21788
rect 6096 21786 6120 21788
rect 6176 21786 6200 21788
rect 6256 21786 6262 21788
rect 6016 21734 6018 21786
rect 6198 21734 6200 21786
rect 5954 21732 5960 21734
rect 6016 21732 6040 21734
rect 6096 21732 6120 21734
rect 6176 21732 6200 21734
rect 6256 21732 6262 21734
rect 5954 21723 6262 21732
rect 2908 21448 2960 21454
rect 2906 21416 2908 21425
rect 2960 21416 2962 21425
rect 2906 21351 2962 21360
rect 7140 21380 7192 21386
rect 7140 21322 7192 21328
rect 7152 21289 7180 21322
rect 7138 21280 7194 21289
rect 6690 21244 6998 21253
rect 6690 21242 6696 21244
rect 6752 21242 6776 21244
rect 6832 21242 6856 21244
rect 6912 21242 6936 21244
rect 6992 21242 6998 21244
rect 6752 21190 6754 21242
rect 6934 21190 6936 21242
rect 7138 21215 7194 21224
rect 6690 21188 6696 21190
rect 6752 21188 6776 21190
rect 6832 21188 6856 21190
rect 6912 21188 6936 21190
rect 6992 21188 6998 21190
rect 6690 21179 6998 21188
rect 5954 20700 6262 20709
rect 5954 20698 5960 20700
rect 6016 20698 6040 20700
rect 6096 20698 6120 20700
rect 6176 20698 6200 20700
rect 6256 20698 6262 20700
rect 6016 20646 6018 20698
rect 6198 20646 6200 20698
rect 5954 20644 5960 20646
rect 6016 20644 6040 20646
rect 6096 20644 6120 20646
rect 6176 20644 6200 20646
rect 6256 20644 6262 20646
rect 5954 20635 6262 20644
rect 2908 20360 2960 20366
rect 2908 20302 2960 20308
rect 2920 20065 2948 20302
rect 7140 20292 7192 20298
rect 7140 20234 7192 20240
rect 7152 20201 7180 20234
rect 7138 20192 7194 20201
rect 6690 20156 6998 20165
rect 6690 20154 6696 20156
rect 6752 20154 6776 20156
rect 6832 20154 6856 20156
rect 6912 20154 6936 20156
rect 6992 20154 6998 20156
rect 6752 20102 6754 20154
rect 6934 20102 6936 20154
rect 7138 20127 7194 20136
rect 6690 20100 6696 20102
rect 6752 20100 6776 20102
rect 6832 20100 6856 20102
rect 6912 20100 6936 20102
rect 6992 20100 6998 20102
rect 6690 20091 6998 20100
rect 2906 20056 2962 20065
rect 2906 19991 2962 20000
rect 4932 19918 4984 19924
rect 4932 19860 4984 19866
rect 4944 19385 4972 19860
rect 5954 19612 6262 19621
rect 5954 19610 5960 19612
rect 6016 19610 6040 19612
rect 6096 19610 6120 19612
rect 6176 19610 6200 19612
rect 6256 19610 6262 19612
rect 6016 19558 6018 19610
rect 6198 19558 6200 19610
rect 5954 19556 5960 19558
rect 6016 19556 6040 19558
rect 6096 19556 6120 19558
rect 6176 19556 6200 19558
rect 6256 19556 6262 19558
rect 5954 19547 6262 19556
rect 4930 19376 4986 19385
rect 4930 19311 4986 19320
rect 6690 19068 6998 19077
rect 6690 19066 6696 19068
rect 6752 19066 6776 19068
rect 6832 19066 6856 19068
rect 6912 19066 6936 19068
rect 6992 19066 6998 19068
rect 6752 19014 6754 19066
rect 6934 19014 6936 19066
rect 6690 19012 6696 19014
rect 6752 19012 6776 19014
rect 6832 19012 6856 19014
rect 6912 19012 6936 19014
rect 6992 19012 6998 19014
rect 6690 19003 6998 19012
rect 5954 18524 6262 18533
rect 5954 18522 5960 18524
rect 6016 18522 6040 18524
rect 6096 18522 6120 18524
rect 6176 18522 6200 18524
rect 6256 18522 6262 18524
rect 6016 18470 6018 18522
rect 6198 18470 6200 18522
rect 5954 18468 5960 18470
rect 6016 18468 6040 18470
rect 6096 18468 6120 18470
rect 6176 18468 6200 18470
rect 6256 18468 6262 18470
rect 5954 18459 6262 18468
rect 5116 18218 5168 18224
rect 5116 18160 5168 18166
rect 5128 18025 5156 18160
rect 5114 18016 5170 18025
rect 5114 17951 5170 17960
rect 6690 17980 6998 17989
rect 6690 17978 6696 17980
rect 6752 17978 6776 17980
rect 6832 17978 6856 17980
rect 6912 17978 6936 17980
rect 6992 17978 6998 17980
rect 6752 17926 6754 17978
rect 6934 17926 6936 17978
rect 6690 17924 6696 17926
rect 6752 17924 6776 17926
rect 6832 17924 6856 17926
rect 6912 17924 6936 17926
rect 6992 17924 6998 17926
rect 6690 17915 6998 17924
rect 5954 17436 6262 17445
rect 5954 17434 5960 17436
rect 6016 17434 6040 17436
rect 6096 17434 6120 17436
rect 6176 17434 6200 17436
rect 6256 17434 6262 17436
rect 6016 17382 6018 17434
rect 6198 17382 6200 17434
rect 5954 17380 5960 17382
rect 6016 17380 6040 17382
rect 6096 17380 6120 17382
rect 6176 17380 6200 17382
rect 6256 17380 6262 17382
rect 5954 17371 6262 17380
rect 5208 17130 5260 17136
rect 5208 17072 5260 17078
rect 5220 16665 5248 17072
rect 7140 17028 7192 17034
rect 7140 16970 7192 16976
rect 7152 16937 7180 16970
rect 7138 16928 7194 16937
rect 6690 16892 6998 16901
rect 6690 16890 6696 16892
rect 6752 16890 6776 16892
rect 6832 16890 6856 16892
rect 6912 16890 6936 16892
rect 6992 16890 6998 16892
rect 6752 16838 6754 16890
rect 6934 16838 6936 16890
rect 7138 16863 7194 16872
rect 6690 16836 6696 16838
rect 6752 16836 6776 16838
rect 6832 16836 6856 16838
rect 6912 16836 6936 16838
rect 6992 16836 6998 16838
rect 6690 16827 6998 16836
rect 5206 16656 5262 16665
rect 5206 16591 5262 16600
rect 5954 16348 6262 16357
rect 5954 16346 5960 16348
rect 6016 16346 6040 16348
rect 6096 16346 6120 16348
rect 6176 16346 6200 16348
rect 6256 16346 6262 16348
rect 6016 16294 6018 16346
rect 6198 16294 6200 16346
rect 5954 16292 5960 16294
rect 6016 16292 6040 16294
rect 6096 16292 6120 16294
rect 6176 16292 6200 16294
rect 6256 16292 6262 16294
rect 5954 16283 6262 16292
rect 2908 16008 2960 16014
rect 2906 15976 2908 15985
rect 2960 15976 2962 15985
rect 2906 15911 2962 15920
rect 7600 15940 7652 15946
rect 7600 15882 7652 15888
rect 7612 15849 7640 15882
rect 7598 15840 7654 15849
rect 6690 15804 6998 15813
rect 6690 15802 6696 15804
rect 6752 15802 6776 15804
rect 6832 15802 6856 15804
rect 6912 15802 6936 15804
rect 6992 15802 6998 15804
rect 6752 15750 6754 15802
rect 6934 15750 6936 15802
rect 7598 15775 7654 15784
rect 6690 15748 6696 15750
rect 6752 15748 6776 15750
rect 6832 15748 6856 15750
rect 6912 15748 6936 15750
rect 6992 15748 6998 15750
rect 6690 15739 6998 15748
rect 5954 15260 6262 15269
rect 5954 15258 5960 15260
rect 6016 15258 6040 15260
rect 6096 15258 6120 15260
rect 6176 15258 6200 15260
rect 6256 15258 6262 15260
rect 6016 15206 6018 15258
rect 6198 15206 6200 15258
rect 5954 15204 5960 15206
rect 6016 15204 6040 15206
rect 6096 15204 6120 15206
rect 6176 15204 6200 15206
rect 6256 15204 6262 15206
rect 5954 15195 6262 15204
rect 2908 14920 2960 14926
rect 2908 14862 2960 14868
rect 2920 14625 2948 14862
rect 7600 14852 7652 14858
rect 7600 14794 7652 14800
rect 7612 14761 7640 14794
rect 7598 14752 7654 14761
rect 6690 14716 6998 14725
rect 6690 14714 6696 14716
rect 6752 14714 6776 14716
rect 6832 14714 6856 14716
rect 6912 14714 6936 14716
rect 6992 14714 6998 14716
rect 6752 14662 6754 14714
rect 6934 14662 6936 14714
rect 7598 14687 7654 14696
rect 6690 14660 6696 14662
rect 6752 14660 6776 14662
rect 6832 14660 6856 14662
rect 6912 14660 6936 14662
rect 6992 14660 6998 14662
rect 6690 14651 6998 14660
rect 2906 14616 2962 14625
rect 2906 14551 2962 14560
rect 4932 14478 4984 14484
rect 4932 14420 4984 14426
rect 4944 13945 4972 14420
rect 5668 14308 5720 14314
rect 5668 14250 5720 14256
rect 4930 13936 4986 13945
rect 4930 13871 4986 13880
rect 5680 13809 5708 14250
rect 5954 14172 6262 14181
rect 5954 14170 5960 14172
rect 6016 14170 6040 14172
rect 6096 14170 6120 14172
rect 6176 14170 6200 14172
rect 6256 14170 6262 14172
rect 6016 14118 6018 14170
rect 6198 14118 6200 14170
rect 5954 14116 5960 14118
rect 6016 14116 6040 14118
rect 6096 14116 6120 14118
rect 6176 14116 6200 14118
rect 6256 14116 6262 14118
rect 5954 14107 6262 14116
rect 5666 13800 5722 13809
rect 5666 13735 5722 13744
rect 6690 13628 6998 13637
rect 6690 13626 6696 13628
rect 6752 13626 6776 13628
rect 6832 13626 6856 13628
rect 6912 13626 6936 13628
rect 6992 13626 6998 13628
rect 6752 13574 6754 13626
rect 6934 13574 6936 13626
rect 6690 13572 6696 13574
rect 6752 13572 6776 13574
rect 6832 13572 6856 13574
rect 6912 13572 6936 13574
rect 6992 13572 6998 13574
rect 6690 13563 6998 13572
rect 5954 13084 6262 13093
rect 5954 13082 5960 13084
rect 6016 13082 6040 13084
rect 6096 13082 6120 13084
rect 6176 13082 6200 13084
rect 6256 13082 6262 13084
rect 6016 13030 6018 13082
rect 6198 13030 6200 13082
rect 5954 13028 5960 13030
rect 6016 13028 6040 13030
rect 6096 13028 6120 13030
rect 6176 13028 6200 13030
rect 6256 13028 6262 13030
rect 5954 13019 6262 13028
rect 6690 12540 6998 12549
rect 6690 12538 6696 12540
rect 6752 12538 6776 12540
rect 6832 12538 6856 12540
rect 6912 12538 6936 12540
rect 6992 12538 6998 12540
rect 6752 12486 6754 12538
rect 6934 12486 6936 12538
rect 6690 12484 6696 12486
rect 6752 12484 6776 12486
rect 6832 12484 6856 12486
rect 6912 12484 6936 12486
rect 6992 12484 6998 12486
rect 6690 12475 6998 12484
rect 5954 11996 6262 12005
rect 5954 11994 5960 11996
rect 6016 11994 6040 11996
rect 6096 11994 6120 11996
rect 6176 11994 6200 11996
rect 6256 11994 6262 11996
rect 6016 11942 6018 11994
rect 6198 11942 6200 11994
rect 5954 11940 5960 11942
rect 6016 11940 6040 11942
rect 6096 11940 6120 11942
rect 6176 11940 6200 11942
rect 6256 11940 6262 11942
rect 5954 11931 6262 11940
rect 6690 11452 6998 11461
rect 6690 11450 6696 11452
rect 6752 11450 6776 11452
rect 6832 11450 6856 11452
rect 6912 11450 6936 11452
rect 6992 11450 6998 11452
rect 6752 11398 6754 11450
rect 6934 11398 6936 11450
rect 6690 11396 6696 11398
rect 6752 11396 6776 11398
rect 6832 11396 6856 11398
rect 6912 11396 6936 11398
rect 6992 11396 6998 11398
rect 6690 11387 6998 11396
rect 5954 10908 6262 10917
rect 5954 10906 5960 10908
rect 6016 10906 6040 10908
rect 6096 10906 6120 10908
rect 6176 10906 6200 10908
rect 6256 10906 6262 10908
rect 6016 10854 6018 10906
rect 6198 10854 6200 10906
rect 5954 10852 5960 10854
rect 6016 10852 6040 10854
rect 6096 10852 6120 10854
rect 6176 10852 6200 10854
rect 6256 10852 6262 10854
rect 5954 10843 6262 10852
rect 7888 10545 7916 47162
rect 7874 10536 7930 10545
rect 7874 10471 7930 10480
rect 6690 10364 6998 10373
rect 6690 10362 6696 10364
rect 6752 10362 6776 10364
rect 6832 10362 6856 10364
rect 6912 10362 6936 10364
rect 6992 10362 6998 10364
rect 6752 10310 6754 10362
rect 6934 10310 6936 10362
rect 6690 10308 6696 10310
rect 6752 10308 6776 10310
rect 6832 10308 6856 10310
rect 6912 10308 6936 10310
rect 6992 10308 6998 10310
rect 6690 10299 6998 10308
rect 8164 10273 8192 47230
rect 8334 47191 8390 47200
rect 8348 10409 8376 47191
rect 8334 10400 8390 10409
rect 8334 10335 8390 10344
rect 8150 10264 8206 10273
rect 8150 10199 8206 10208
rect 5954 9820 6262 9829
rect 5954 9818 5960 9820
rect 6016 9818 6040 9820
rect 6096 9818 6120 9820
rect 6176 9818 6200 9820
rect 6256 9818 6262 9820
rect 6016 9766 6018 9818
rect 6198 9766 6200 9818
rect 5954 9764 5960 9766
rect 6016 9764 6040 9766
rect 6096 9764 6120 9766
rect 6176 9764 6200 9766
rect 6256 9764 6262 9766
rect 5954 9755 6262 9764
rect 6690 9276 6998 9285
rect 6690 9274 6696 9276
rect 6752 9274 6776 9276
rect 6832 9274 6856 9276
rect 6912 9274 6936 9276
rect 6992 9274 6998 9276
rect 6752 9222 6754 9274
rect 6934 9222 6936 9274
rect 6690 9220 6696 9222
rect 6752 9220 6776 9222
rect 6832 9220 6856 9222
rect 6912 9220 6936 9222
rect 6992 9220 6998 9222
rect 6690 9211 6998 9220
rect 5954 8732 6262 8741
rect 5954 8730 5960 8732
rect 6016 8730 6040 8732
rect 6096 8730 6120 8732
rect 6176 8730 6200 8732
rect 6256 8730 6262 8732
rect 6016 8678 6018 8730
rect 6198 8678 6200 8730
rect 5954 8676 5960 8678
rect 6016 8676 6040 8678
rect 6096 8676 6120 8678
rect 6176 8676 6200 8678
rect 6256 8676 6262 8678
rect 5954 8667 6262 8676
rect 8440 8505 8468 84319
rect 13672 84280 13724 84286
rect 9806 84248 9862 84257
rect 12226 84218 12608 84234
rect 13330 84228 13672 84234
rect 13330 84222 13724 84228
rect 12226 84212 12620 84218
rect 12226 84206 12568 84212
rect 9806 84183 9862 84192
rect 9624 62384 9676 62390
rect 9624 62326 9676 62332
rect 9636 61921 9664 62326
rect 9622 61912 9678 61921
rect 9622 61847 9678 61856
rect 9624 61092 9676 61098
rect 9624 61034 9676 61040
rect 9636 60833 9664 61034
rect 9622 60824 9678 60833
rect 9622 60759 9678 60768
rect 9820 48081 9848 84183
rect 13330 84206 13712 84222
rect 12568 84154 12620 84160
rect 31716 84150 31744 86602
rect 32084 84356 32112 88880
rect 33188 84356 33216 88880
rect 34292 84356 34320 88880
rect 35396 84356 35424 88880
rect 36500 84356 36528 88880
rect 37604 84356 37632 88880
rect 38382 88700 38690 88709
rect 38382 88698 38388 88700
rect 38444 88698 38468 88700
rect 38524 88698 38548 88700
rect 38604 88698 38628 88700
rect 38684 88698 38690 88700
rect 38444 88646 38446 88698
rect 38626 88646 38628 88698
rect 38382 88644 38388 88646
rect 38444 88644 38468 88646
rect 38524 88644 38548 88646
rect 38604 88644 38628 88646
rect 38684 88644 38690 88646
rect 38382 88635 38690 88644
rect 37722 88156 38030 88165
rect 37722 88154 37728 88156
rect 37784 88154 37808 88156
rect 37864 88154 37888 88156
rect 37944 88154 37968 88156
rect 38024 88154 38030 88156
rect 37784 88102 37786 88154
rect 37966 88102 37968 88154
rect 37722 88100 37728 88102
rect 37784 88100 37808 88102
rect 37864 88100 37888 88102
rect 37944 88100 37968 88102
rect 38024 88100 38030 88102
rect 37722 88091 38030 88100
rect 38382 87612 38690 87621
rect 38382 87610 38388 87612
rect 38444 87610 38468 87612
rect 38524 87610 38548 87612
rect 38604 87610 38628 87612
rect 38684 87610 38690 87612
rect 38444 87558 38446 87610
rect 38626 87558 38628 87610
rect 38382 87556 38388 87558
rect 38444 87556 38468 87558
rect 38524 87556 38548 87558
rect 38604 87556 38628 87558
rect 38684 87556 38690 87558
rect 38382 87547 38690 87556
rect 37722 87068 38030 87077
rect 37722 87066 37728 87068
rect 37784 87066 37808 87068
rect 37864 87066 37888 87068
rect 37944 87066 37968 87068
rect 38024 87066 38030 87068
rect 37784 87014 37786 87066
rect 37966 87014 37968 87066
rect 37722 87012 37728 87014
rect 37784 87012 37808 87014
rect 37864 87012 37888 87014
rect 37944 87012 37968 87014
rect 38024 87012 38030 87014
rect 37722 87003 38030 87012
rect 38382 86524 38690 86533
rect 38382 86522 38388 86524
rect 38444 86522 38468 86524
rect 38524 86522 38548 86524
rect 38604 86522 38628 86524
rect 38684 86522 38690 86524
rect 38444 86470 38446 86522
rect 38626 86470 38628 86522
rect 38382 86468 38388 86470
rect 38444 86468 38468 86470
rect 38524 86468 38548 86470
rect 38604 86468 38628 86470
rect 38684 86468 38690 86470
rect 38382 86459 38690 86468
rect 38800 85794 38828 88880
rect 38708 85766 38828 85794
rect 38708 84356 38736 85766
rect 39812 84356 39840 88880
rect 40916 84356 40944 88880
rect 42020 84356 42048 88880
rect 43124 84356 43152 88880
rect 44228 84356 44256 88880
rect 45332 84356 45360 88880
rect 48000 86734 48028 91800
rect 48644 88468 48672 91800
rect 49932 88939 49960 91800
rect 52508 88944 52536 91800
rect 53796 88944 53824 91800
rect 49920 88933 49972 88939
rect 52496 88938 52548 88944
rect 49920 88875 49972 88881
rect 50012 88904 50064 88910
rect 52496 88880 52548 88886
rect 53784 88938 53836 88944
rect 54440 88910 54468 91800
rect 55728 88944 55756 91800
rect 56372 89114 56400 91800
rect 57016 90354 57044 91800
rect 57016 90326 57136 90354
rect 56722 89244 57030 89253
rect 56722 89242 56728 89244
rect 56784 89242 56808 89244
rect 56864 89242 56888 89244
rect 56944 89242 56968 89244
rect 57024 89242 57030 89244
rect 56784 89190 56786 89242
rect 56966 89190 56968 89242
rect 56722 89188 56728 89190
rect 56784 89188 56808 89190
rect 56864 89188 56888 89190
rect 56944 89188 56968 89190
rect 57024 89188 57030 89190
rect 56722 89179 57030 89188
rect 56360 89108 56412 89114
rect 56360 89050 56412 89056
rect 57108 88944 57136 90326
rect 57660 89114 57688 91800
rect 57648 89108 57700 89114
rect 57648 89050 57700 89056
rect 55716 88938 55768 88944
rect 53784 88880 53836 88886
rect 54428 88904 54480 88910
rect 50012 88846 50064 88852
rect 55716 88880 55768 88886
rect 57096 88938 57148 88944
rect 58304 88910 58332 91800
rect 58948 88944 58976 91800
rect 60236 88944 60264 91800
rect 61524 88944 61552 91800
rect 62168 88978 62196 91800
rect 62156 88972 62208 88978
rect 58936 88938 58988 88944
rect 57096 88880 57148 88886
rect 58292 88904 58344 88910
rect 54428 88846 54480 88852
rect 58936 88880 58988 88886
rect 60224 88938 60276 88944
rect 60224 88880 60276 88886
rect 61512 88938 61564 88944
rect 62156 88914 62208 88920
rect 63456 88910 63484 91800
rect 64744 88910 64772 91800
rect 66032 88944 66060 91800
rect 66676 88944 66704 91800
rect 67964 89114 67992 91800
rect 69252 89114 69280 91800
rect 69896 89114 69924 91800
rect 71184 89114 71212 91800
rect 72472 89114 72500 91800
rect 73760 89114 73788 91800
rect 74404 89114 74432 91800
rect 75692 89402 75720 91800
rect 75600 89374 75720 89402
rect 75600 89114 75628 89374
rect 75722 89244 76030 89253
rect 75722 89242 75728 89244
rect 75784 89242 75808 89244
rect 75864 89242 75888 89244
rect 75944 89242 75968 89244
rect 76024 89242 76030 89244
rect 75784 89190 75786 89242
rect 75966 89190 75968 89242
rect 75722 89188 75728 89190
rect 75784 89188 75808 89190
rect 75864 89188 75888 89190
rect 75944 89188 75968 89190
rect 76024 89188 76030 89190
rect 75722 89179 76030 89188
rect 76980 89114 77008 91800
rect 77624 89114 77652 91800
rect 78912 89114 78940 91800
rect 80200 89114 80228 91800
rect 81488 89114 81516 91800
rect 82132 89114 82160 91800
rect 67952 89108 68004 89114
rect 67952 89050 68004 89056
rect 69240 89108 69292 89114
rect 69240 89050 69292 89056
rect 69884 89108 69936 89114
rect 69884 89050 69936 89056
rect 71172 89108 71224 89114
rect 71172 89050 71224 89056
rect 72460 89108 72512 89114
rect 72460 89050 72512 89056
rect 73748 89108 73800 89114
rect 73748 89050 73800 89056
rect 74392 89108 74444 89114
rect 74392 89050 74444 89056
rect 75588 89108 75640 89114
rect 75588 89050 75640 89056
rect 76968 89108 77020 89114
rect 76968 89050 77020 89056
rect 77612 89108 77664 89114
rect 77612 89050 77664 89056
rect 78900 89108 78952 89114
rect 78900 89050 78952 89056
rect 80188 89108 80240 89114
rect 80188 89050 80240 89056
rect 81476 89108 81528 89114
rect 81476 89050 81528 89056
rect 82120 89108 82172 89114
rect 82120 89050 82172 89056
rect 66020 88938 66072 88944
rect 61512 88880 61564 88886
rect 63444 88904 63496 88910
rect 58292 88846 58344 88852
rect 63444 88846 63496 88852
rect 64732 88904 64784 88910
rect 66020 88880 66072 88886
rect 66664 88938 66716 88944
rect 66664 88880 66716 88886
rect 68044 88938 68096 88944
rect 68044 88880 68096 88886
rect 69424 88938 69476 88944
rect 69424 88880 69476 88886
rect 70252 88938 70304 88944
rect 70252 88880 70304 88886
rect 71356 88938 71408 88944
rect 71356 88880 71408 88886
rect 72460 88938 72512 88944
rect 72460 88880 72512 88886
rect 73564 88938 73616 88944
rect 73564 88880 73616 88886
rect 74668 88938 74720 88944
rect 74668 88880 74720 88886
rect 75496 88938 75548 88944
rect 75496 88880 75548 88886
rect 76876 88938 76928 88944
rect 76876 88880 76928 88886
rect 77980 88938 78032 88944
rect 77980 88880 78032 88886
rect 79084 88938 79136 88944
rect 79084 88880 79136 88886
rect 80280 88938 80332 88944
rect 80280 88880 80332 88886
rect 81292 88938 81344 88944
rect 81292 88880 81344 88886
rect 82396 88938 82448 88944
rect 82396 88880 82448 88886
rect 64732 88846 64784 88852
rect 48632 88462 48684 88468
rect 48632 88404 48684 88410
rect 49644 88428 49696 88434
rect 49644 88370 49696 88376
rect 49656 87380 49684 88370
rect 49276 87374 49328 87380
rect 49276 87316 49328 87322
rect 49644 87374 49696 87380
rect 49644 87316 49696 87322
rect 47988 86728 48040 86734
rect 47988 86670 48040 86676
rect 49288 84506 49316 87316
rect 50024 86763 50052 88846
rect 52772 88836 52824 88842
rect 52772 88778 52824 88784
rect 54152 88836 54204 88842
rect 54152 88778 54204 88784
rect 54796 88836 54848 88842
rect 54796 88778 54848 88784
rect 55992 88836 56044 88842
rect 55992 88778 56044 88784
rect 57096 88836 57148 88842
rect 57096 88778 57148 88784
rect 58384 88836 58436 88842
rect 58384 88778 58436 88784
rect 59304 88836 59356 88842
rect 59304 88778 59356 88784
rect 60316 88836 60368 88842
rect 60316 88778 60368 88784
rect 61420 88836 61472 88842
rect 61420 88778 61472 88784
rect 62524 88836 62576 88842
rect 62524 88778 62576 88784
rect 63720 88836 63772 88842
rect 63720 88778 63772 88784
rect 65100 88836 65152 88842
rect 65100 88778 65152 88784
rect 65836 88836 65888 88842
rect 65836 88778 65888 88784
rect 66940 88836 66992 88842
rect 66940 88778 66992 88784
rect 50012 86757 50064 86763
rect 50012 86699 50064 86705
rect 49242 84478 49316 84506
rect 49242 84370 49270 84478
rect 48920 84356 49270 84370
rect 48920 84342 49256 84356
rect 48920 84218 48948 84342
rect 50024 84286 50052 86699
rect 52784 85794 52812 88778
rect 54164 85794 54192 88778
rect 52692 85766 52812 85794
rect 54072 85766 54192 85794
rect 52692 84370 52720 85766
rect 54072 84370 54100 85766
rect 54808 84642 54836 88778
rect 56004 85794 56032 88778
rect 56722 88156 57030 88165
rect 56722 88154 56728 88156
rect 56784 88154 56808 88156
rect 56864 88154 56888 88156
rect 56944 88154 56968 88156
rect 57024 88154 57030 88156
rect 56784 88102 56786 88154
rect 56966 88102 56968 88154
rect 56722 88100 56728 88102
rect 56784 88100 56808 88102
rect 56864 88100 56888 88102
rect 56944 88100 56968 88102
rect 57024 88100 57030 88102
rect 56722 88091 57030 88100
rect 56722 87068 57030 87077
rect 56722 87066 56728 87068
rect 56784 87066 56808 87068
rect 56864 87066 56888 87068
rect 56944 87066 56968 87068
rect 57024 87066 57030 87068
rect 56784 87014 56786 87066
rect 56966 87014 56968 87066
rect 56722 87012 56728 87014
rect 56784 87012 56808 87014
rect 56864 87012 56888 87014
rect 56944 87012 56968 87014
rect 57024 87012 57030 87014
rect 56722 87003 57030 87012
rect 55912 85766 56032 85794
rect 55912 84642 55940 85766
rect 52568 84342 52720 84370
rect 53672 84342 54100 84370
rect 54762 84614 54836 84642
rect 55866 84614 55940 84642
rect 54762 84356 54790 84614
rect 55866 84356 55894 84614
rect 57108 84370 57136 88778
rect 57382 88700 57690 88709
rect 57382 88698 57388 88700
rect 57444 88698 57468 88700
rect 57524 88698 57548 88700
rect 57604 88698 57628 88700
rect 57684 88698 57690 88700
rect 57444 88646 57446 88698
rect 57626 88646 57628 88698
rect 57382 88644 57388 88646
rect 57444 88644 57468 88646
rect 57524 88644 57548 88646
rect 57604 88644 57628 88646
rect 57684 88644 57690 88646
rect 57382 88635 57690 88644
rect 57382 87612 57690 87621
rect 57382 87610 57388 87612
rect 57444 87610 57468 87612
rect 57524 87610 57548 87612
rect 57604 87610 57628 87612
rect 57684 87610 57690 87612
rect 57444 87558 57446 87610
rect 57626 87558 57628 87610
rect 57382 87556 57388 87558
rect 57444 87556 57468 87558
rect 57524 87556 57548 87558
rect 57604 87556 57628 87558
rect 57684 87556 57690 87558
rect 57382 87547 57690 87556
rect 57382 86524 57690 86533
rect 57382 86522 57388 86524
rect 57444 86522 57468 86524
rect 57524 86522 57548 86524
rect 57604 86522 57628 86524
rect 57684 86522 57690 86524
rect 57444 86470 57446 86522
rect 57626 86470 57628 86522
rect 57382 86468 57388 86470
rect 57444 86468 57468 86470
rect 57524 86468 57548 86470
rect 57604 86468 57628 86470
rect 57684 86468 57690 86470
rect 57382 86459 57690 86468
rect 58396 84370 58424 88778
rect 59316 85794 59344 88778
rect 59224 85766 59344 85794
rect 59224 84642 59252 85766
rect 60328 84642 60356 88778
rect 61432 84642 61460 88778
rect 62536 84642 62564 88778
rect 56984 84342 57136 84370
rect 58088 84342 58424 84370
rect 59178 84614 59252 84642
rect 60282 84614 60356 84642
rect 61386 84614 61460 84642
rect 62490 84614 62564 84642
rect 59178 84356 59206 84614
rect 60282 84356 60310 84614
rect 61386 84356 61414 84614
rect 62490 84356 62518 84614
rect 63732 84370 63760 88778
rect 65112 84370 65140 88778
rect 65848 84642 65876 88778
rect 66952 84642 66980 88778
rect 68056 84642 68084 88880
rect 63608 84342 63760 84370
rect 64712 84342 65140 84370
rect 65802 84614 65876 84642
rect 66906 84614 66980 84642
rect 68010 84614 68084 84642
rect 65802 84356 65830 84614
rect 66906 84356 66934 84614
rect 68010 84356 68038 84614
rect 69436 84370 69464 88880
rect 70264 84642 70292 88880
rect 71368 84642 71396 88880
rect 72472 84642 72500 88880
rect 73576 84642 73604 88880
rect 74680 84642 74708 88880
rect 69128 84342 69464 84370
rect 70218 84614 70292 84642
rect 71322 84614 71396 84642
rect 72426 84614 72500 84642
rect 73530 84614 73604 84642
rect 74634 84614 74708 84642
rect 70218 84356 70246 84614
rect 71322 84356 71350 84614
rect 72426 84356 72454 84614
rect 73530 84356 73558 84614
rect 74634 84356 74662 84614
rect 75508 84370 75536 88880
rect 76382 88700 76690 88709
rect 76382 88698 76388 88700
rect 76444 88698 76468 88700
rect 76524 88698 76548 88700
rect 76604 88698 76628 88700
rect 76684 88698 76690 88700
rect 76444 88646 76446 88698
rect 76626 88646 76628 88698
rect 76382 88644 76388 88646
rect 76444 88644 76468 88646
rect 76524 88644 76548 88646
rect 76604 88644 76628 88646
rect 76684 88644 76690 88646
rect 76382 88635 76690 88644
rect 75722 88156 76030 88165
rect 75722 88154 75728 88156
rect 75784 88154 75808 88156
rect 75864 88154 75888 88156
rect 75944 88154 75968 88156
rect 76024 88154 76030 88156
rect 75784 88102 75786 88154
rect 75966 88102 75968 88154
rect 75722 88100 75728 88102
rect 75784 88100 75808 88102
rect 75864 88100 75888 88102
rect 75944 88100 75968 88102
rect 76024 88100 76030 88102
rect 75722 88091 76030 88100
rect 76382 87612 76690 87621
rect 76382 87610 76388 87612
rect 76444 87610 76468 87612
rect 76524 87610 76548 87612
rect 76604 87610 76628 87612
rect 76684 87610 76690 87612
rect 76444 87558 76446 87610
rect 76626 87558 76628 87610
rect 76382 87556 76388 87558
rect 76444 87556 76468 87558
rect 76524 87556 76548 87558
rect 76604 87556 76628 87558
rect 76684 87556 76690 87558
rect 76382 87547 76690 87556
rect 75722 87068 76030 87077
rect 75722 87066 75728 87068
rect 75784 87066 75808 87068
rect 75864 87066 75888 87068
rect 75944 87066 75968 87068
rect 76024 87066 76030 87068
rect 75784 87014 75786 87066
rect 75966 87014 75968 87066
rect 75722 87012 75728 87014
rect 75784 87012 75808 87014
rect 75864 87012 75888 87014
rect 75944 87012 75968 87014
rect 76024 87012 76030 87014
rect 75722 87003 76030 87012
rect 76382 86524 76690 86533
rect 76382 86522 76388 86524
rect 76444 86522 76468 86524
rect 76524 86522 76548 86524
rect 76604 86522 76628 86524
rect 76684 86522 76690 86524
rect 76444 86470 76446 86522
rect 76626 86470 76628 86522
rect 76382 86468 76388 86470
rect 76444 86468 76468 86470
rect 76524 86468 76548 86470
rect 76604 86468 76628 86470
rect 76684 86468 76690 86470
rect 76382 86459 76690 86468
rect 76888 84642 76916 88880
rect 77992 84642 78020 88880
rect 79096 84642 79124 88880
rect 76842 84614 76916 84642
rect 77946 84614 78020 84642
rect 79050 84614 79124 84642
rect 75508 84342 75752 84370
rect 76842 84356 76870 84614
rect 77946 84356 77974 84614
rect 79050 84356 79078 84614
rect 80292 84370 80320 88880
rect 81304 84642 81332 88880
rect 82408 84642 82436 88880
rect 83684 87340 83736 87346
rect 83684 87282 83736 87288
rect 80168 84342 80320 84370
rect 81258 84614 81332 84642
rect 82362 84614 82436 84642
rect 81258 84356 81286 84614
rect 82362 84356 82390 84614
rect 50012 84280 50064 84286
rect 51436 84248 51492 84257
rect 50064 84228 50360 84234
rect 50012 84222 50360 84228
rect 48908 84212 48960 84218
rect 50024 84206 50360 84222
rect 51436 84183 51492 84192
rect 48908 84154 48960 84160
rect 11280 84144 11332 84150
rect 11122 84092 11280 84098
rect 11122 84086 11332 84092
rect 31704 84144 31756 84150
rect 31704 84086 31756 84092
rect 47804 84144 47856 84150
rect 47856 84092 48152 84098
rect 47804 84086 48152 84092
rect 11122 84070 11320 84086
rect 47816 84070 48152 84086
rect 9806 48072 9862 48081
rect 9806 48007 9862 48016
rect 11122 48072 11178 48081
rect 11122 48007 11178 48016
rect 12240 47362 12268 47500
rect 12228 47356 12280 47362
rect 12228 47298 12280 47304
rect 12240 47242 12268 47298
rect 13344 47265 13372 47500
rect 14448 47294 14476 47500
rect 14436 47288 14488 47294
rect 12212 47226 12268 47242
rect 12200 47220 12268 47226
rect 12252 47214 12268 47220
rect 13330 47256 13386 47265
rect 15552 47276 15580 47500
rect 16656 47276 16684 47500
rect 17760 47276 17788 47500
rect 14436 47230 14488 47236
rect 15524 47248 15580 47276
rect 16628 47248 16684 47276
rect 17732 47248 17788 47276
rect 13330 47191 13386 47200
rect 12200 47162 12252 47168
rect 11004 47152 11056 47158
rect 11004 47094 11056 47100
rect 9806 46848 9862 46857
rect 9806 46783 9862 46792
rect 9624 19748 9676 19754
rect 9624 19690 9676 19696
rect 9636 19081 9664 19690
rect 9622 19072 9678 19081
rect 9622 19007 9678 19016
rect 9624 18252 9676 18258
rect 9624 18194 9676 18200
rect 9636 17993 9664 18194
rect 9622 17984 9678 17993
rect 9622 17919 9678 17928
rect 9820 10681 9848 46783
rect 11016 46750 11044 47094
rect 14144 46954 14434 46970
rect 15524 46956 15552 47248
rect 16628 46956 16656 47248
rect 17732 46956 17760 47248
rect 18864 47242 18892 47500
rect 19968 47242 19996 47500
rect 21072 47242 21100 47500
rect 22176 47242 22204 47500
rect 23280 47242 23308 47500
rect 24384 47242 24412 47500
rect 25488 47242 25516 47500
rect 26592 47242 26620 47500
rect 27696 47242 27724 47500
rect 28800 47242 28828 47500
rect 29904 47242 29932 47500
rect 31008 47242 31036 47500
rect 32112 47242 32140 47500
rect 33216 47242 33244 47500
rect 34320 47242 34348 47500
rect 35424 47242 35452 47500
rect 36528 47242 36556 47500
rect 37632 47242 37660 47500
rect 38736 47242 38764 47500
rect 39840 47242 39868 47500
rect 40944 47242 40972 47500
rect 42048 47242 42076 47500
rect 43152 47242 43180 47500
rect 44256 47242 44284 47500
rect 45360 47242 45388 47500
rect 18836 47214 18892 47242
rect 19940 47214 19996 47242
rect 21044 47214 21100 47242
rect 22148 47214 22204 47242
rect 23252 47214 23308 47242
rect 24356 47214 24412 47242
rect 25460 47214 25516 47242
rect 26564 47214 26620 47242
rect 27668 47214 27724 47242
rect 28772 47214 28828 47242
rect 29876 47214 29932 47242
rect 30980 47214 31036 47242
rect 32084 47214 32140 47242
rect 33188 47214 33244 47242
rect 34292 47214 34348 47242
rect 35396 47214 35452 47242
rect 36500 47214 36556 47242
rect 37604 47214 37660 47242
rect 38708 47214 38764 47242
rect 39812 47214 39868 47242
rect 40916 47214 40972 47242
rect 42020 47214 42076 47242
rect 43124 47214 43180 47242
rect 44228 47214 44284 47242
rect 45332 47214 45388 47242
rect 48138 47242 48166 47500
rect 49242 47362 49270 47500
rect 49230 47356 49282 47362
rect 49230 47298 49282 47304
rect 50346 47265 50374 47500
rect 51450 47362 51478 47500
rect 51438 47356 51490 47362
rect 51438 47298 51490 47304
rect 50332 47256 50388 47265
rect 48138 47226 48212 47242
rect 48138 47220 48224 47226
rect 48138 47214 48172 47220
rect 18836 46956 18864 47214
rect 19940 46956 19968 47214
rect 21044 46956 21072 47214
rect 22148 46956 22176 47214
rect 23252 46956 23280 47214
rect 24356 46956 24384 47214
rect 25460 46956 25488 47214
rect 26564 46956 26592 47214
rect 27668 46956 27696 47214
rect 28772 46956 28800 47214
rect 29876 46956 29904 47214
rect 30980 46956 31008 47214
rect 32084 46956 32112 47214
rect 33188 46956 33216 47214
rect 34292 46956 34320 47214
rect 35396 46956 35424 47214
rect 36500 46956 36528 47214
rect 37604 46956 37632 47214
rect 38708 46956 38736 47214
rect 39812 46956 39840 47214
rect 40916 46956 40944 47214
rect 42020 46956 42048 47214
rect 43124 46956 43152 47214
rect 44228 46956 44256 47214
rect 45332 46956 45360 47214
rect 50332 47191 50388 47200
rect 48172 47162 48224 47168
rect 52554 46956 52582 47500
rect 53658 46956 53686 47500
rect 54762 46956 54790 47500
rect 55866 46956 55894 47500
rect 56970 46956 56998 47500
rect 58074 46956 58102 47500
rect 59178 46956 59206 47500
rect 60282 46956 60310 47500
rect 61386 46956 61414 47500
rect 62490 46956 62518 47500
rect 63594 46956 63622 47500
rect 64698 46956 64726 47500
rect 65802 46956 65830 47500
rect 66906 46956 66934 47500
rect 68010 46956 68038 47500
rect 69114 46956 69142 47500
rect 70218 46956 70246 47500
rect 71322 46956 71350 47500
rect 72426 46956 72454 47500
rect 73530 46956 73558 47500
rect 74634 46956 74662 47500
rect 75738 46956 75766 47500
rect 76842 46956 76870 47500
rect 77946 46956 77974 47500
rect 79050 46956 79078 47500
rect 80154 46956 80182 47500
rect 81258 46956 81286 47500
rect 82362 46956 82390 47500
rect 14132 46948 14434 46954
rect 14184 46942 14434 46948
rect 14132 46890 14184 46896
rect 13580 46880 13632 46886
rect 12226 46818 12516 46834
rect 13330 46828 13580 46834
rect 13330 46822 13632 46828
rect 50196 46880 50248 46886
rect 51436 46848 51492 46857
rect 50248 46828 50696 46834
rect 50196 46822 50696 46828
rect 12226 46812 12528 46818
rect 12226 46806 12476 46812
rect 13330 46806 13620 46822
rect 50208 46818 50696 46822
rect 49092 46812 49144 46818
rect 12476 46754 12528 46760
rect 50208 46812 50708 46818
rect 50208 46806 50656 46812
rect 49092 46754 49144 46760
rect 51436 46783 51492 46792
rect 50656 46754 50708 46760
rect 11004 46744 11056 46750
rect 47804 46744 47856 46750
rect 11056 46692 11122 46698
rect 11004 46686 11122 46692
rect 49104 46698 49132 46754
rect 83696 46750 83724 87282
rect 87098 87068 87406 87077
rect 87098 87066 87104 87068
rect 87160 87066 87184 87068
rect 87240 87066 87264 87068
rect 87320 87066 87344 87068
rect 87400 87066 87406 87068
rect 87160 87014 87162 87066
rect 87342 87014 87344 87066
rect 87098 87012 87104 87014
rect 87160 87012 87184 87014
rect 87240 87012 87264 87014
rect 87320 87012 87344 87014
rect 87400 87012 87406 87014
rect 87098 87003 87406 87012
rect 84052 86728 84104 86734
rect 84052 86670 84104 86676
rect 84064 46818 84092 86670
rect 87834 86524 88142 86533
rect 87834 86522 87840 86524
rect 87896 86522 87920 86524
rect 87976 86522 88000 86524
rect 88056 86522 88080 86524
rect 88136 86522 88142 86524
rect 87896 86470 87898 86522
rect 88078 86470 88080 86522
rect 87834 86468 87840 86470
rect 87896 86468 87920 86470
rect 87976 86468 88000 86470
rect 88056 86468 88080 86470
rect 88136 86468 88142 86470
rect 87834 86459 88142 86468
rect 87098 85980 87406 85989
rect 87098 85978 87104 85980
rect 87160 85978 87184 85980
rect 87240 85978 87264 85980
rect 87320 85978 87344 85980
rect 87400 85978 87406 85980
rect 87160 85926 87162 85978
rect 87342 85926 87344 85978
rect 87098 85924 87104 85926
rect 87160 85924 87184 85926
rect 87240 85924 87264 85926
rect 87320 85924 87344 85926
rect 87400 85924 87406 85926
rect 87098 85915 87406 85924
rect 87834 85436 88142 85445
rect 87834 85434 87840 85436
rect 87896 85434 87920 85436
rect 87976 85434 88000 85436
rect 88056 85434 88080 85436
rect 88136 85434 88142 85436
rect 87896 85382 87898 85434
rect 88078 85382 88080 85434
rect 87834 85380 87840 85382
rect 87896 85380 87920 85382
rect 87976 85380 88000 85382
rect 88056 85380 88080 85382
rect 88136 85380 88142 85382
rect 87834 85371 88142 85380
rect 87098 84892 87406 84901
rect 87098 84890 87104 84892
rect 87160 84890 87184 84892
rect 87240 84890 87264 84892
rect 87320 84890 87344 84892
rect 87400 84890 87406 84892
rect 87160 84838 87162 84890
rect 87342 84838 87344 84890
rect 87098 84836 87104 84838
rect 87160 84836 87184 84838
rect 87240 84836 87264 84838
rect 87320 84836 87344 84838
rect 87400 84836 87406 84838
rect 87098 84827 87406 84836
rect 87834 84348 88142 84357
rect 87834 84346 87840 84348
rect 87896 84346 87920 84348
rect 87976 84346 88000 84348
rect 88056 84346 88080 84348
rect 88136 84346 88142 84348
rect 87896 84294 87898 84346
rect 88078 84294 88080 84346
rect 87834 84292 87840 84294
rect 87896 84292 87920 84294
rect 87976 84292 88000 84294
rect 88056 84292 88080 84294
rect 88136 84292 88142 84294
rect 87834 84283 88142 84292
rect 87098 83804 87406 83813
rect 87098 83802 87104 83804
rect 87160 83802 87184 83804
rect 87240 83802 87264 83804
rect 87320 83802 87344 83804
rect 87400 83802 87406 83804
rect 87160 83750 87162 83802
rect 87342 83750 87344 83802
rect 87098 83748 87104 83750
rect 87160 83748 87184 83750
rect 87240 83748 87264 83750
rect 87320 83748 87344 83750
rect 87400 83748 87406 83750
rect 87098 83739 87406 83748
rect 87834 83260 88142 83269
rect 87834 83258 87840 83260
rect 87896 83258 87920 83260
rect 87976 83258 88000 83260
rect 88056 83258 88080 83260
rect 88136 83258 88142 83260
rect 87896 83206 87898 83258
rect 88078 83206 88080 83258
rect 87834 83204 87840 83206
rect 87896 83204 87920 83206
rect 87976 83204 88000 83206
rect 88056 83204 88080 83206
rect 88136 83204 88142 83206
rect 87834 83195 88142 83204
rect 87098 82716 87406 82725
rect 87098 82714 87104 82716
rect 87160 82714 87184 82716
rect 87240 82714 87264 82716
rect 87320 82714 87344 82716
rect 87400 82714 87406 82716
rect 87160 82662 87162 82714
rect 87342 82662 87344 82714
rect 87098 82660 87104 82662
rect 87160 82660 87184 82662
rect 87240 82660 87264 82662
rect 87320 82660 87344 82662
rect 87400 82660 87406 82662
rect 87098 82651 87406 82660
rect 87834 82172 88142 82181
rect 87834 82170 87840 82172
rect 87896 82170 87920 82172
rect 87976 82170 88000 82172
rect 88056 82170 88080 82172
rect 88136 82170 88142 82172
rect 87896 82118 87898 82170
rect 88078 82118 88080 82170
rect 87834 82116 87840 82118
rect 87896 82116 87920 82118
rect 87976 82116 88000 82118
rect 88056 82116 88080 82118
rect 88136 82116 88142 82118
rect 87834 82107 88142 82116
rect 87098 81628 87406 81637
rect 87098 81626 87104 81628
rect 87160 81626 87184 81628
rect 87240 81626 87264 81628
rect 87320 81626 87344 81628
rect 87400 81626 87406 81628
rect 87160 81574 87162 81626
rect 87342 81574 87344 81626
rect 87098 81572 87104 81574
rect 87160 81572 87184 81574
rect 87240 81572 87264 81574
rect 87320 81572 87344 81574
rect 87400 81572 87406 81574
rect 87098 81563 87406 81572
rect 87834 81084 88142 81093
rect 87834 81082 87840 81084
rect 87896 81082 87920 81084
rect 87976 81082 88000 81084
rect 88056 81082 88080 81084
rect 88136 81082 88142 81084
rect 87896 81030 87898 81082
rect 88078 81030 88080 81082
rect 87834 81028 87840 81030
rect 87896 81028 87920 81030
rect 87976 81028 88000 81030
rect 88056 81028 88080 81030
rect 88136 81028 88142 81030
rect 87834 81019 88142 81028
rect 88652 80812 88704 80818
rect 88652 80754 88704 80760
rect 84328 80676 84380 80682
rect 84328 80618 84380 80624
rect 84340 80449 84368 80618
rect 88664 80585 88692 80754
rect 88650 80576 88706 80585
rect 87098 80540 87406 80549
rect 87098 80538 87104 80540
rect 87160 80538 87184 80540
rect 87240 80538 87264 80540
rect 87320 80538 87344 80540
rect 87400 80538 87406 80540
rect 87160 80486 87162 80538
rect 87342 80486 87344 80538
rect 88650 80511 88706 80520
rect 87098 80484 87104 80486
rect 87160 80484 87184 80486
rect 87240 80484 87264 80486
rect 87320 80484 87344 80486
rect 87400 80484 87406 80486
rect 87098 80475 87406 80484
rect 84326 80440 84382 80449
rect 84326 80375 84382 80384
rect 87834 79996 88142 80005
rect 87834 79994 87840 79996
rect 87896 79994 87920 79996
rect 87976 79994 88000 79996
rect 88056 79994 88080 79996
rect 88136 79994 88142 79996
rect 87896 79942 87898 79994
rect 88078 79942 88080 79994
rect 87834 79940 87840 79942
rect 87896 79940 87920 79942
rect 87976 79940 88000 79942
rect 88056 79940 88080 79942
rect 88136 79940 88142 79942
rect 87834 79931 88142 79940
rect 88652 79758 88704 79764
rect 88652 79700 88704 79706
rect 84328 79588 84380 79594
rect 84328 79530 84380 79536
rect 84340 79361 84368 79530
rect 87098 79452 87406 79461
rect 87098 79450 87104 79452
rect 87160 79450 87184 79452
rect 87240 79450 87264 79452
rect 87320 79450 87344 79452
rect 87400 79450 87406 79452
rect 87160 79398 87162 79450
rect 87342 79398 87344 79450
rect 87098 79396 87104 79398
rect 87160 79396 87184 79398
rect 87240 79396 87264 79398
rect 87320 79396 87344 79398
rect 87400 79396 87406 79398
rect 87098 79387 87406 79396
rect 84326 79352 84382 79361
rect 84326 79287 84382 79296
rect 88664 79225 88692 79700
rect 88650 79216 88706 79225
rect 88650 79151 88706 79160
rect 87834 78908 88142 78917
rect 87834 78906 87840 78908
rect 87896 78906 87920 78908
rect 87976 78906 88000 78908
rect 88056 78906 88080 78908
rect 88136 78906 88142 78908
rect 87896 78854 87898 78906
rect 88078 78854 88080 78906
rect 87834 78852 87840 78854
rect 87896 78852 87920 78854
rect 87976 78852 88000 78854
rect 88056 78852 88080 78854
rect 88136 78852 88142 78854
rect 87834 78843 88142 78852
rect 88652 78670 88704 78676
rect 88652 78612 88704 78618
rect 88664 78545 88692 78612
rect 88650 78536 88706 78545
rect 84328 78500 84380 78506
rect 88650 78471 88706 78480
rect 84328 78442 84380 78448
rect 84340 78273 84368 78442
rect 87098 78364 87406 78373
rect 87098 78362 87104 78364
rect 87160 78362 87184 78364
rect 87240 78362 87264 78364
rect 87320 78362 87344 78364
rect 87400 78362 87406 78364
rect 87160 78310 87162 78362
rect 87342 78310 87344 78362
rect 87098 78308 87104 78310
rect 87160 78308 87184 78310
rect 87240 78308 87264 78310
rect 87320 78308 87344 78310
rect 87400 78308 87406 78310
rect 87098 78299 87406 78308
rect 84326 78264 84382 78273
rect 84326 78199 84382 78208
rect 87834 77820 88142 77829
rect 87834 77818 87840 77820
rect 87896 77818 87920 77820
rect 87976 77818 88000 77820
rect 88056 77818 88080 77820
rect 88136 77818 88142 77820
rect 87896 77766 87898 77818
rect 88078 77766 88080 77818
rect 87834 77764 87840 77766
rect 87896 77764 87920 77766
rect 87976 77764 88000 77766
rect 88056 77764 88080 77766
rect 88136 77764 88142 77766
rect 87834 77755 88142 77764
rect 90032 77616 90084 77622
rect 90032 77558 90084 77564
rect 84328 77480 84380 77486
rect 84328 77422 84380 77428
rect 84340 77185 84368 77422
rect 87098 77276 87406 77285
rect 87098 77274 87104 77276
rect 87160 77274 87184 77276
rect 87240 77274 87264 77276
rect 87320 77274 87344 77276
rect 87400 77274 87406 77276
rect 87160 77222 87162 77274
rect 87342 77222 87344 77274
rect 87098 77220 87104 77222
rect 87160 77220 87184 77222
rect 87240 77220 87264 77222
rect 87320 77220 87344 77222
rect 87400 77220 87406 77222
rect 87098 77211 87406 77220
rect 90044 77185 90072 77558
rect 84326 77176 84382 77185
rect 84326 77111 84382 77120
rect 90030 77176 90086 77185
rect 90030 77111 90086 77120
rect 87834 76732 88142 76741
rect 87834 76730 87840 76732
rect 87896 76730 87920 76732
rect 87976 76730 88000 76732
rect 88056 76730 88080 76732
rect 88136 76730 88142 76732
rect 87896 76678 87898 76730
rect 88078 76678 88080 76730
rect 87834 76676 87840 76678
rect 87896 76676 87920 76678
rect 87976 76676 88000 76678
rect 88056 76676 88080 76678
rect 88136 76676 88142 76678
rect 87834 76667 88142 76676
rect 87098 76188 87406 76197
rect 87098 76186 87104 76188
rect 87160 76186 87184 76188
rect 87240 76186 87264 76188
rect 87320 76186 87344 76188
rect 87400 76186 87406 76188
rect 87160 76134 87162 76186
rect 87342 76134 87344 76186
rect 87098 76132 87104 76134
rect 87160 76132 87184 76134
rect 87240 76132 87264 76134
rect 87320 76132 87344 76134
rect 87400 76132 87406 76134
rect 87098 76123 87406 76132
rect 84326 76020 84382 76029
rect 84326 75955 84328 75964
rect 84380 75955 84382 75964
rect 84328 75926 84380 75932
rect 88744 75848 88796 75854
rect 88742 75816 88744 75825
rect 88796 75816 88798 75825
rect 88742 75751 88798 75760
rect 87834 75644 88142 75653
rect 87834 75642 87840 75644
rect 87896 75642 87920 75644
rect 87976 75642 88000 75644
rect 88056 75642 88080 75644
rect 88136 75642 88142 75644
rect 87896 75590 87898 75642
rect 88078 75590 88080 75642
rect 87834 75588 87840 75590
rect 87896 75588 87920 75590
rect 87976 75588 88000 75590
rect 88056 75588 88080 75590
rect 88136 75588 88142 75590
rect 87834 75579 88142 75588
rect 88560 75440 88612 75446
rect 88560 75382 88612 75388
rect 84328 75304 84380 75310
rect 84328 75246 84380 75252
rect 84340 75009 84368 75246
rect 88572 75145 88600 75382
rect 88558 75136 88614 75145
rect 87098 75100 87406 75109
rect 87098 75098 87104 75100
rect 87160 75098 87184 75100
rect 87240 75098 87264 75100
rect 87320 75098 87344 75100
rect 87400 75098 87406 75100
rect 87160 75046 87162 75098
rect 87342 75046 87344 75098
rect 88558 75071 88614 75080
rect 87098 75044 87104 75046
rect 87160 75044 87184 75046
rect 87240 75044 87264 75046
rect 87320 75044 87344 75046
rect 87400 75044 87406 75046
rect 87098 75035 87406 75044
rect 84326 75000 84382 75009
rect 84326 74935 84382 74944
rect 87834 74556 88142 74565
rect 87834 74554 87840 74556
rect 87896 74554 87920 74556
rect 87976 74554 88000 74556
rect 88056 74554 88080 74556
rect 88136 74554 88142 74556
rect 87896 74502 87898 74554
rect 88078 74502 88080 74554
rect 87834 74500 87840 74502
rect 87896 74500 87920 74502
rect 87976 74500 88000 74502
rect 88056 74500 88080 74502
rect 88136 74500 88142 74502
rect 87834 74491 88142 74500
rect 88560 74352 88612 74358
rect 88560 74294 88612 74300
rect 84328 74216 84380 74222
rect 84328 74158 84380 74164
rect 84340 73921 84368 74158
rect 87098 74012 87406 74021
rect 87098 74010 87104 74012
rect 87160 74010 87184 74012
rect 87240 74010 87264 74012
rect 87320 74010 87344 74012
rect 87400 74010 87406 74012
rect 87160 73958 87162 74010
rect 87342 73958 87344 74010
rect 87098 73956 87104 73958
rect 87160 73956 87184 73958
rect 87240 73956 87264 73958
rect 87320 73956 87344 73958
rect 87400 73956 87406 73958
rect 87098 73947 87406 73956
rect 84326 73912 84382 73921
rect 84326 73847 84382 73856
rect 88572 73785 88600 74294
rect 88558 73776 88614 73785
rect 88558 73711 88614 73720
rect 87834 73468 88142 73477
rect 87834 73466 87840 73468
rect 87896 73466 87920 73468
rect 87976 73466 88000 73468
rect 88056 73466 88080 73468
rect 88136 73466 88142 73468
rect 87896 73414 87898 73466
rect 88078 73414 88080 73466
rect 87834 73412 87840 73414
rect 87896 73412 87920 73414
rect 87976 73412 88000 73414
rect 88056 73412 88080 73414
rect 88136 73412 88142 73414
rect 87834 73403 88142 73412
rect 88652 73230 88704 73236
rect 88652 73172 88704 73178
rect 88664 73105 88692 73172
rect 88650 73096 88706 73105
rect 84328 73060 84380 73066
rect 88650 73031 88706 73040
rect 84328 73002 84380 73008
rect 84340 72833 84368 73002
rect 87098 72924 87406 72933
rect 87098 72922 87104 72924
rect 87160 72922 87184 72924
rect 87240 72922 87264 72924
rect 87320 72922 87344 72924
rect 87400 72922 87406 72924
rect 87160 72870 87162 72922
rect 87342 72870 87344 72922
rect 87098 72868 87104 72870
rect 87160 72868 87184 72870
rect 87240 72868 87264 72870
rect 87320 72868 87344 72870
rect 87400 72868 87406 72870
rect 87098 72859 87406 72868
rect 84326 72824 84382 72833
rect 84326 72759 84382 72768
rect 87834 72380 88142 72389
rect 87834 72378 87840 72380
rect 87896 72378 87920 72380
rect 87976 72378 88000 72380
rect 88056 72378 88080 72380
rect 88136 72378 88142 72380
rect 87896 72326 87898 72378
rect 88078 72326 88080 72378
rect 87834 72324 87840 72326
rect 87896 72324 87920 72326
rect 87976 72324 88000 72326
rect 88056 72324 88080 72326
rect 88136 72324 88142 72326
rect 87834 72315 88142 72324
rect 90124 72108 90176 72114
rect 90124 72050 90176 72056
rect 87180 72040 87232 72046
rect 87178 72008 87180 72017
rect 87232 72008 87234 72017
rect 87178 71943 87234 71952
rect 87098 71836 87406 71845
rect 87098 71834 87104 71836
rect 87160 71834 87184 71836
rect 87240 71834 87264 71836
rect 87320 71834 87344 71836
rect 87400 71834 87406 71836
rect 87160 71782 87162 71834
rect 87342 71782 87344 71834
rect 87098 71780 87104 71782
rect 87160 71780 87184 71782
rect 87240 71780 87264 71782
rect 87320 71780 87344 71782
rect 87400 71780 87406 71782
rect 87098 71771 87406 71780
rect 90136 71745 90164 72050
rect 90122 71736 90178 71745
rect 90122 71671 90178 71680
rect 87834 71292 88142 71301
rect 87834 71290 87840 71292
rect 87896 71290 87920 71292
rect 87976 71290 88000 71292
rect 88056 71290 88080 71292
rect 88136 71290 88142 71292
rect 87896 71238 87898 71290
rect 88078 71238 88080 71290
rect 87834 71236 87840 71238
rect 87896 71236 87920 71238
rect 87976 71236 88000 71238
rect 88056 71236 88080 71238
rect 88136 71236 88142 71238
rect 87834 71227 88142 71236
rect 87098 70748 87406 70757
rect 87098 70746 87104 70748
rect 87160 70746 87184 70748
rect 87240 70746 87264 70748
rect 87320 70746 87344 70748
rect 87400 70746 87406 70748
rect 87160 70694 87162 70746
rect 87342 70694 87344 70746
rect 87098 70692 87104 70694
rect 87160 70692 87184 70694
rect 87240 70692 87264 70694
rect 87320 70692 87344 70694
rect 87400 70692 87406 70694
rect 87098 70683 87406 70692
rect 84326 70648 84382 70657
rect 84326 70583 84382 70592
rect 84340 70550 84368 70583
rect 84328 70544 84380 70550
rect 84328 70486 84380 70492
rect 89940 70408 89992 70414
rect 89938 70376 89940 70385
rect 89992 70376 89994 70385
rect 89938 70311 89994 70320
rect 87834 70204 88142 70213
rect 87834 70202 87840 70204
rect 87896 70202 87920 70204
rect 87976 70202 88000 70204
rect 88056 70202 88080 70204
rect 88136 70202 88142 70204
rect 87896 70150 87898 70202
rect 88078 70150 88080 70202
rect 87834 70148 87840 70150
rect 87896 70148 87920 70150
rect 87976 70148 88000 70150
rect 88056 70148 88080 70150
rect 88136 70148 88142 70150
rect 87834 70139 88142 70148
rect 88560 70000 88612 70006
rect 88560 69942 88612 69948
rect 84328 69864 84380 69870
rect 84328 69806 84380 69812
rect 84340 69569 84368 69806
rect 88572 69705 88600 69942
rect 88558 69696 88614 69705
rect 87098 69660 87406 69669
rect 87098 69658 87104 69660
rect 87160 69658 87184 69660
rect 87240 69658 87264 69660
rect 87320 69658 87344 69660
rect 87400 69658 87406 69660
rect 87160 69606 87162 69658
rect 87342 69606 87344 69658
rect 88558 69631 88614 69640
rect 87098 69604 87104 69606
rect 87160 69604 87184 69606
rect 87240 69604 87264 69606
rect 87320 69604 87344 69606
rect 87400 69604 87406 69606
rect 87098 69595 87406 69604
rect 84326 69560 84382 69569
rect 84326 69495 84382 69504
rect 89940 69320 89992 69326
rect 89940 69262 89992 69268
rect 87834 69116 88142 69125
rect 87834 69114 87840 69116
rect 87896 69114 87920 69116
rect 87976 69114 88000 69116
rect 88056 69114 88080 69116
rect 88136 69114 88142 69116
rect 87896 69062 87898 69114
rect 88078 69062 88080 69114
rect 87834 69060 87840 69062
rect 87896 69060 87920 69062
rect 87976 69060 88000 69062
rect 88056 69060 88080 69062
rect 88136 69060 88142 69062
rect 87834 69051 88142 69060
rect 89952 69025 89980 69262
rect 89938 69016 89994 69025
rect 89938 68951 89994 68960
rect 88652 68878 88704 68884
rect 88652 68820 88704 68826
rect 84328 68708 84380 68714
rect 84328 68650 84380 68656
rect 84340 68481 84368 68650
rect 87098 68572 87406 68581
rect 87098 68570 87104 68572
rect 87160 68570 87184 68572
rect 87240 68570 87264 68572
rect 87320 68570 87344 68572
rect 87400 68570 87406 68572
rect 87160 68518 87162 68570
rect 87342 68518 87344 68570
rect 87098 68516 87104 68518
rect 87160 68516 87184 68518
rect 87240 68516 87264 68518
rect 87320 68516 87344 68518
rect 87400 68516 87406 68518
rect 87098 68507 87406 68516
rect 84326 68472 84382 68481
rect 84326 68407 84382 68416
rect 88664 68345 88692 68820
rect 88650 68336 88706 68345
rect 88650 68271 88706 68280
rect 87834 68028 88142 68037
rect 87834 68026 87840 68028
rect 87896 68026 87920 68028
rect 87976 68026 88000 68028
rect 88056 68026 88080 68028
rect 88136 68026 88142 68028
rect 87896 67974 87898 68026
rect 88078 67974 88080 68026
rect 87834 67972 87840 67974
rect 87896 67972 87920 67974
rect 87976 67972 88000 67974
rect 88056 67972 88080 67974
rect 88136 67972 88142 67974
rect 87834 67963 88142 67972
rect 88652 67790 88704 67796
rect 88652 67732 88704 67738
rect 88664 67665 88692 67732
rect 88650 67656 88706 67665
rect 84328 67620 84380 67626
rect 88650 67591 88706 67600
rect 84328 67562 84380 67568
rect 84340 67393 84368 67562
rect 87098 67484 87406 67493
rect 87098 67482 87104 67484
rect 87160 67482 87184 67484
rect 87240 67482 87264 67484
rect 87320 67482 87344 67484
rect 87400 67482 87406 67484
rect 87160 67430 87162 67482
rect 87342 67430 87344 67482
rect 87098 67428 87104 67430
rect 87160 67428 87184 67430
rect 87240 67428 87264 67430
rect 87320 67428 87344 67430
rect 87400 67428 87406 67430
rect 87098 67419 87406 67428
rect 84326 67384 84382 67393
rect 84326 67319 84382 67328
rect 87834 66940 88142 66949
rect 87834 66938 87840 66940
rect 87896 66938 87920 66940
rect 87976 66938 88000 66940
rect 88056 66938 88080 66940
rect 88136 66938 88142 66940
rect 87896 66886 87898 66938
rect 88078 66886 88080 66938
rect 87834 66884 87840 66886
rect 87896 66884 87920 66886
rect 87976 66884 88000 66886
rect 88056 66884 88080 66886
rect 88136 66884 88142 66886
rect 87834 66875 88142 66884
rect 90124 66668 90176 66674
rect 90124 66610 90176 66616
rect 87456 66532 87508 66538
rect 87456 66474 87508 66480
rect 87098 66396 87406 66405
rect 87098 66394 87104 66396
rect 87160 66394 87184 66396
rect 87240 66394 87264 66396
rect 87320 66394 87344 66396
rect 87400 66394 87406 66396
rect 87160 66342 87162 66394
rect 87342 66342 87344 66394
rect 87098 66340 87104 66342
rect 87160 66340 87184 66342
rect 87240 66340 87264 66342
rect 87320 66340 87344 66342
rect 87400 66340 87406 66342
rect 87098 66331 87406 66340
rect 87468 66169 87496 66474
rect 90136 66305 90164 66610
rect 90122 66296 90178 66305
rect 90122 66231 90178 66240
rect 87454 66160 87510 66169
rect 87454 66095 87510 66104
rect 87834 65852 88142 65861
rect 87834 65850 87840 65852
rect 87896 65850 87920 65852
rect 87976 65850 88000 65852
rect 88056 65850 88080 65852
rect 88136 65850 88142 65852
rect 87896 65798 87898 65850
rect 88078 65798 88080 65850
rect 87834 65796 87840 65798
rect 87896 65796 87920 65798
rect 87976 65796 88000 65798
rect 88056 65796 88080 65798
rect 88136 65796 88142 65798
rect 87834 65787 88142 65796
rect 87098 65308 87406 65317
rect 87098 65306 87104 65308
rect 87160 65306 87184 65308
rect 87240 65306 87264 65308
rect 87320 65306 87344 65308
rect 87400 65306 87406 65308
rect 87160 65254 87162 65306
rect 87342 65254 87344 65306
rect 87098 65252 87104 65254
rect 87160 65252 87184 65254
rect 87240 65252 87264 65254
rect 87320 65252 87344 65254
rect 87400 65252 87406 65254
rect 87098 65243 87406 65252
rect 84326 65140 84382 65149
rect 84326 65075 84382 65084
rect 84340 65042 84368 65075
rect 84328 65036 84380 65042
rect 84328 64978 84380 64984
rect 89938 64936 89994 64945
rect 89938 64871 89940 64880
rect 89992 64871 89994 64880
rect 89940 64842 89992 64848
rect 87834 64764 88142 64773
rect 87834 64762 87840 64764
rect 87896 64762 87920 64764
rect 87976 64762 88000 64764
rect 88056 64762 88080 64764
rect 88136 64762 88142 64764
rect 87896 64710 87898 64762
rect 88078 64710 88080 64762
rect 87834 64708 87840 64710
rect 87896 64708 87920 64710
rect 87976 64708 88000 64710
rect 88056 64708 88080 64710
rect 88136 64708 88142 64710
rect 87834 64699 88142 64708
rect 84328 64492 84380 64498
rect 84328 64434 84380 64440
rect 84340 64129 84368 64434
rect 88560 64356 88612 64362
rect 88560 64298 88612 64304
rect 88572 64265 88600 64298
rect 88558 64256 88614 64265
rect 87098 64220 87406 64229
rect 87098 64218 87104 64220
rect 87160 64218 87184 64220
rect 87240 64218 87264 64220
rect 87320 64218 87344 64220
rect 87400 64218 87406 64220
rect 87160 64166 87162 64218
rect 87342 64166 87344 64218
rect 88558 64191 88614 64200
rect 87098 64164 87104 64166
rect 87160 64164 87184 64166
rect 87240 64164 87264 64166
rect 87320 64164 87344 64166
rect 87400 64164 87406 64166
rect 87098 64155 87406 64164
rect 84326 64120 84382 64129
rect 84326 64055 84382 64064
rect 87834 63676 88142 63685
rect 87834 63674 87840 63676
rect 87896 63674 87920 63676
rect 87976 63674 88000 63676
rect 88056 63674 88080 63676
rect 88136 63674 88142 63676
rect 87896 63622 87898 63674
rect 88078 63622 88080 63674
rect 87834 63620 87840 63622
rect 87896 63620 87920 63622
rect 87976 63620 88000 63622
rect 88056 63620 88080 63622
rect 88136 63620 88142 63622
rect 87834 63611 88142 63620
rect 84328 63404 84380 63410
rect 84328 63346 84380 63352
rect 84340 63041 84368 63346
rect 88560 63268 88612 63274
rect 88560 63210 88612 63216
rect 87098 63132 87406 63141
rect 87098 63130 87104 63132
rect 87160 63130 87184 63132
rect 87240 63130 87264 63132
rect 87320 63130 87344 63132
rect 87400 63130 87406 63132
rect 87160 63078 87162 63130
rect 87342 63078 87344 63130
rect 87098 63076 87104 63078
rect 87160 63076 87184 63078
rect 87240 63076 87264 63078
rect 87320 63076 87344 63078
rect 87400 63076 87406 63078
rect 87098 63067 87406 63076
rect 84326 63032 84382 63041
rect 84326 62967 84382 62976
rect 88572 62905 88600 63210
rect 88558 62896 88614 62905
rect 88558 62831 88614 62840
rect 87834 62588 88142 62597
rect 87834 62586 87840 62588
rect 87896 62586 87920 62588
rect 87976 62586 88000 62588
rect 88056 62586 88080 62588
rect 88136 62586 88142 62588
rect 87896 62534 87898 62586
rect 88078 62534 88080 62586
rect 87834 62532 87840 62534
rect 87896 62532 87920 62534
rect 87976 62532 88000 62534
rect 88056 62532 88080 62534
rect 88136 62532 88142 62534
rect 87834 62523 88142 62532
rect 89940 62384 89992 62390
rect 88376 62350 88428 62356
rect 89940 62326 89992 62332
rect 88376 62292 88428 62298
rect 88388 62225 88416 62292
rect 89952 62225 89980 62326
rect 88374 62216 88430 62225
rect 88374 62151 88430 62160
rect 89938 62216 89994 62225
rect 89938 62151 89994 62160
rect 87098 62044 87406 62053
rect 87098 62042 87104 62044
rect 87160 62042 87184 62044
rect 87240 62042 87264 62044
rect 87320 62042 87344 62044
rect 87400 62042 87406 62044
rect 87160 61990 87162 62042
rect 87342 61990 87344 62042
rect 87098 61988 87104 61990
rect 87160 61988 87184 61990
rect 87240 61988 87264 61990
rect 87320 61988 87344 61990
rect 87400 61988 87406 61990
rect 87098 61979 87406 61988
rect 87834 61500 88142 61509
rect 87834 61498 87840 61500
rect 87896 61498 87920 61500
rect 87976 61498 88000 61500
rect 88056 61498 88080 61500
rect 88136 61498 88142 61500
rect 87896 61446 87898 61498
rect 88078 61446 88080 61498
rect 87834 61444 87840 61446
rect 87896 61444 87920 61446
rect 87976 61444 88000 61446
rect 88056 61444 88080 61446
rect 88136 61444 88142 61446
rect 87834 61435 88142 61444
rect 88376 61262 88428 61268
rect 88376 61204 88428 61210
rect 87098 60956 87406 60965
rect 87098 60954 87104 60956
rect 87160 60954 87184 60956
rect 87240 60954 87264 60956
rect 87320 60954 87344 60956
rect 87400 60954 87406 60956
rect 87160 60902 87162 60954
rect 87342 60902 87344 60954
rect 87098 60900 87104 60902
rect 87160 60900 87184 60902
rect 87240 60900 87264 60902
rect 87320 60900 87344 60902
rect 87400 60900 87406 60902
rect 87098 60891 87406 60900
rect 88388 60729 88416 61204
rect 89940 61092 89992 61098
rect 89940 61034 89992 61040
rect 89952 60865 89980 61034
rect 89938 60856 89994 60865
rect 89938 60791 89994 60800
rect 88374 60720 88430 60729
rect 88374 60655 88430 60664
rect 87834 60412 88142 60421
rect 87834 60410 87840 60412
rect 87896 60410 87920 60412
rect 87976 60410 88000 60412
rect 88056 60410 88080 60412
rect 88136 60410 88142 60412
rect 87896 60358 87898 60410
rect 88078 60358 88080 60410
rect 87834 60356 87840 60358
rect 87896 60356 87920 60358
rect 87976 60356 88000 60358
rect 88056 60356 88080 60358
rect 88136 60356 88142 60358
rect 87834 60347 88142 60356
rect 87098 59868 87406 59877
rect 87098 59866 87104 59868
rect 87160 59866 87184 59868
rect 87240 59866 87264 59868
rect 87320 59866 87344 59868
rect 87400 59866 87406 59868
rect 87160 59814 87162 59866
rect 87342 59814 87344 59866
rect 87098 59812 87104 59814
rect 87160 59812 87184 59814
rect 87240 59812 87264 59814
rect 87320 59812 87344 59814
rect 87400 59812 87406 59814
rect 87098 59803 87406 59812
rect 84326 59700 84382 59709
rect 84326 59635 84382 59644
rect 84340 59534 84368 59635
rect 84328 59528 84380 59534
rect 84328 59470 84380 59476
rect 89938 59496 89994 59505
rect 89938 59431 89940 59440
rect 89992 59431 89994 59440
rect 89940 59402 89992 59408
rect 87834 59324 88142 59333
rect 87834 59322 87840 59324
rect 87896 59322 87920 59324
rect 87976 59322 88000 59324
rect 88056 59322 88080 59324
rect 88136 59322 88142 59324
rect 87896 59270 87898 59322
rect 88078 59270 88080 59322
rect 87834 59268 87840 59270
rect 87896 59268 87920 59270
rect 87976 59268 88000 59270
rect 88056 59268 88080 59270
rect 88136 59268 88142 59270
rect 87834 59259 88142 59268
rect 84328 59052 84380 59058
rect 84328 58994 84380 59000
rect 84340 58689 84368 58994
rect 88560 58916 88612 58922
rect 88560 58858 88612 58864
rect 88572 58825 88600 58858
rect 88558 58816 88614 58825
rect 87098 58780 87406 58789
rect 87098 58778 87104 58780
rect 87160 58778 87184 58780
rect 87240 58778 87264 58780
rect 87320 58778 87344 58780
rect 87400 58778 87406 58780
rect 87160 58726 87162 58778
rect 87342 58726 87344 58778
rect 88558 58751 88614 58760
rect 87098 58724 87104 58726
rect 87160 58724 87184 58726
rect 87240 58724 87264 58726
rect 87320 58724 87344 58726
rect 87400 58724 87406 58726
rect 87098 58715 87406 58724
rect 84326 58680 84382 58689
rect 84326 58615 84382 58624
rect 87834 58236 88142 58245
rect 87834 58234 87840 58236
rect 87896 58234 87920 58236
rect 87976 58234 88000 58236
rect 88056 58234 88080 58236
rect 88136 58234 88142 58236
rect 87896 58182 87898 58234
rect 88078 58182 88080 58234
rect 87834 58180 87840 58182
rect 87896 58180 87920 58182
rect 87976 58180 88000 58182
rect 88056 58180 88080 58182
rect 88136 58180 88142 58182
rect 87834 58171 88142 58180
rect 84328 57964 84380 57970
rect 84328 57906 84380 57912
rect 84340 57601 84368 57906
rect 88560 57828 88612 57834
rect 88560 57770 88612 57776
rect 87098 57692 87406 57701
rect 87098 57690 87104 57692
rect 87160 57690 87184 57692
rect 87240 57690 87264 57692
rect 87320 57690 87344 57692
rect 87400 57690 87406 57692
rect 87160 57638 87162 57690
rect 87342 57638 87344 57690
rect 87098 57636 87104 57638
rect 87160 57636 87184 57638
rect 87240 57636 87264 57638
rect 87320 57636 87344 57638
rect 87400 57636 87406 57638
rect 87098 57627 87406 57636
rect 84326 57592 84382 57601
rect 84326 57527 84382 57536
rect 88572 57465 88600 57770
rect 88558 57456 88614 57465
rect 88558 57391 88614 57400
rect 87834 57148 88142 57157
rect 87834 57146 87840 57148
rect 87896 57146 87920 57148
rect 87976 57146 88000 57148
rect 88056 57146 88080 57148
rect 88136 57146 88142 57148
rect 87896 57094 87898 57146
rect 88078 57094 88080 57146
rect 87834 57092 87840 57094
rect 87896 57092 87920 57094
rect 87976 57092 88000 57094
rect 88056 57092 88080 57094
rect 88136 57092 88142 57094
rect 87834 57083 88142 57092
rect 88284 56910 88336 56916
rect 88284 56852 88336 56858
rect 89940 56876 89992 56882
rect 88296 56785 88324 56852
rect 89940 56818 89992 56824
rect 89952 56785 89980 56818
rect 88282 56776 88338 56785
rect 88282 56711 88338 56720
rect 89938 56776 89994 56785
rect 89938 56711 89994 56720
rect 87098 56604 87406 56613
rect 87098 56602 87104 56604
rect 87160 56602 87184 56604
rect 87240 56602 87264 56604
rect 87320 56602 87344 56604
rect 87400 56602 87406 56604
rect 87160 56550 87162 56602
rect 87342 56550 87344 56602
rect 87098 56548 87104 56550
rect 87160 56548 87184 56550
rect 87240 56548 87264 56550
rect 87320 56548 87344 56550
rect 87400 56548 87406 56550
rect 87098 56539 87406 56548
rect 87834 56060 88142 56069
rect 87834 56058 87840 56060
rect 87896 56058 87920 56060
rect 87976 56058 88000 56060
rect 88056 56058 88080 56060
rect 88136 56058 88142 56060
rect 87896 56006 87898 56058
rect 88078 56006 88080 56058
rect 87834 56004 87840 56006
rect 87896 56004 87920 56006
rect 87976 56004 88000 56006
rect 88056 56004 88080 56006
rect 88136 56004 88142 56006
rect 87834 55995 88142 56004
rect 88376 55822 88428 55828
rect 88376 55764 88428 55770
rect 87098 55516 87406 55525
rect 87098 55514 87104 55516
rect 87160 55514 87184 55516
rect 87240 55514 87264 55516
rect 87320 55514 87344 55516
rect 87400 55514 87406 55516
rect 87160 55462 87162 55514
rect 87342 55462 87344 55514
rect 87098 55460 87104 55462
rect 87160 55460 87184 55462
rect 87240 55460 87264 55462
rect 87320 55460 87344 55462
rect 87400 55460 87406 55462
rect 87098 55451 87406 55460
rect 88388 55289 88416 55764
rect 89940 55652 89992 55658
rect 89940 55594 89992 55600
rect 89952 55425 89980 55594
rect 89938 55416 89994 55425
rect 89938 55351 89994 55360
rect 88374 55280 88430 55289
rect 88374 55215 88430 55224
rect 87834 54972 88142 54981
rect 87834 54970 87840 54972
rect 87896 54970 87920 54972
rect 87976 54970 88000 54972
rect 88056 54970 88080 54972
rect 88136 54970 88142 54972
rect 87896 54918 87898 54970
rect 88078 54918 88080 54970
rect 87834 54916 87840 54918
rect 87896 54916 87920 54918
rect 87976 54916 88000 54918
rect 88056 54916 88080 54918
rect 88136 54916 88142 54918
rect 87834 54907 88142 54916
rect 87098 54428 87406 54437
rect 87098 54426 87104 54428
rect 87160 54426 87184 54428
rect 87240 54426 87264 54428
rect 87320 54426 87344 54428
rect 87400 54426 87406 54428
rect 87160 54374 87162 54426
rect 87342 54374 87344 54426
rect 87098 54372 87104 54374
rect 87160 54372 87184 54374
rect 87240 54372 87264 54374
rect 87320 54372 87344 54374
rect 87400 54372 87406 54374
rect 87098 54363 87406 54372
rect 84326 54260 84382 54269
rect 84326 54195 84382 54204
rect 84340 54162 84368 54195
rect 84328 54156 84380 54162
rect 84328 54098 84380 54104
rect 89940 54088 89992 54094
rect 89938 54056 89940 54065
rect 89992 54056 89994 54065
rect 89938 53991 89994 54000
rect 87834 53884 88142 53893
rect 87834 53882 87840 53884
rect 87896 53882 87920 53884
rect 87976 53882 88000 53884
rect 88056 53882 88080 53884
rect 88136 53882 88142 53884
rect 87896 53830 87898 53882
rect 88078 53830 88080 53882
rect 87834 53828 87840 53830
rect 87896 53828 87920 53830
rect 87976 53828 88000 53830
rect 88056 53828 88080 53830
rect 88136 53828 88142 53830
rect 87834 53819 88142 53828
rect 84328 53612 84380 53618
rect 84328 53554 84380 53560
rect 84340 53249 84368 53554
rect 88560 53476 88612 53482
rect 88560 53418 88612 53424
rect 88572 53385 88600 53418
rect 88558 53376 88614 53385
rect 87098 53340 87406 53349
rect 87098 53338 87104 53340
rect 87160 53338 87184 53340
rect 87240 53338 87264 53340
rect 87320 53338 87344 53340
rect 87400 53338 87406 53340
rect 87160 53286 87162 53338
rect 87342 53286 87344 53338
rect 88558 53311 88614 53320
rect 87098 53284 87104 53286
rect 87160 53284 87184 53286
rect 87240 53284 87264 53286
rect 87320 53284 87344 53286
rect 87400 53284 87406 53286
rect 87098 53275 87406 53284
rect 84326 53240 84382 53249
rect 84326 53175 84382 53184
rect 89940 53000 89992 53006
rect 89940 52942 89992 52948
rect 87834 52796 88142 52805
rect 87834 52794 87840 52796
rect 87896 52794 87920 52796
rect 87976 52794 88000 52796
rect 88056 52794 88080 52796
rect 88136 52794 88142 52796
rect 87896 52742 87898 52794
rect 88078 52742 88080 52794
rect 87834 52740 87840 52742
rect 87896 52740 87920 52742
rect 87976 52740 88000 52742
rect 88056 52740 88080 52742
rect 88136 52740 88142 52742
rect 87834 52731 88142 52740
rect 89952 52705 89980 52942
rect 89938 52696 89994 52705
rect 89938 52631 89994 52640
rect 84328 52524 84380 52530
rect 84328 52466 84380 52472
rect 84340 52161 84368 52466
rect 88560 52388 88612 52394
rect 88560 52330 88612 52336
rect 87098 52252 87406 52261
rect 87098 52250 87104 52252
rect 87160 52250 87184 52252
rect 87240 52250 87264 52252
rect 87320 52250 87344 52252
rect 87400 52250 87406 52252
rect 87160 52198 87162 52250
rect 87342 52198 87344 52250
rect 87098 52196 87104 52198
rect 87160 52196 87184 52198
rect 87240 52196 87264 52198
rect 87320 52196 87344 52198
rect 87400 52196 87406 52198
rect 87098 52187 87406 52196
rect 84326 52152 84382 52161
rect 84326 52087 84382 52096
rect 88572 52025 88600 52330
rect 88558 52016 88614 52025
rect 88558 51951 88614 51960
rect 87834 51708 88142 51717
rect 87834 51706 87840 51708
rect 87896 51706 87920 51708
rect 87976 51706 88000 51708
rect 88056 51706 88080 51708
rect 88136 51706 88142 51708
rect 87896 51654 87898 51706
rect 88078 51654 88080 51706
rect 87834 51652 87840 51654
rect 87896 51652 87920 51654
rect 87976 51652 88000 51654
rect 88056 51652 88080 51654
rect 88136 51652 88142 51654
rect 87834 51643 88142 51652
rect 88376 51470 88428 51476
rect 88376 51412 88428 51418
rect 87098 51164 87406 51173
rect 87098 51162 87104 51164
rect 87160 51162 87184 51164
rect 87240 51162 87264 51164
rect 87320 51162 87344 51164
rect 87400 51162 87406 51164
rect 87160 51110 87162 51162
rect 87342 51110 87344 51162
rect 87098 51108 87104 51110
rect 87160 51108 87184 51110
rect 87240 51108 87264 51110
rect 87320 51108 87344 51110
rect 87400 51108 87406 51110
rect 87098 51099 87406 51108
rect 88388 50937 88416 51412
rect 88560 51368 88612 51374
rect 88558 51336 88560 51345
rect 88612 51336 88614 51345
rect 88558 51271 88614 51280
rect 88374 50928 88430 50937
rect 88374 50863 88430 50872
rect 87834 50620 88142 50629
rect 87834 50618 87840 50620
rect 87896 50618 87920 50620
rect 87976 50618 88000 50620
rect 88056 50618 88080 50620
rect 88136 50618 88142 50620
rect 87896 50566 87898 50618
rect 88078 50566 88080 50618
rect 87834 50564 87840 50566
rect 87896 50564 87920 50566
rect 87976 50564 88000 50566
rect 88056 50564 88080 50566
rect 88136 50564 88142 50566
rect 87834 50555 88142 50564
rect 87098 50076 87406 50085
rect 87098 50074 87104 50076
rect 87160 50074 87184 50076
rect 87240 50074 87264 50076
rect 87320 50074 87344 50076
rect 87400 50074 87406 50076
rect 87160 50022 87162 50074
rect 87342 50022 87344 50074
rect 87098 50020 87104 50022
rect 87160 50020 87184 50022
rect 87240 50020 87264 50022
rect 87320 50020 87344 50022
rect 87400 50020 87406 50022
rect 87098 50011 87406 50020
rect 89940 49736 89992 49742
rect 89940 49678 89992 49684
rect 87834 49532 88142 49541
rect 87834 49530 87840 49532
rect 87896 49530 87920 49532
rect 87976 49530 88000 49532
rect 88056 49530 88080 49532
rect 88136 49530 88142 49532
rect 87896 49478 87898 49530
rect 88078 49478 88080 49530
rect 87834 49476 87840 49478
rect 87896 49476 87920 49478
rect 87976 49476 88000 49478
rect 88056 49476 88080 49478
rect 88136 49476 88142 49478
rect 87834 49467 88142 49476
rect 89952 49305 89980 49678
rect 89938 49296 89994 49305
rect 89938 49231 89994 49240
rect 87098 48988 87406 48997
rect 87098 48986 87104 48988
rect 87160 48986 87184 48988
rect 87240 48986 87264 48988
rect 87320 48986 87344 48988
rect 87400 48986 87406 48988
rect 87160 48934 87162 48986
rect 87342 48934 87344 48986
rect 87098 48932 87104 48934
rect 87160 48932 87184 48934
rect 87240 48932 87264 48934
rect 87320 48932 87344 48934
rect 87400 48932 87406 48934
rect 87098 48923 87406 48932
rect 89940 48648 89992 48654
rect 89938 48616 89940 48625
rect 89992 48616 89994 48625
rect 89938 48551 89994 48560
rect 87834 48444 88142 48453
rect 87834 48442 87840 48444
rect 87896 48442 87920 48444
rect 87976 48442 88000 48444
rect 88056 48442 88080 48444
rect 88136 48442 88142 48444
rect 87896 48390 87898 48442
rect 88078 48390 88080 48442
rect 87834 48388 87840 48390
rect 87896 48388 87920 48390
rect 87976 48388 88000 48390
rect 88056 48388 88080 48390
rect 88136 48388 88142 48390
rect 87834 48379 88142 48388
rect 88560 48036 88612 48042
rect 88560 47978 88612 47984
rect 88572 47945 88600 47978
rect 88558 47936 88614 47945
rect 87098 47900 87406 47909
rect 87098 47898 87104 47900
rect 87160 47898 87184 47900
rect 87240 47898 87264 47900
rect 87320 47898 87344 47900
rect 87400 47898 87406 47900
rect 87160 47846 87162 47898
rect 87342 47846 87344 47898
rect 88558 47871 88614 47880
rect 87098 47844 87104 47846
rect 87160 47844 87184 47846
rect 87240 47844 87264 47846
rect 87320 47844 87344 47846
rect 87400 47844 87406 47846
rect 87098 47835 87406 47844
rect 84420 47356 84472 47362
rect 84420 47298 84472 47304
rect 87834 47356 88142 47365
rect 87834 47354 87840 47356
rect 87896 47354 87920 47356
rect 87976 47354 88000 47356
rect 88056 47354 88080 47356
rect 88136 47354 88142 47356
rect 87896 47302 87898 47354
rect 88078 47302 88080 47354
rect 87834 47300 87840 47302
rect 87896 47300 87920 47302
rect 87976 47300 88000 47302
rect 88056 47300 88080 47302
rect 88136 47300 88142 47302
rect 84052 46812 84104 46818
rect 84052 46754 84104 46760
rect 49552 46744 49604 46750
rect 47856 46692 48152 46698
rect 47804 46686 48152 46692
rect 11016 46670 11122 46686
rect 47816 46670 48152 46686
rect 49104 46692 49552 46698
rect 49104 46686 49604 46692
rect 83684 46744 83736 46750
rect 83684 46686 83736 46692
rect 49104 46670 49592 46686
rect 84328 43140 84380 43146
rect 84328 43082 84380 43088
rect 84340 43049 84368 43082
rect 84326 43040 84382 43049
rect 84326 42975 84382 42984
rect 84328 42052 84380 42058
rect 84328 41994 84380 42000
rect 84340 41961 84368 41994
rect 84326 41952 84382 41961
rect 84326 41887 84382 41896
rect 84328 39944 84380 39950
rect 84328 39886 84380 39892
rect 84340 39785 84368 39886
rect 84326 39776 84382 39785
rect 84326 39711 84382 39720
rect 84328 37768 84380 37774
rect 84328 37710 84380 37716
rect 84340 37609 84368 37710
rect 84326 37600 84382 37609
rect 84326 37535 84382 37544
rect 84328 36680 84380 36686
rect 84328 36622 84380 36628
rect 84340 36521 84368 36622
rect 84326 36512 84382 36521
rect 84326 36447 84382 36456
rect 84328 34436 84380 34442
rect 84328 34378 84380 34384
rect 84340 34345 84368 34378
rect 84326 34336 84382 34345
rect 84326 34271 84382 34280
rect 84328 32328 84380 32334
rect 84328 32270 84380 32276
rect 84340 32169 84368 32270
rect 84326 32160 84382 32169
rect 84326 32095 84382 32104
rect 84328 31172 84380 31178
rect 84328 31114 84380 31120
rect 84340 31081 84368 31114
rect 84326 31072 84382 31081
rect 84326 31007 84382 31016
rect 84328 28996 84380 29002
rect 84328 28938 84380 28944
rect 84340 28905 84368 28938
rect 84326 28896 84382 28905
rect 84326 28831 84382 28840
rect 84328 26888 84380 26894
rect 84328 26830 84380 26836
rect 84340 26729 84368 26830
rect 84326 26720 84382 26729
rect 84326 26655 84382 26664
rect 84328 25800 84380 25806
rect 84328 25742 84380 25748
rect 84340 25641 84368 25742
rect 84326 25632 84382 25641
rect 84326 25567 84382 25576
rect 84328 23624 84380 23630
rect 84328 23566 84380 23572
rect 84340 23465 84368 23566
rect 84326 23456 84382 23465
rect 84326 23391 84382 23400
rect 84328 22536 84380 22542
rect 84328 22478 84380 22484
rect 84340 22377 84368 22478
rect 84326 22368 84382 22377
rect 84326 22303 84382 22312
rect 84328 21448 84380 21454
rect 84328 21390 84380 21396
rect 84340 21289 84368 21390
rect 84326 21280 84382 21289
rect 84326 21215 84382 21224
rect 84328 20360 84380 20366
rect 84328 20302 84380 20308
rect 84340 20201 84368 20302
rect 84326 20192 84382 20201
rect 84326 20127 84382 20136
rect 84328 17096 84380 17102
rect 84328 17038 84380 17044
rect 84340 16937 84368 17038
rect 84326 16928 84382 16937
rect 84326 16863 84382 16872
rect 84328 16008 84380 16014
rect 84328 15950 84380 15956
rect 84340 15849 84368 15950
rect 84326 15840 84382 15849
rect 84326 15775 84382 15784
rect 84328 14920 84380 14926
rect 84328 14862 84380 14868
rect 84340 14761 84368 14862
rect 84326 14752 84382 14761
rect 84326 14687 84382 14696
rect 9806 10672 9862 10681
rect 9806 10607 9862 10616
rect 11122 10672 11178 10681
rect 11122 10607 11178 10616
rect 12226 10536 12282 10545
rect 12226 10471 12282 10480
rect 12240 10137 12268 10471
rect 13330 10400 13386 10409
rect 13330 10335 13386 10344
rect 46698 10400 46754 10409
rect 46698 10335 46754 10344
rect 13344 10137 13372 10335
rect 14434 10264 14490 10273
rect 14434 10199 14490 10208
rect 12226 10128 12282 10137
rect 12226 10063 12282 10072
rect 13330 10128 13386 10137
rect 13330 10063 13386 10072
rect 12658 9992 12714 10001
rect 12658 9927 12714 9936
rect 14682 9992 14738 10001
rect 14682 9927 14738 9936
rect 15418 9992 15474 10001
rect 15418 9927 15474 9936
rect 8426 8496 8482 8505
rect 8426 8431 8482 8440
rect 6690 8188 6998 8197
rect 6690 8186 6696 8188
rect 6752 8186 6776 8188
rect 6832 8186 6856 8188
rect 6912 8186 6936 8188
rect 6992 8186 6998 8188
rect 6752 8134 6754 8186
rect 6934 8134 6936 8186
rect 6690 8132 6696 8134
rect 6752 8132 6776 8134
rect 6832 8132 6856 8134
rect 6912 8132 6936 8134
rect 6992 8132 6998 8134
rect 6690 8123 6998 8132
rect 5954 7644 6262 7653
rect 5954 7642 5960 7644
rect 6016 7642 6040 7644
rect 6096 7642 6120 7644
rect 6176 7642 6200 7644
rect 6256 7642 6262 7644
rect 6016 7590 6018 7642
rect 6198 7590 6200 7642
rect 5954 7588 5960 7590
rect 6016 7588 6040 7590
rect 6096 7588 6120 7590
rect 6176 7588 6200 7590
rect 6256 7588 6262 7590
rect 5954 7579 6262 7588
rect 6690 7100 6998 7109
rect 6690 7098 6696 7100
rect 6752 7098 6776 7100
rect 6832 7098 6856 7100
rect 6912 7098 6936 7100
rect 6992 7098 6998 7100
rect 6752 7046 6754 7098
rect 6934 7046 6936 7098
rect 6690 7044 6696 7046
rect 6752 7044 6776 7046
rect 6832 7044 6856 7046
rect 6912 7044 6936 7046
rect 6992 7044 6998 7046
rect 6690 7035 6998 7044
rect 12672 5338 12700 9927
rect 14696 5338 14724 9927
rect 12660 5332 12712 5338
rect 12660 5274 12712 5280
rect 14684 5332 14736 5338
rect 14684 5274 14736 5280
rect 15432 5134 15460 9927
rect 15552 9842 15580 10100
rect 16656 9842 16684 10100
rect 17760 9842 17788 10100
rect 15524 9814 15580 9842
rect 16628 9814 16684 9842
rect 17732 9814 17788 9842
rect 18864 9842 18892 10100
rect 19968 9842 19996 10100
rect 21072 9842 21100 10100
rect 22176 9842 22204 10100
rect 18864 9814 19140 9842
rect 15524 5202 15552 9814
rect 15512 5196 15564 5202
rect 16628 5168 16656 9814
rect 17732 5168 17760 9814
rect 18722 7644 19030 7653
rect 18722 7642 18728 7644
rect 18784 7642 18808 7644
rect 18864 7642 18888 7644
rect 18944 7642 18968 7644
rect 19024 7642 19030 7644
rect 18784 7590 18786 7642
rect 18966 7590 18968 7642
rect 18722 7588 18728 7590
rect 18784 7588 18808 7590
rect 18864 7588 18888 7590
rect 18944 7588 18968 7590
rect 19024 7588 19030 7590
rect 18722 7579 19030 7588
rect 18722 6556 19030 6565
rect 18722 6554 18728 6556
rect 18784 6554 18808 6556
rect 18864 6554 18888 6556
rect 18944 6554 18968 6556
rect 19024 6554 19030 6556
rect 18784 6502 18786 6554
rect 18966 6502 18968 6554
rect 18722 6500 18728 6502
rect 18784 6500 18808 6502
rect 18864 6500 18888 6502
rect 18944 6500 18968 6502
rect 19024 6500 19030 6502
rect 18722 6491 19030 6500
rect 18722 5468 19030 5477
rect 18722 5466 18728 5468
rect 18784 5466 18808 5468
rect 18864 5466 18888 5468
rect 18944 5466 18968 5468
rect 19024 5466 19030 5468
rect 18784 5414 18786 5466
rect 18966 5414 18968 5466
rect 18722 5412 18728 5414
rect 18784 5412 18808 5414
rect 18864 5412 18888 5414
rect 18944 5412 18968 5414
rect 19024 5412 19030 5414
rect 18722 5403 19030 5412
rect 19112 5168 19140 9814
rect 19940 9814 19996 9842
rect 21044 9814 21100 9842
rect 22148 9814 22204 9842
rect 23280 9842 23308 10100
rect 24384 9842 24412 10100
rect 25488 9842 25516 10100
rect 26592 9842 26620 10100
rect 27696 9842 27724 10100
rect 28800 9842 28828 10100
rect 29904 9842 29932 10100
rect 31008 9842 31036 10100
rect 32112 9842 32140 10100
rect 33216 9842 33244 10100
rect 34320 9842 34348 10100
rect 35424 9842 35452 10100
rect 36528 9842 36556 10100
rect 37632 9842 37660 10100
rect 23280 9814 23372 9842
rect 19382 7100 19690 7109
rect 19382 7098 19388 7100
rect 19444 7098 19468 7100
rect 19524 7098 19548 7100
rect 19604 7098 19628 7100
rect 19684 7098 19690 7100
rect 19444 7046 19446 7098
rect 19626 7046 19628 7098
rect 19382 7044 19388 7046
rect 19444 7044 19468 7046
rect 19524 7044 19548 7046
rect 19604 7044 19628 7046
rect 19684 7044 19690 7046
rect 19382 7035 19690 7044
rect 19382 6012 19690 6021
rect 19382 6010 19388 6012
rect 19444 6010 19468 6012
rect 19524 6010 19548 6012
rect 19604 6010 19628 6012
rect 19684 6010 19690 6012
rect 19444 5958 19446 6010
rect 19626 5958 19628 6010
rect 19382 5956 19388 5958
rect 19444 5956 19468 5958
rect 19524 5956 19548 5958
rect 19604 5956 19628 5958
rect 19684 5956 19690 5958
rect 19382 5947 19690 5956
rect 19940 5168 19968 9814
rect 21044 5168 21072 9814
rect 22148 5168 22176 9814
rect 23344 5168 23372 9814
rect 24356 9814 24412 9842
rect 25460 9814 25516 9842
rect 26564 9814 26620 9842
rect 27668 9814 27724 9842
rect 28772 9814 28828 9842
rect 29876 9814 29932 9842
rect 30980 9814 31036 9842
rect 32084 9814 32140 9842
rect 33188 9814 33244 9842
rect 34292 9814 34348 9842
rect 35396 9814 35452 9842
rect 36500 9814 36556 9842
rect 37604 9814 37660 9842
rect 38736 9842 38764 10100
rect 39840 9842 39868 10100
rect 40944 9842 40972 10100
rect 42048 9842 42076 10100
rect 43152 9842 43180 10100
rect 44256 9842 44284 10100
rect 45360 9842 45388 10100
rect 46712 10001 46740 10335
rect 84432 10273 84460 47298
rect 87834 47291 88142 47300
rect 88560 46948 88612 46954
rect 88560 46890 88612 46896
rect 87098 46812 87406 46821
rect 87098 46810 87104 46812
rect 87160 46810 87184 46812
rect 87240 46810 87264 46812
rect 87320 46810 87344 46812
rect 87400 46810 87406 46812
rect 87160 46758 87162 46810
rect 87342 46758 87344 46810
rect 87098 46756 87104 46758
rect 87160 46756 87184 46758
rect 87240 46756 87264 46758
rect 87320 46756 87344 46758
rect 87400 46756 87406 46758
rect 87098 46747 87406 46756
rect 88572 46585 88600 46890
rect 88558 46576 88614 46585
rect 88558 46511 88614 46520
rect 87834 46268 88142 46277
rect 87834 46266 87840 46268
rect 87896 46266 87920 46268
rect 87976 46266 88000 46268
rect 88056 46266 88080 46268
rect 88136 46266 88142 46268
rect 87896 46214 87898 46266
rect 88078 46214 88080 46266
rect 87834 46212 87840 46214
rect 87896 46212 87920 46214
rect 87976 46212 88000 46214
rect 88056 46212 88080 46214
rect 88136 46212 88142 46214
rect 87834 46203 88142 46212
rect 87098 45724 87406 45733
rect 87098 45722 87104 45724
rect 87160 45722 87184 45724
rect 87240 45722 87264 45724
rect 87320 45722 87344 45724
rect 87400 45722 87406 45724
rect 87160 45670 87162 45722
rect 87342 45670 87344 45722
rect 87098 45668 87104 45670
rect 87160 45668 87184 45670
rect 87240 45668 87264 45670
rect 87320 45668 87344 45670
rect 87400 45668 87406 45670
rect 87098 45659 87406 45668
rect 87834 45180 88142 45189
rect 87834 45178 87840 45180
rect 87896 45178 87920 45180
rect 87976 45178 88000 45180
rect 88056 45178 88080 45180
rect 88136 45178 88142 45180
rect 87896 45126 87898 45178
rect 88078 45126 88080 45178
rect 87834 45124 87840 45126
rect 87896 45124 87920 45126
rect 87976 45124 88000 45126
rect 88056 45124 88080 45126
rect 88136 45124 88142 45126
rect 87834 45115 88142 45124
rect 87098 44636 87406 44645
rect 87098 44634 87104 44636
rect 87160 44634 87184 44636
rect 87240 44634 87264 44636
rect 87320 44634 87344 44636
rect 87400 44634 87406 44636
rect 87160 44582 87162 44634
rect 87342 44582 87344 44634
rect 87098 44580 87104 44582
rect 87160 44580 87184 44582
rect 87240 44580 87264 44582
rect 87320 44580 87344 44582
rect 87400 44580 87406 44582
rect 87098 44571 87406 44580
rect 87834 44092 88142 44101
rect 87834 44090 87840 44092
rect 87896 44090 87920 44092
rect 87976 44090 88000 44092
rect 88056 44090 88080 44092
rect 88136 44090 88142 44092
rect 87896 44038 87898 44090
rect 88078 44038 88080 44090
rect 87834 44036 87840 44038
rect 87896 44036 87920 44038
rect 87976 44036 88000 44038
rect 88056 44036 88080 44038
rect 88136 44036 88142 44038
rect 87834 44027 88142 44036
rect 87098 43548 87406 43557
rect 87098 43546 87104 43548
rect 87160 43546 87184 43548
rect 87240 43546 87264 43548
rect 87320 43546 87344 43548
rect 87400 43546 87406 43548
rect 87160 43494 87162 43546
rect 87342 43494 87344 43546
rect 87098 43492 87104 43494
rect 87160 43492 87184 43494
rect 87240 43492 87264 43494
rect 87320 43492 87344 43494
rect 87400 43492 87406 43494
rect 87098 43483 87406 43492
rect 89940 43276 89992 43282
rect 89940 43218 89992 43224
rect 89952 43185 89980 43218
rect 89938 43176 89994 43185
rect 89938 43111 89994 43120
rect 87834 43004 88142 43013
rect 87834 43002 87840 43004
rect 87896 43002 87920 43004
rect 87976 43002 88000 43004
rect 88056 43002 88080 43004
rect 88136 43002 88142 43004
rect 87896 42950 87898 43002
rect 88078 42950 88080 43002
rect 87834 42948 87840 42950
rect 87896 42948 87920 42950
rect 87976 42948 88000 42950
rect 88056 42948 88080 42950
rect 88136 42948 88142 42950
rect 87834 42939 88142 42948
rect 87098 42460 87406 42469
rect 87098 42458 87104 42460
rect 87160 42458 87184 42460
rect 87240 42458 87264 42460
rect 87320 42458 87344 42460
rect 87400 42458 87406 42460
rect 87160 42406 87162 42458
rect 87342 42406 87344 42458
rect 87098 42404 87104 42406
rect 87160 42404 87184 42406
rect 87240 42404 87264 42406
rect 87320 42404 87344 42406
rect 87400 42404 87406 42406
rect 87098 42395 87406 42404
rect 88560 42154 88612 42160
rect 88560 42096 88612 42102
rect 87834 41916 88142 41925
rect 87834 41914 87840 41916
rect 87896 41914 87920 41916
rect 87976 41914 88000 41916
rect 88056 41914 88080 41916
rect 88136 41914 88142 41916
rect 87896 41862 87898 41914
rect 88078 41862 88080 41914
rect 87834 41860 87840 41862
rect 87896 41860 87920 41862
rect 87976 41860 88000 41862
rect 88056 41860 88080 41862
rect 88136 41860 88142 41862
rect 87834 41851 88142 41860
rect 88572 41825 88600 42096
rect 88558 41816 88614 41825
rect 87456 41780 87508 41786
rect 88558 41751 88614 41760
rect 87456 41722 87508 41728
rect 87098 41372 87406 41381
rect 87098 41370 87104 41372
rect 87160 41370 87184 41372
rect 87240 41370 87264 41372
rect 87320 41370 87344 41372
rect 87400 41370 87406 41372
rect 87160 41318 87162 41370
rect 87342 41318 87344 41370
rect 87098 41316 87104 41318
rect 87160 41316 87184 41318
rect 87240 41316 87264 41318
rect 87320 41316 87344 41318
rect 87400 41316 87406 41318
rect 87098 41307 87406 41316
rect 87468 40873 87496 41722
rect 89940 41712 89992 41718
rect 89940 41654 89992 41660
rect 89952 41145 89980 41654
rect 89938 41136 89994 41145
rect 89938 41071 89994 41080
rect 87454 40864 87510 40873
rect 87454 40799 87510 40808
rect 87834 40828 88142 40837
rect 87834 40826 87840 40828
rect 87896 40826 87920 40828
rect 87976 40826 88000 40828
rect 88056 40826 88080 40828
rect 88136 40826 88142 40828
rect 87896 40774 87898 40826
rect 88078 40774 88080 40826
rect 87834 40772 87840 40774
rect 87896 40772 87920 40774
rect 87976 40772 88000 40774
rect 88056 40772 88080 40774
rect 88136 40772 88142 40774
rect 87834 40763 88142 40772
rect 87098 40284 87406 40293
rect 87098 40282 87104 40284
rect 87160 40282 87184 40284
rect 87240 40282 87264 40284
rect 87320 40282 87344 40284
rect 87400 40282 87406 40284
rect 87160 40230 87162 40282
rect 87342 40230 87344 40282
rect 87098 40228 87104 40230
rect 87160 40228 87184 40230
rect 87240 40228 87264 40230
rect 87320 40228 87344 40230
rect 87400 40228 87406 40230
rect 87098 40219 87406 40228
rect 89940 39944 89992 39950
rect 89940 39886 89992 39892
rect 89952 39785 89980 39886
rect 89938 39776 89994 39785
rect 87834 39740 88142 39749
rect 87834 39738 87840 39740
rect 87896 39738 87920 39740
rect 87976 39738 88000 39740
rect 88056 39738 88080 39740
rect 88136 39738 88142 39740
rect 87896 39686 87898 39738
rect 88078 39686 88080 39738
rect 89938 39711 89994 39720
rect 87834 39684 87840 39686
rect 87896 39684 87920 39686
rect 87976 39684 88000 39686
rect 88056 39684 88080 39686
rect 88136 39684 88142 39686
rect 87834 39675 88142 39684
rect 87098 39196 87406 39205
rect 87098 39194 87104 39196
rect 87160 39194 87184 39196
rect 87240 39194 87264 39196
rect 87320 39194 87344 39196
rect 87400 39194 87406 39196
rect 87160 39142 87162 39194
rect 87342 39142 87344 39194
rect 87098 39140 87104 39142
rect 87160 39140 87184 39142
rect 87240 39140 87264 39142
rect 87320 39140 87344 39142
rect 87400 39140 87406 39142
rect 87098 39131 87406 39140
rect 87180 38992 87232 38998
rect 87180 38934 87232 38940
rect 87192 38697 87220 38934
rect 89296 38856 89348 38862
rect 89296 38798 89348 38804
rect 87178 38688 87234 38697
rect 87178 38623 87234 38632
rect 87834 38652 88142 38661
rect 87834 38650 87840 38652
rect 87896 38650 87920 38652
rect 87976 38650 88000 38652
rect 88056 38650 88080 38652
rect 88136 38650 88142 38652
rect 87896 38598 87898 38650
rect 88078 38598 88080 38650
rect 87834 38596 87840 38598
rect 87896 38596 87920 38598
rect 87976 38596 88000 38598
rect 88056 38596 88080 38598
rect 88136 38596 88142 38598
rect 87834 38587 88142 38596
rect 89308 38425 89336 38798
rect 89294 38416 89350 38425
rect 89294 38351 89350 38360
rect 87098 38108 87406 38117
rect 87098 38106 87104 38108
rect 87160 38106 87184 38108
rect 87240 38106 87264 38108
rect 87320 38106 87344 38108
rect 87400 38106 87406 38108
rect 87160 38054 87162 38106
rect 87342 38054 87344 38106
rect 87098 38052 87104 38054
rect 87160 38052 87184 38054
rect 87240 38052 87264 38054
rect 87320 38052 87344 38054
rect 87400 38052 87406 38054
rect 87098 38043 87406 38052
rect 89940 37768 89992 37774
rect 89938 37736 89940 37745
rect 89992 37736 89994 37745
rect 89938 37671 89994 37680
rect 87834 37564 88142 37573
rect 87834 37562 87840 37564
rect 87896 37562 87920 37564
rect 87976 37562 88000 37564
rect 88056 37562 88080 37564
rect 88136 37562 88142 37564
rect 87896 37510 87898 37562
rect 88078 37510 88080 37562
rect 87834 37508 87840 37510
rect 87896 37508 87920 37510
rect 87976 37508 88000 37510
rect 88056 37508 88080 37510
rect 88136 37508 88142 37510
rect 87834 37499 88142 37508
rect 87098 37020 87406 37029
rect 87098 37018 87104 37020
rect 87160 37018 87184 37020
rect 87240 37018 87264 37020
rect 87320 37018 87344 37020
rect 87400 37018 87406 37020
rect 87160 36966 87162 37018
rect 87342 36966 87344 37018
rect 87098 36964 87104 36966
rect 87160 36964 87184 36966
rect 87240 36964 87264 36966
rect 87320 36964 87344 36966
rect 87400 36964 87406 36966
rect 87098 36955 87406 36964
rect 89940 36680 89992 36686
rect 89940 36622 89992 36628
rect 87834 36476 88142 36485
rect 87834 36474 87840 36476
rect 87896 36474 87920 36476
rect 87976 36474 88000 36476
rect 88056 36474 88080 36476
rect 88136 36474 88142 36476
rect 87896 36422 87898 36474
rect 88078 36422 88080 36474
rect 87834 36420 87840 36422
rect 87896 36420 87920 36422
rect 87976 36420 88000 36422
rect 88056 36420 88080 36422
rect 88136 36420 88142 36422
rect 87834 36411 88142 36420
rect 89952 36385 89980 36622
rect 89938 36376 89994 36385
rect 89938 36311 89994 36320
rect 90124 36204 90176 36210
rect 90124 36146 90176 36152
rect 87456 36136 87508 36142
rect 87456 36078 87508 36084
rect 87098 35932 87406 35941
rect 87098 35930 87104 35932
rect 87160 35930 87184 35932
rect 87240 35930 87264 35932
rect 87320 35930 87344 35932
rect 87400 35930 87406 35932
rect 87160 35878 87162 35930
rect 87342 35878 87344 35930
rect 87098 35876 87104 35878
rect 87160 35876 87184 35878
rect 87240 35876 87264 35878
rect 87320 35876 87344 35878
rect 87400 35876 87406 35878
rect 87098 35867 87406 35876
rect 87468 35433 87496 36078
rect 90136 35705 90164 36146
rect 90122 35696 90178 35705
rect 90122 35631 90178 35640
rect 87454 35424 87510 35433
rect 87454 35359 87510 35368
rect 87834 35388 88142 35397
rect 87834 35386 87840 35388
rect 87896 35386 87920 35388
rect 87976 35386 88000 35388
rect 88056 35386 88080 35388
rect 88136 35386 88142 35388
rect 87896 35334 87898 35386
rect 88078 35334 88080 35386
rect 87834 35332 87840 35334
rect 87896 35332 87920 35334
rect 87976 35332 88000 35334
rect 88056 35332 88080 35334
rect 88136 35332 88142 35334
rect 87834 35323 88142 35332
rect 87098 34844 87406 34853
rect 87098 34842 87104 34844
rect 87160 34842 87184 34844
rect 87240 34842 87264 34844
rect 87320 34842 87344 34844
rect 87400 34842 87406 34844
rect 87160 34790 87162 34842
rect 87342 34790 87344 34842
rect 87098 34788 87104 34790
rect 87160 34788 87184 34790
rect 87240 34788 87264 34790
rect 87320 34788 87344 34790
rect 87400 34788 87406 34790
rect 87098 34779 87406 34788
rect 88560 34532 88612 34538
rect 88560 34474 88612 34480
rect 88572 34345 88600 34474
rect 88558 34336 88614 34345
rect 87834 34300 88142 34309
rect 87834 34298 87840 34300
rect 87896 34298 87920 34300
rect 87976 34298 88000 34300
rect 88056 34298 88080 34300
rect 88136 34298 88142 34300
rect 87896 34246 87898 34298
rect 88078 34246 88080 34298
rect 88558 34271 88614 34280
rect 87834 34244 87840 34246
rect 87896 34244 87920 34246
rect 87976 34244 88000 34246
rect 88056 34244 88080 34246
rect 88136 34244 88142 34246
rect 87834 34235 88142 34244
rect 87098 33756 87406 33765
rect 87098 33754 87104 33756
rect 87160 33754 87184 33756
rect 87240 33754 87264 33756
rect 87320 33754 87344 33756
rect 87400 33754 87406 33756
rect 87160 33702 87162 33754
rect 87342 33702 87344 33754
rect 87098 33700 87104 33702
rect 87160 33700 87184 33702
rect 87240 33700 87264 33702
rect 87320 33700 87344 33702
rect 87400 33700 87406 33702
rect 87098 33691 87406 33700
rect 87180 33416 87232 33422
rect 87180 33358 87232 33364
rect 89940 33416 89992 33422
rect 89940 33358 89992 33364
rect 87192 33257 87220 33358
rect 87178 33248 87234 33257
rect 87178 33183 87234 33192
rect 87834 33212 88142 33221
rect 87834 33210 87840 33212
rect 87896 33210 87920 33212
rect 87976 33210 88000 33212
rect 88056 33210 88080 33212
rect 88136 33210 88142 33212
rect 87896 33158 87898 33210
rect 88078 33158 88080 33210
rect 87834 33156 87840 33158
rect 87896 33156 87920 33158
rect 87976 33156 88000 33158
rect 88056 33156 88080 33158
rect 88136 33156 88142 33158
rect 87834 33147 88142 33156
rect 89952 32985 89980 33358
rect 89938 32976 89994 32985
rect 89938 32911 89994 32920
rect 87098 32668 87406 32677
rect 87098 32666 87104 32668
rect 87160 32666 87184 32668
rect 87240 32666 87264 32668
rect 87320 32666 87344 32668
rect 87400 32666 87406 32668
rect 87160 32614 87162 32666
rect 87342 32614 87344 32666
rect 87098 32612 87104 32614
rect 87160 32612 87184 32614
rect 87240 32612 87264 32614
rect 87320 32612 87344 32614
rect 87400 32612 87406 32614
rect 87098 32603 87406 32612
rect 89940 32328 89992 32334
rect 89938 32296 89940 32305
rect 89992 32296 89994 32305
rect 89938 32231 89994 32240
rect 87834 32124 88142 32133
rect 87834 32122 87840 32124
rect 87896 32122 87920 32124
rect 87976 32122 88000 32124
rect 88056 32122 88080 32124
rect 88136 32122 88142 32124
rect 87896 32070 87898 32122
rect 88078 32070 88080 32122
rect 87834 32068 87840 32070
rect 87896 32068 87920 32070
rect 87976 32068 88000 32070
rect 88056 32068 88080 32070
rect 88136 32068 88142 32070
rect 87834 32059 88142 32068
rect 87098 31580 87406 31589
rect 87098 31578 87104 31580
rect 87160 31578 87184 31580
rect 87240 31578 87264 31580
rect 87320 31578 87344 31580
rect 87400 31578 87406 31580
rect 87160 31526 87162 31578
rect 87342 31526 87344 31578
rect 87098 31524 87104 31526
rect 87160 31524 87184 31526
rect 87240 31524 87264 31526
rect 87320 31524 87344 31526
rect 87400 31524 87406 31526
rect 87098 31515 87406 31524
rect 88560 31268 88612 31274
rect 88560 31210 88612 31216
rect 87834 31036 88142 31045
rect 87834 31034 87840 31036
rect 87896 31034 87920 31036
rect 87976 31034 88000 31036
rect 88056 31034 88080 31036
rect 88136 31034 88142 31036
rect 87896 30982 87898 31034
rect 88078 30982 88080 31034
rect 87834 30980 87840 30982
rect 87896 30980 87920 30982
rect 87976 30980 88000 30982
rect 88056 30980 88080 30982
rect 88136 30980 88142 30982
rect 87834 30971 88142 30980
rect 88572 30945 88600 31210
rect 88558 30936 88614 30945
rect 88558 30871 88614 30880
rect 89940 30764 89992 30770
rect 89940 30706 89992 30712
rect 87456 30628 87508 30634
rect 87456 30570 87508 30576
rect 87098 30492 87406 30501
rect 87098 30490 87104 30492
rect 87160 30490 87184 30492
rect 87240 30490 87264 30492
rect 87320 30490 87344 30492
rect 87400 30490 87406 30492
rect 87160 30438 87162 30490
rect 87342 30438 87344 30490
rect 87098 30436 87104 30438
rect 87160 30436 87184 30438
rect 87240 30436 87264 30438
rect 87320 30436 87344 30438
rect 87400 30436 87406 30438
rect 87098 30427 87406 30436
rect 87468 30265 87496 30570
rect 89952 30265 89980 30706
rect 87454 30256 87510 30265
rect 87454 30191 87510 30200
rect 89938 30256 89994 30265
rect 89938 30191 89994 30200
rect 87834 29948 88142 29957
rect 87834 29946 87840 29948
rect 87896 29946 87920 29948
rect 87976 29946 88000 29948
rect 88056 29946 88080 29948
rect 88136 29946 88142 29948
rect 87896 29894 87898 29946
rect 88078 29894 88080 29946
rect 87834 29892 87840 29894
rect 87896 29892 87920 29894
rect 87976 29892 88000 29894
rect 88056 29892 88080 29894
rect 88136 29892 88142 29894
rect 87834 29883 88142 29892
rect 87098 29404 87406 29413
rect 87098 29402 87104 29404
rect 87160 29402 87184 29404
rect 87240 29402 87264 29404
rect 87320 29402 87344 29404
rect 87400 29402 87406 29404
rect 87160 29350 87162 29402
rect 87342 29350 87344 29402
rect 87098 29348 87104 29350
rect 87160 29348 87184 29350
rect 87240 29348 87264 29350
rect 87320 29348 87344 29350
rect 87400 29348 87406 29350
rect 87098 29339 87406 29348
rect 88560 29092 88612 29098
rect 88560 29034 88612 29040
rect 88572 28905 88600 29034
rect 88558 28896 88614 28905
rect 87834 28860 88142 28869
rect 87834 28858 87840 28860
rect 87896 28858 87920 28860
rect 87976 28858 88000 28860
rect 88056 28858 88080 28860
rect 88136 28858 88142 28860
rect 87896 28806 87898 28858
rect 88078 28806 88080 28858
rect 88558 28831 88614 28840
rect 87834 28804 87840 28806
rect 87896 28804 87920 28806
rect 87976 28804 88000 28806
rect 88056 28804 88080 28806
rect 88136 28804 88142 28806
rect 87834 28795 88142 28804
rect 87098 28316 87406 28325
rect 87098 28314 87104 28316
rect 87160 28314 87184 28316
rect 87240 28314 87264 28316
rect 87320 28314 87344 28316
rect 87400 28314 87406 28316
rect 87160 28262 87162 28314
rect 87342 28262 87344 28314
rect 87098 28260 87104 28262
rect 87160 28260 87184 28262
rect 87240 28260 87264 28262
rect 87320 28260 87344 28262
rect 87400 28260 87406 28262
rect 87098 28251 87406 28260
rect 87548 27976 87600 27982
rect 87548 27918 87600 27924
rect 87560 27817 87588 27918
rect 89940 27908 89992 27914
rect 89940 27850 89992 27856
rect 87546 27808 87602 27817
rect 87546 27743 87602 27752
rect 87834 27772 88142 27781
rect 87834 27770 87840 27772
rect 87896 27770 87920 27772
rect 87976 27770 88000 27772
rect 88056 27770 88080 27772
rect 88136 27770 88142 27772
rect 87896 27718 87898 27770
rect 88078 27718 88080 27770
rect 87834 27716 87840 27718
rect 87896 27716 87920 27718
rect 87976 27716 88000 27718
rect 88056 27716 88080 27718
rect 88136 27716 88142 27718
rect 87834 27707 88142 27716
rect 89952 27545 89980 27850
rect 89938 27536 89994 27545
rect 89938 27471 89994 27480
rect 87098 27228 87406 27237
rect 87098 27226 87104 27228
rect 87160 27226 87184 27228
rect 87240 27226 87264 27228
rect 87320 27226 87344 27228
rect 87400 27226 87406 27228
rect 87160 27174 87162 27226
rect 87342 27174 87344 27226
rect 87098 27172 87104 27174
rect 87160 27172 87184 27174
rect 87240 27172 87264 27174
rect 87320 27172 87344 27174
rect 87400 27172 87406 27174
rect 87098 27163 87406 27172
rect 89938 26856 89994 26865
rect 89938 26791 89940 26800
rect 89992 26791 89994 26800
rect 89940 26762 89992 26768
rect 87834 26684 88142 26693
rect 87834 26682 87840 26684
rect 87896 26682 87920 26684
rect 87976 26682 88000 26684
rect 88056 26682 88080 26684
rect 88136 26682 88142 26684
rect 87896 26630 87898 26682
rect 88078 26630 88080 26682
rect 87834 26628 87840 26630
rect 87896 26628 87920 26630
rect 87976 26628 88000 26630
rect 88056 26628 88080 26630
rect 88136 26628 88142 26630
rect 87834 26619 88142 26628
rect 87098 26140 87406 26149
rect 87098 26138 87104 26140
rect 87160 26138 87184 26140
rect 87240 26138 87264 26140
rect 87320 26138 87344 26140
rect 87400 26138 87406 26140
rect 87160 26086 87162 26138
rect 87342 26086 87344 26138
rect 87098 26084 87104 26086
rect 87160 26084 87184 26086
rect 87240 26084 87264 26086
rect 87320 26084 87344 26086
rect 87400 26084 87406 26086
rect 87098 26075 87406 26084
rect 89940 25732 89992 25738
rect 89940 25674 89992 25680
rect 87834 25596 88142 25605
rect 87834 25594 87840 25596
rect 87896 25594 87920 25596
rect 87976 25594 88000 25596
rect 88056 25594 88080 25596
rect 88136 25594 88142 25596
rect 87896 25542 87898 25594
rect 88078 25542 88080 25594
rect 87834 25540 87840 25542
rect 87896 25540 87920 25542
rect 87976 25540 88000 25542
rect 88056 25540 88080 25542
rect 88136 25540 88142 25542
rect 87834 25531 88142 25540
rect 89952 25505 89980 25674
rect 89938 25496 89994 25505
rect 89938 25431 89994 25440
rect 88376 25358 88428 25364
rect 88376 25300 88428 25306
rect 87098 25052 87406 25061
rect 87098 25050 87104 25052
rect 87160 25050 87184 25052
rect 87240 25050 87264 25052
rect 87320 25050 87344 25052
rect 87400 25050 87406 25052
rect 87160 24998 87162 25050
rect 87342 24998 87344 25050
rect 87098 24996 87104 24998
rect 87160 24996 87184 24998
rect 87240 24996 87264 24998
rect 87320 24996 87344 24998
rect 87400 24996 87406 24998
rect 87098 24987 87406 24996
rect 88388 24825 88416 25300
rect 89940 25188 89992 25194
rect 89940 25130 89992 25136
rect 89952 24825 89980 25130
rect 88374 24816 88430 24825
rect 88374 24751 88430 24760
rect 89938 24816 89994 24825
rect 89938 24751 89994 24760
rect 87834 24508 88142 24517
rect 87834 24506 87840 24508
rect 87896 24506 87920 24508
rect 87976 24506 88000 24508
rect 88056 24506 88080 24508
rect 88136 24506 88142 24508
rect 87896 24454 87898 24506
rect 88078 24454 88080 24506
rect 87834 24452 87840 24454
rect 87896 24452 87920 24454
rect 87976 24452 88000 24454
rect 88056 24452 88080 24454
rect 88136 24452 88142 24454
rect 87834 24443 88142 24452
rect 87098 23964 87406 23973
rect 87098 23962 87104 23964
rect 87160 23962 87184 23964
rect 87240 23962 87264 23964
rect 87320 23962 87344 23964
rect 87400 23962 87406 23964
rect 87160 23910 87162 23962
rect 87342 23910 87344 23962
rect 87098 23908 87104 23910
rect 87160 23908 87184 23910
rect 87240 23908 87264 23910
rect 87320 23908 87344 23910
rect 87400 23908 87406 23910
rect 87098 23899 87406 23908
rect 89940 23556 89992 23562
rect 89940 23498 89992 23504
rect 89952 23465 89980 23498
rect 89938 23456 89994 23465
rect 87834 23420 88142 23429
rect 87834 23418 87840 23420
rect 87896 23418 87920 23420
rect 87976 23418 88000 23420
rect 88056 23418 88080 23420
rect 88136 23418 88142 23420
rect 87896 23366 87898 23418
rect 88078 23366 88080 23418
rect 89938 23391 89994 23400
rect 87834 23364 87840 23366
rect 87896 23364 87920 23366
rect 87976 23364 88000 23366
rect 88056 23364 88080 23366
rect 88136 23364 88142 23366
rect 87834 23355 88142 23364
rect 87098 22876 87406 22885
rect 87098 22874 87104 22876
rect 87160 22874 87184 22876
rect 87240 22874 87264 22876
rect 87320 22874 87344 22876
rect 87400 22874 87406 22876
rect 87160 22822 87162 22874
rect 87342 22822 87344 22874
rect 87098 22820 87104 22822
rect 87160 22820 87184 22822
rect 87240 22820 87264 22822
rect 87320 22820 87344 22822
rect 87400 22820 87406 22822
rect 87098 22811 87406 22820
rect 89940 22468 89992 22474
rect 89940 22410 89992 22416
rect 87834 22332 88142 22341
rect 87834 22330 87840 22332
rect 87896 22330 87920 22332
rect 87976 22330 88000 22332
rect 88056 22330 88080 22332
rect 88136 22330 88142 22332
rect 87896 22278 87898 22330
rect 88078 22278 88080 22330
rect 87834 22276 87840 22278
rect 87896 22276 87920 22278
rect 87976 22276 88000 22278
rect 88056 22276 88080 22278
rect 88136 22276 88142 22278
rect 87834 22267 88142 22276
rect 89952 22105 89980 22410
rect 89938 22096 89994 22105
rect 89938 22031 89994 22040
rect 87098 21788 87406 21797
rect 87098 21786 87104 21788
rect 87160 21786 87184 21788
rect 87240 21786 87264 21788
rect 87320 21786 87344 21788
rect 87400 21786 87406 21788
rect 87160 21734 87162 21786
rect 87342 21734 87344 21786
rect 87098 21732 87104 21734
rect 87160 21732 87184 21734
rect 87240 21732 87264 21734
rect 87320 21732 87344 21734
rect 87400 21732 87406 21734
rect 87098 21723 87406 21732
rect 89938 21416 89994 21425
rect 89938 21351 89940 21360
rect 89992 21351 89994 21360
rect 89940 21322 89992 21328
rect 87834 21244 88142 21253
rect 87834 21242 87840 21244
rect 87896 21242 87920 21244
rect 87976 21242 88000 21244
rect 88056 21242 88080 21244
rect 88136 21242 88142 21244
rect 87896 21190 87898 21242
rect 88078 21190 88080 21242
rect 87834 21188 87840 21190
rect 87896 21188 87920 21190
rect 87976 21188 88000 21190
rect 88056 21188 88080 21190
rect 88136 21188 88142 21190
rect 87834 21179 88142 21188
rect 87098 20700 87406 20709
rect 87098 20698 87104 20700
rect 87160 20698 87184 20700
rect 87240 20698 87264 20700
rect 87320 20698 87344 20700
rect 87400 20698 87406 20700
rect 87160 20646 87162 20698
rect 87342 20646 87344 20698
rect 87098 20644 87104 20646
rect 87160 20644 87184 20646
rect 87240 20644 87264 20646
rect 87320 20644 87344 20646
rect 87400 20644 87406 20646
rect 87098 20635 87406 20644
rect 89940 20292 89992 20298
rect 89940 20234 89992 20240
rect 87834 20156 88142 20165
rect 87834 20154 87840 20156
rect 87896 20154 87920 20156
rect 87976 20154 88000 20156
rect 88056 20154 88080 20156
rect 88136 20154 88142 20156
rect 87896 20102 87898 20154
rect 88078 20102 88080 20154
rect 87834 20100 87840 20102
rect 87896 20100 87920 20102
rect 87976 20100 88000 20102
rect 88056 20100 88080 20102
rect 88136 20100 88142 20102
rect 87834 20091 88142 20100
rect 89952 20065 89980 20234
rect 89938 20056 89994 20065
rect 89938 19991 89994 20000
rect 88376 19918 88428 19924
rect 88376 19860 88428 19866
rect 87098 19612 87406 19621
rect 87098 19610 87104 19612
rect 87160 19610 87184 19612
rect 87240 19610 87264 19612
rect 87320 19610 87344 19612
rect 87400 19610 87406 19612
rect 87160 19558 87162 19610
rect 87342 19558 87344 19610
rect 87098 19556 87104 19558
rect 87160 19556 87184 19558
rect 87240 19556 87264 19558
rect 87320 19556 87344 19558
rect 87400 19556 87406 19558
rect 87098 19547 87406 19556
rect 88388 19385 88416 19860
rect 90032 19748 90084 19754
rect 90032 19690 90084 19696
rect 90044 19385 90072 19690
rect 88374 19376 88430 19385
rect 88374 19311 88430 19320
rect 90030 19376 90086 19385
rect 90030 19311 90086 19320
rect 87834 19068 88142 19077
rect 87834 19066 87840 19068
rect 87896 19066 87920 19068
rect 87976 19066 88000 19068
rect 88056 19066 88080 19068
rect 88136 19066 88142 19068
rect 87896 19014 87898 19066
rect 88078 19014 88080 19066
rect 87834 19012 87840 19014
rect 87896 19012 87920 19014
rect 87976 19012 88000 19014
rect 88056 19012 88080 19014
rect 88136 19012 88142 19014
rect 87834 19003 88142 19012
rect 87098 18524 87406 18533
rect 87098 18522 87104 18524
rect 87160 18522 87184 18524
rect 87240 18522 87264 18524
rect 87320 18522 87344 18524
rect 87400 18522 87406 18524
rect 87160 18470 87162 18522
rect 87342 18470 87344 18522
rect 87098 18468 87104 18470
rect 87160 18468 87184 18470
rect 87240 18468 87264 18470
rect 87320 18468 87344 18470
rect 87400 18468 87406 18470
rect 87098 18459 87406 18468
rect 89940 18252 89992 18258
rect 88192 18218 88244 18224
rect 89940 18194 89992 18200
rect 88192 18161 88244 18166
rect 88190 18152 88246 18161
rect 88190 18087 88246 18096
rect 89952 18025 89980 18194
rect 89938 18016 89994 18025
rect 87834 17980 88142 17989
rect 87834 17978 87840 17980
rect 87896 17978 87920 17980
rect 87976 17978 88000 17980
rect 88056 17978 88080 17980
rect 88136 17978 88142 17980
rect 87896 17926 87898 17978
rect 88078 17926 88080 17978
rect 89938 17951 89994 17960
rect 87834 17924 87840 17926
rect 87896 17924 87920 17926
rect 87976 17924 88000 17926
rect 88056 17924 88080 17926
rect 88136 17924 88142 17926
rect 87834 17915 88142 17924
rect 87098 17436 87406 17445
rect 87098 17434 87104 17436
rect 87160 17434 87184 17436
rect 87240 17434 87264 17436
rect 87320 17434 87344 17436
rect 87400 17434 87406 17436
rect 87160 17382 87162 17434
rect 87342 17382 87344 17434
rect 87098 17380 87104 17382
rect 87160 17380 87184 17382
rect 87240 17380 87264 17382
rect 87320 17380 87344 17382
rect 87400 17380 87406 17382
rect 87098 17371 87406 17380
rect 89940 17028 89992 17034
rect 89940 16970 89992 16976
rect 87834 16892 88142 16901
rect 87834 16890 87840 16892
rect 87896 16890 87920 16892
rect 87976 16890 88000 16892
rect 88056 16890 88080 16892
rect 88136 16890 88142 16892
rect 87896 16838 87898 16890
rect 88078 16838 88080 16890
rect 87834 16836 87840 16838
rect 87896 16836 87920 16838
rect 87976 16836 88000 16838
rect 88056 16836 88080 16838
rect 88136 16836 88142 16838
rect 87834 16827 88142 16836
rect 89952 16665 89980 16970
rect 89938 16656 89994 16665
rect 89938 16591 89994 16600
rect 87098 16348 87406 16357
rect 87098 16346 87104 16348
rect 87160 16346 87184 16348
rect 87240 16346 87264 16348
rect 87320 16346 87344 16348
rect 87400 16346 87406 16348
rect 87160 16294 87162 16346
rect 87342 16294 87344 16346
rect 87098 16292 87104 16294
rect 87160 16292 87184 16294
rect 87240 16292 87264 16294
rect 87320 16292 87344 16294
rect 87400 16292 87406 16294
rect 87098 16283 87406 16292
rect 89938 15976 89994 15985
rect 89938 15911 89940 15920
rect 89992 15911 89994 15920
rect 89940 15882 89992 15888
rect 87834 15804 88142 15813
rect 87834 15802 87840 15804
rect 87896 15802 87920 15804
rect 87976 15802 88000 15804
rect 88056 15802 88080 15804
rect 88136 15802 88142 15804
rect 87896 15750 87898 15802
rect 88078 15750 88080 15802
rect 87834 15748 87840 15750
rect 87896 15748 87920 15750
rect 87976 15748 88000 15750
rect 88056 15748 88080 15750
rect 88136 15748 88142 15750
rect 87834 15739 88142 15748
rect 87098 15260 87406 15269
rect 87098 15258 87104 15260
rect 87160 15258 87184 15260
rect 87240 15258 87264 15260
rect 87320 15258 87344 15260
rect 87400 15258 87406 15260
rect 87160 15206 87162 15258
rect 87342 15206 87344 15258
rect 87098 15204 87104 15206
rect 87160 15204 87184 15206
rect 87240 15204 87264 15206
rect 87320 15204 87344 15206
rect 87400 15204 87406 15206
rect 87098 15195 87406 15204
rect 89940 14852 89992 14858
rect 89940 14794 89992 14800
rect 87834 14716 88142 14725
rect 87834 14714 87840 14716
rect 87896 14714 87920 14716
rect 87976 14714 88000 14716
rect 88056 14714 88080 14716
rect 88136 14714 88142 14716
rect 87896 14662 87898 14714
rect 88078 14662 88080 14714
rect 87834 14660 87840 14662
rect 87896 14660 87920 14662
rect 87976 14660 88000 14662
rect 88056 14660 88080 14662
rect 88136 14660 88142 14662
rect 87834 14651 88142 14660
rect 89952 14625 89980 14794
rect 89938 14616 89994 14625
rect 89938 14551 89994 14560
rect 88376 14478 88428 14484
rect 88376 14420 88428 14426
rect 87098 14172 87406 14181
rect 87098 14170 87104 14172
rect 87160 14170 87184 14172
rect 87240 14170 87264 14172
rect 87320 14170 87344 14172
rect 87400 14170 87406 14172
rect 87160 14118 87162 14170
rect 87342 14118 87344 14170
rect 87098 14116 87104 14118
rect 87160 14116 87184 14118
rect 87240 14116 87264 14118
rect 87320 14116 87344 14118
rect 87400 14116 87406 14118
rect 87098 14107 87406 14116
rect 88388 13945 88416 14420
rect 89940 14308 89992 14314
rect 89940 14250 89992 14256
rect 89952 13945 89980 14250
rect 88374 13936 88430 13945
rect 88374 13871 88430 13880
rect 89938 13936 89994 13945
rect 89938 13871 89994 13880
rect 87834 13628 88142 13637
rect 87834 13626 87840 13628
rect 87896 13626 87920 13628
rect 87976 13626 88000 13628
rect 88056 13626 88080 13628
rect 88136 13626 88142 13628
rect 87896 13574 87898 13626
rect 88078 13574 88080 13626
rect 87834 13572 87840 13574
rect 87896 13572 87920 13574
rect 87976 13572 88000 13574
rect 88056 13572 88080 13574
rect 88136 13572 88142 13574
rect 87834 13563 88142 13572
rect 87098 13084 87406 13093
rect 87098 13082 87104 13084
rect 87160 13082 87184 13084
rect 87240 13082 87264 13084
rect 87320 13082 87344 13084
rect 87400 13082 87406 13084
rect 87160 13030 87162 13082
rect 87342 13030 87344 13082
rect 87098 13028 87104 13030
rect 87160 13028 87184 13030
rect 87240 13028 87264 13030
rect 87320 13028 87344 13030
rect 87400 13028 87406 13030
rect 87098 13019 87406 13028
rect 87834 12540 88142 12549
rect 87834 12538 87840 12540
rect 87896 12538 87920 12540
rect 87976 12538 88000 12540
rect 88056 12538 88080 12540
rect 88136 12538 88142 12540
rect 87896 12486 87898 12538
rect 88078 12486 88080 12538
rect 87834 12484 87840 12486
rect 87896 12484 87920 12486
rect 87976 12484 88000 12486
rect 88056 12484 88080 12486
rect 88136 12484 88142 12486
rect 87834 12475 88142 12484
rect 87098 11996 87406 12005
rect 87098 11994 87104 11996
rect 87160 11994 87184 11996
rect 87240 11994 87264 11996
rect 87320 11994 87344 11996
rect 87400 11994 87406 11996
rect 87160 11942 87162 11994
rect 87342 11942 87344 11994
rect 87098 11940 87104 11942
rect 87160 11940 87184 11942
rect 87240 11940 87264 11942
rect 87320 11940 87344 11942
rect 87400 11940 87406 11942
rect 87098 11931 87406 11940
rect 87834 11452 88142 11461
rect 87834 11450 87840 11452
rect 87896 11450 87920 11452
rect 87976 11450 88000 11452
rect 88056 11450 88080 11452
rect 88136 11450 88142 11452
rect 87896 11398 87898 11450
rect 88078 11398 88080 11450
rect 87834 11396 87840 11398
rect 87896 11396 87920 11398
rect 87976 11396 88000 11398
rect 88056 11396 88080 11398
rect 88136 11396 88142 11398
rect 87834 11387 88142 11396
rect 87098 10908 87406 10917
rect 87098 10906 87104 10908
rect 87160 10906 87184 10908
rect 87240 10906 87264 10908
rect 87320 10906 87344 10908
rect 87400 10906 87406 10908
rect 87160 10854 87162 10906
rect 87342 10854 87344 10906
rect 87098 10852 87104 10854
rect 87160 10852 87184 10854
rect 87240 10852 87264 10854
rect 87320 10852 87344 10854
rect 87400 10852 87406 10854
rect 87098 10843 87406 10852
rect 87834 10364 88142 10373
rect 87834 10362 87840 10364
rect 87896 10362 87920 10364
rect 87976 10362 88000 10364
rect 88056 10362 88080 10364
rect 88136 10362 88142 10364
rect 87896 10310 87898 10362
rect 88078 10310 88080 10362
rect 87834 10308 87840 10310
rect 87896 10308 87920 10310
rect 87976 10308 88000 10310
rect 88056 10308 88080 10310
rect 88136 10308 88142 10310
rect 87834 10299 88142 10308
rect 84418 10264 84474 10273
rect 84418 10199 84474 10208
rect 46698 9992 46754 10001
rect 46698 9927 46754 9936
rect 48138 9842 48166 10100
rect 49090 9992 49146 10001
rect 49090 9927 49146 9936
rect 38736 9814 38828 9842
rect 24356 5168 24384 9814
rect 25460 5168 25488 9814
rect 26564 5168 26592 9814
rect 27668 5168 27696 9814
rect 28772 5168 28800 9814
rect 29876 5168 29904 9814
rect 30980 5338 31008 9814
rect 30968 5332 31020 5338
rect 30968 5274 31020 5280
rect 32084 5270 32112 9814
rect 33188 5338 33216 9814
rect 34292 5338 34320 9814
rect 35396 5338 35424 9814
rect 36500 5338 36528 9814
rect 37604 5338 37632 9814
rect 37722 7644 38030 7653
rect 37722 7642 37728 7644
rect 37784 7642 37808 7644
rect 37864 7642 37888 7644
rect 37944 7642 37968 7644
rect 38024 7642 38030 7644
rect 37784 7590 37786 7642
rect 37966 7590 37968 7642
rect 37722 7588 37728 7590
rect 37784 7588 37808 7590
rect 37864 7588 37888 7590
rect 37944 7588 37968 7590
rect 38024 7588 38030 7590
rect 37722 7579 38030 7588
rect 38382 7100 38690 7109
rect 38382 7098 38388 7100
rect 38444 7098 38468 7100
rect 38524 7098 38548 7100
rect 38604 7098 38628 7100
rect 38684 7098 38690 7100
rect 38444 7046 38446 7098
rect 38626 7046 38628 7098
rect 38382 7044 38388 7046
rect 38444 7044 38468 7046
rect 38524 7044 38548 7046
rect 38604 7044 38628 7046
rect 38684 7044 38690 7046
rect 38382 7035 38690 7044
rect 37722 6556 38030 6565
rect 37722 6554 37728 6556
rect 37784 6554 37808 6556
rect 37864 6554 37888 6556
rect 37944 6554 37968 6556
rect 38024 6554 38030 6556
rect 37784 6502 37786 6554
rect 37966 6502 37968 6554
rect 37722 6500 37728 6502
rect 37784 6500 37808 6502
rect 37864 6500 37888 6502
rect 37944 6500 37968 6502
rect 38024 6500 38030 6502
rect 37722 6491 38030 6500
rect 38382 6012 38690 6021
rect 38382 6010 38388 6012
rect 38444 6010 38468 6012
rect 38524 6010 38548 6012
rect 38604 6010 38628 6012
rect 38684 6010 38690 6012
rect 38444 5958 38446 6010
rect 38626 5958 38628 6010
rect 38382 5956 38388 5958
rect 38444 5956 38468 5958
rect 38524 5956 38548 5958
rect 38604 5956 38628 5958
rect 38684 5956 38690 5958
rect 38382 5947 38690 5956
rect 37722 5468 38030 5477
rect 37722 5466 37728 5468
rect 37784 5466 37808 5468
rect 37864 5466 37888 5468
rect 37944 5466 37968 5468
rect 38024 5466 38030 5468
rect 37784 5414 37786 5466
rect 37966 5414 37968 5466
rect 37722 5412 37728 5414
rect 37784 5412 37808 5414
rect 37864 5412 37888 5414
rect 37944 5412 37968 5414
rect 38024 5412 38030 5414
rect 37722 5403 38030 5412
rect 38800 5338 38828 9814
rect 39812 9814 39868 9842
rect 40916 9814 40972 9842
rect 42020 9814 42076 9842
rect 43124 9814 43180 9842
rect 44228 9814 44284 9842
rect 45332 9814 45388 9842
rect 48092 9814 48166 9842
rect 49104 9842 49132 9927
rect 49242 9842 49270 10100
rect 50194 9992 50250 10001
rect 50194 9927 50250 9936
rect 49104 9814 49270 9842
rect 50208 9842 50236 9927
rect 50346 9842 50374 10100
rect 50208 9814 50374 9842
rect 51450 9842 51478 10100
rect 51574 9992 51630 10001
rect 51574 9927 51630 9936
rect 51588 9842 51616 9927
rect 51450 9814 51616 9842
rect 52554 9842 52582 10100
rect 53658 9842 53686 10100
rect 54762 9842 54790 10100
rect 55866 9842 55894 10100
rect 52554 9814 52628 9842
rect 53658 9814 53732 9842
rect 54762 9814 54836 9842
rect 33176 5332 33228 5338
rect 33176 5274 33228 5280
rect 34280 5332 34332 5338
rect 34280 5274 34332 5280
rect 35384 5332 35436 5338
rect 35384 5274 35436 5280
rect 36488 5332 36540 5338
rect 36488 5274 36540 5280
rect 37592 5332 37644 5338
rect 37592 5274 37644 5280
rect 38788 5332 38840 5338
rect 38788 5274 38840 5280
rect 39812 5270 39840 9814
rect 40916 5338 40944 9814
rect 40904 5332 40956 5338
rect 40904 5274 40956 5280
rect 42020 5270 42048 9814
rect 43124 5270 43152 9814
rect 44228 5338 44256 9814
rect 45332 5338 45360 9814
rect 48092 8505 48120 9814
rect 48078 8496 48134 8505
rect 48078 8431 48134 8440
rect 44216 5332 44268 5338
rect 44216 5274 44268 5280
rect 45320 5332 45372 5338
rect 45320 5274 45372 5280
rect 32072 5264 32124 5270
rect 32072 5206 32124 5212
rect 39800 5264 39852 5270
rect 39800 5206 39852 5212
rect 42008 5264 42060 5270
rect 42008 5206 42060 5212
rect 43112 5264 43164 5270
rect 43112 5206 43164 5212
rect 44124 5196 44176 5202
rect 15512 5138 15564 5144
rect 16616 5162 16668 5168
rect 12568 5128 12620 5134
rect 12568 5070 12620 5076
rect 13856 5128 13908 5134
rect 13856 5070 13908 5076
rect 14500 5128 14552 5134
rect 14500 5070 14552 5076
rect 15420 5128 15472 5134
rect 16616 5104 16668 5110
rect 17720 5162 17772 5168
rect 17720 5104 17772 5110
rect 19100 5162 19152 5168
rect 19100 5104 19152 5110
rect 19928 5162 19980 5168
rect 19928 5104 19980 5110
rect 21032 5162 21084 5168
rect 21032 5104 21084 5110
rect 22136 5162 22188 5168
rect 22136 5104 22188 5110
rect 23332 5162 23384 5168
rect 23332 5104 23384 5110
rect 24344 5162 24396 5168
rect 24344 5104 24396 5110
rect 25448 5162 25500 5168
rect 25448 5104 25500 5110
rect 26552 5162 26604 5168
rect 26552 5104 26604 5110
rect 27656 5162 27708 5168
rect 27656 5104 27708 5110
rect 28760 5162 28812 5168
rect 28760 5104 28812 5110
rect 29864 5162 29916 5168
rect 31888 5162 31940 5168
rect 29864 5104 29916 5110
rect 31244 5156 31296 5162
rect 35108 5162 35160 5168
rect 34464 5136 34516 5142
rect 31888 5104 31940 5110
rect 33176 5128 33228 5134
rect 31244 5098 31296 5104
rect 15420 5070 15472 5076
rect 12580 2400 12608 5070
rect 13868 2400 13896 5070
rect 14512 2400 14540 5070
rect 15788 5060 15840 5066
rect 15788 5002 15840 5008
rect 16432 5060 16484 5066
rect 16432 5002 16484 5008
rect 17720 5060 17772 5066
rect 17720 5002 17772 5008
rect 19008 5060 19060 5066
rect 19008 5002 19060 5008
rect 19744 5060 19796 5066
rect 19744 5002 19796 5008
rect 20940 5060 20992 5066
rect 20940 5002 20992 5008
rect 22228 5060 22280 5066
rect 22228 5002 22280 5008
rect 23516 5060 23568 5066
rect 23516 5002 23568 5008
rect 24160 5060 24212 5066
rect 24160 5002 24212 5008
rect 25448 5060 25500 5066
rect 25448 5002 25500 5008
rect 26736 5060 26788 5066
rect 26736 5002 26788 5008
rect 27380 5060 27432 5066
rect 27380 5002 27432 5008
rect 28668 5060 28720 5066
rect 28668 5002 28720 5008
rect 29956 5060 30008 5066
rect 29956 5002 30008 5008
rect 15800 2400 15828 5002
rect 16444 2400 16472 5002
rect 17732 2400 17760 5002
rect 19020 2400 19048 5002
rect 19382 4924 19690 4933
rect 19382 4922 19388 4924
rect 19444 4922 19468 4924
rect 19524 4922 19548 4924
rect 19604 4922 19628 4924
rect 19684 4922 19690 4924
rect 19444 4870 19446 4922
rect 19626 4870 19628 4922
rect 19382 4868 19388 4870
rect 19444 4868 19468 4870
rect 19524 4868 19548 4870
rect 19604 4868 19628 4870
rect 19684 4868 19690 4870
rect 19382 4859 19690 4868
rect 19756 3314 19784 5002
rect 19664 3286 19784 3314
rect 19664 2400 19692 3286
rect 20952 2400 20980 5002
rect 22240 2400 22268 5002
rect 23528 2400 23556 5002
rect 24172 2400 24200 5002
rect 25460 2400 25488 5002
rect 26748 2400 26776 5002
rect 27392 2400 27420 5002
rect 28680 2400 28708 5002
rect 29968 2400 29996 5002
rect 31256 2400 31284 5098
rect 31900 2400 31928 5104
rect 35108 5104 35160 5110
rect 36396 5162 36448 5168
rect 39616 5162 39668 5168
rect 36396 5104 36448 5110
rect 37684 5156 37736 5162
rect 34464 5078 34516 5084
rect 33176 5070 33228 5076
rect 33188 2400 33216 5070
rect 34476 2400 34504 5078
rect 35120 2400 35148 5104
rect 36408 2400 36436 5104
rect 37684 5098 37736 5104
rect 38972 5156 39024 5162
rect 44124 5138 44176 5144
rect 45412 5196 45464 5202
rect 52600 5168 52628 9814
rect 53704 5168 53732 9814
rect 54808 5168 54836 9814
rect 55820 9814 55894 9842
rect 56970 9842 56998 10100
rect 58074 9842 58102 10100
rect 59178 9842 59206 10100
rect 56970 9814 57136 9842
rect 58074 9814 58240 9842
rect 55820 5168 55848 9814
rect 56722 7644 57030 7653
rect 56722 7642 56728 7644
rect 56784 7642 56808 7644
rect 56864 7642 56888 7644
rect 56944 7642 56968 7644
rect 57024 7642 57030 7644
rect 56784 7590 56786 7642
rect 56966 7590 56968 7642
rect 56722 7588 56728 7590
rect 56784 7588 56808 7590
rect 56864 7588 56888 7590
rect 56944 7588 56968 7590
rect 57024 7588 57030 7590
rect 56722 7579 57030 7588
rect 56722 6556 57030 6565
rect 56722 6554 56728 6556
rect 56784 6554 56808 6556
rect 56864 6554 56888 6556
rect 56944 6554 56968 6556
rect 57024 6554 57030 6556
rect 56784 6502 56786 6554
rect 56966 6502 56968 6554
rect 56722 6500 56728 6502
rect 56784 6500 56808 6502
rect 56864 6500 56888 6502
rect 56944 6500 56968 6502
rect 57024 6500 57030 6502
rect 56722 6491 57030 6500
rect 56722 5468 57030 5477
rect 56722 5466 56728 5468
rect 56784 5466 56808 5468
rect 56864 5466 56888 5468
rect 56944 5466 56968 5468
rect 57024 5466 57030 5468
rect 56784 5414 56786 5466
rect 56966 5414 56968 5466
rect 56722 5412 56728 5414
rect 56784 5412 56808 5414
rect 56864 5412 56888 5414
rect 56944 5412 56968 5414
rect 57024 5412 57030 5414
rect 56722 5403 57030 5412
rect 57108 5168 57136 9814
rect 57382 7100 57690 7109
rect 57382 7098 57388 7100
rect 57444 7098 57468 7100
rect 57524 7098 57548 7100
rect 57604 7098 57628 7100
rect 57684 7098 57690 7100
rect 57444 7046 57446 7098
rect 57626 7046 57628 7098
rect 57382 7044 57388 7046
rect 57444 7044 57468 7046
rect 57524 7044 57548 7046
rect 57604 7044 57628 7046
rect 57684 7044 57690 7046
rect 57382 7035 57690 7044
rect 57382 6012 57690 6021
rect 57382 6010 57388 6012
rect 57444 6010 57468 6012
rect 57524 6010 57548 6012
rect 57604 6010 57628 6012
rect 57684 6010 57690 6012
rect 57444 5958 57446 6010
rect 57626 5958 57628 6010
rect 57382 5956 57388 5958
rect 57444 5956 57468 5958
rect 57524 5956 57548 5958
rect 57604 5956 57628 5958
rect 57684 5956 57690 5958
rect 57382 5947 57690 5956
rect 58212 5168 58240 9814
rect 59132 9814 59206 9842
rect 60282 9842 60310 10100
rect 61386 9842 61414 10100
rect 62490 9842 62518 10100
rect 63594 9842 63622 10100
rect 60282 9814 60356 9842
rect 61386 9814 61460 9842
rect 62490 9814 62564 9842
rect 59132 5168 59160 9814
rect 60328 5168 60356 9814
rect 61432 5168 61460 9814
rect 62536 5168 62564 9814
rect 63548 9814 63622 9842
rect 64698 9842 64726 10100
rect 65802 9842 65830 10100
rect 66906 9842 66934 10100
rect 64698 9814 64772 9842
rect 65802 9814 65876 9842
rect 63548 5168 63576 9814
rect 64744 5168 64772 9814
rect 65848 5168 65876 9814
rect 66860 9814 66934 9842
rect 68010 9842 68038 10100
rect 69114 9842 69142 10100
rect 70218 9842 70246 10100
rect 68010 9814 68084 9842
rect 69114 9814 69372 9842
rect 66860 5168 66888 9814
rect 68056 5338 68084 9814
rect 69344 5338 69372 9814
rect 70172 9814 70246 9842
rect 71322 9842 71350 10100
rect 72426 9842 72454 10100
rect 73530 9842 73558 10100
rect 74634 9842 74662 10100
rect 75738 9842 75766 10100
rect 71322 9814 71396 9842
rect 72426 9814 72500 9842
rect 73530 9814 73604 9842
rect 74634 9814 74800 9842
rect 70172 5338 70200 9814
rect 68044 5332 68096 5338
rect 68044 5274 68096 5280
rect 69332 5332 69384 5338
rect 69332 5274 69384 5280
rect 70160 5332 70212 5338
rect 70160 5274 70212 5280
rect 71368 5270 71396 9814
rect 72472 5338 72500 9814
rect 73576 5338 73604 9814
rect 74772 5338 74800 9814
rect 75600 9814 75766 9842
rect 76842 9842 76870 10100
rect 77946 9842 77974 10100
rect 76842 9814 76916 9842
rect 75600 5338 75628 9814
rect 75722 7644 76030 7653
rect 75722 7642 75728 7644
rect 75784 7642 75808 7644
rect 75864 7642 75888 7644
rect 75944 7642 75968 7644
rect 76024 7642 76030 7644
rect 75784 7590 75786 7642
rect 75966 7590 75968 7642
rect 75722 7588 75728 7590
rect 75784 7588 75808 7590
rect 75864 7588 75888 7590
rect 75944 7588 75968 7590
rect 76024 7588 76030 7590
rect 75722 7579 76030 7588
rect 76382 7100 76690 7109
rect 76382 7098 76388 7100
rect 76444 7098 76468 7100
rect 76524 7098 76548 7100
rect 76604 7098 76628 7100
rect 76684 7098 76690 7100
rect 76444 7046 76446 7098
rect 76626 7046 76628 7098
rect 76382 7044 76388 7046
rect 76444 7044 76468 7046
rect 76524 7044 76548 7046
rect 76604 7044 76628 7046
rect 76684 7044 76690 7046
rect 76382 7035 76690 7044
rect 75722 6556 76030 6565
rect 75722 6554 75728 6556
rect 75784 6554 75808 6556
rect 75864 6554 75888 6556
rect 75944 6554 75968 6556
rect 76024 6554 76030 6556
rect 75784 6502 75786 6554
rect 75966 6502 75968 6554
rect 75722 6500 75728 6502
rect 75784 6500 75808 6502
rect 75864 6500 75888 6502
rect 75944 6500 75968 6502
rect 76024 6500 76030 6502
rect 75722 6491 76030 6500
rect 76382 6012 76690 6021
rect 76382 6010 76388 6012
rect 76444 6010 76468 6012
rect 76524 6010 76548 6012
rect 76604 6010 76628 6012
rect 76684 6010 76690 6012
rect 76444 5958 76446 6010
rect 76626 5958 76628 6010
rect 76382 5956 76388 5958
rect 76444 5956 76468 5958
rect 76524 5956 76548 5958
rect 76604 5956 76628 5958
rect 76684 5956 76690 5958
rect 76382 5947 76690 5956
rect 75722 5468 76030 5477
rect 75722 5466 75728 5468
rect 75784 5466 75808 5468
rect 75864 5466 75888 5468
rect 75944 5466 75968 5468
rect 76024 5466 76030 5468
rect 75784 5414 75786 5466
rect 75966 5414 75968 5466
rect 75722 5412 75728 5414
rect 75784 5412 75808 5414
rect 75864 5412 75888 5414
rect 75944 5412 75968 5414
rect 76024 5412 76030 5414
rect 75722 5403 76030 5412
rect 76888 5338 76916 9814
rect 77900 9814 77974 9842
rect 79050 9842 79078 10100
rect 80154 9842 80182 10100
rect 81258 9842 81286 10100
rect 82362 9842 82390 10100
rect 79050 9814 79124 9842
rect 80154 9814 80320 9842
rect 81258 9814 81700 9842
rect 82362 9814 82436 9842
rect 77900 5338 77928 9814
rect 72460 5332 72512 5338
rect 72460 5274 72512 5280
rect 73564 5332 73616 5338
rect 73564 5274 73616 5280
rect 74760 5332 74812 5338
rect 74760 5274 74812 5280
rect 75588 5332 75640 5338
rect 75588 5274 75640 5280
rect 76876 5332 76928 5338
rect 76876 5274 76928 5280
rect 77888 5332 77940 5338
rect 77888 5274 77940 5280
rect 79096 5270 79124 9814
rect 80292 5270 80320 9814
rect 81672 5338 81700 9814
rect 82120 5740 82172 5746
rect 82120 5682 82172 5688
rect 81660 5332 81712 5338
rect 81660 5274 81712 5280
rect 71356 5264 71408 5270
rect 71356 5206 71408 5212
rect 79084 5264 79136 5270
rect 79084 5206 79136 5212
rect 80280 5264 80332 5270
rect 80280 5206 80332 5212
rect 81476 5196 81528 5202
rect 45412 5138 45464 5144
rect 52588 5162 52640 5168
rect 39616 5104 39668 5110
rect 40904 5128 40956 5134
rect 38972 5098 39024 5104
rect 37696 2400 37724 5098
rect 38382 4924 38690 4933
rect 38382 4922 38388 4924
rect 38444 4922 38468 4924
rect 38524 4922 38548 4924
rect 38604 4922 38628 4924
rect 38684 4922 38690 4924
rect 38444 4870 38446 4922
rect 38626 4870 38628 4922
rect 38382 4868 38388 4870
rect 38444 4868 38468 4870
rect 38524 4868 38548 4870
rect 38604 4868 38628 4870
rect 38684 4868 38690 4870
rect 38382 4859 38690 4868
rect 38984 2400 39012 5098
rect 39628 2400 39656 5104
rect 40904 5070 40956 5076
rect 42192 5128 42244 5134
rect 42192 5070 42244 5076
rect 42836 5128 42888 5134
rect 42836 5070 42888 5076
rect 40916 2400 40944 5070
rect 42204 2400 42232 5070
rect 42848 2400 42876 5070
rect 44136 2400 44164 5138
rect 45424 2400 45452 5138
rect 52588 5104 52640 5110
rect 53692 5162 53744 5168
rect 53692 5104 53744 5110
rect 54796 5162 54848 5168
rect 54796 5104 54848 5110
rect 55808 5162 55860 5168
rect 55808 5104 55860 5110
rect 57096 5162 57148 5168
rect 57096 5104 57148 5110
rect 58200 5162 58252 5168
rect 58200 5104 58252 5110
rect 59120 5162 59172 5168
rect 59120 5104 59172 5110
rect 60316 5162 60368 5168
rect 60316 5104 60368 5110
rect 61420 5162 61472 5168
rect 61420 5104 61472 5110
rect 62524 5162 62576 5168
rect 62524 5104 62576 5110
rect 63536 5162 63588 5168
rect 63536 5104 63588 5110
rect 64732 5162 64784 5168
rect 64732 5104 64784 5110
rect 65836 5162 65888 5168
rect 65836 5104 65888 5110
rect 66848 5162 66900 5168
rect 69884 5162 69936 5168
rect 66848 5104 66900 5110
rect 67952 5136 68004 5142
rect 67952 5078 68004 5084
rect 69240 5128 69292 5134
rect 52496 5060 52548 5066
rect 52496 5002 52548 5008
rect 53784 5060 53836 5066
rect 53784 5002 53836 5008
rect 54428 5060 54480 5066
rect 54428 5002 54480 5008
rect 55716 5060 55768 5066
rect 55716 5002 55768 5008
rect 57004 5060 57056 5066
rect 57004 5002 57056 5008
rect 58292 5060 58344 5066
rect 58292 5002 58344 5008
rect 58936 5060 58988 5066
rect 58936 5002 58988 5008
rect 60224 5060 60276 5066
rect 60224 5002 60276 5008
rect 61512 5060 61564 5066
rect 61512 5002 61564 5008
rect 62156 5060 62208 5066
rect 62156 5002 62208 5008
rect 63444 5060 63496 5066
rect 63444 5002 63496 5008
rect 64732 5060 64784 5066
rect 64732 5002 64784 5008
rect 66020 5060 66072 5066
rect 66020 5002 66072 5008
rect 66664 5060 66716 5066
rect 66664 5002 66716 5008
rect 52508 2400 52536 5002
rect 53796 2400 53824 5002
rect 54440 2400 54468 5002
rect 55728 2400 55756 5002
rect 57016 2400 57044 5002
rect 57382 4924 57690 4933
rect 57382 4922 57388 4924
rect 57444 4922 57468 4924
rect 57524 4922 57548 4924
rect 57604 4922 57628 4924
rect 57684 4922 57690 4924
rect 57444 4870 57446 4922
rect 57626 4870 57628 4922
rect 57382 4868 57388 4870
rect 57444 4868 57468 4870
rect 57524 4868 57548 4870
rect 57604 4868 57628 4870
rect 57684 4868 57690 4870
rect 57382 4859 57690 4868
rect 58304 2400 58332 5002
rect 58948 2400 58976 5002
rect 60236 2400 60264 5002
rect 61524 2400 61552 5002
rect 62168 2400 62196 5002
rect 63456 2400 63484 5002
rect 64744 2400 64772 5002
rect 66032 2400 66060 5002
rect 66676 2400 66704 5002
rect 67964 2400 67992 5078
rect 69884 5104 69936 5110
rect 71172 5162 71224 5168
rect 74392 5162 74444 5168
rect 71172 5104 71224 5110
rect 72460 5156 72512 5162
rect 69240 5070 69292 5076
rect 69252 2400 69280 5070
rect 69896 2400 69924 5104
rect 71184 2400 71212 5104
rect 72460 5098 72512 5104
rect 73748 5156 73800 5162
rect 77612 5162 77664 5168
rect 74392 5104 74444 5110
rect 75680 5136 75732 5142
rect 73748 5098 73800 5104
rect 72472 2400 72500 5098
rect 73760 2400 73788 5098
rect 74404 2400 74432 5104
rect 75680 5078 75732 5084
rect 76968 5128 77020 5134
rect 75692 2400 75720 5078
rect 81476 5138 81528 5144
rect 77612 5104 77664 5110
rect 78900 5128 78952 5134
rect 76968 5070 77020 5076
rect 76382 4924 76690 4933
rect 76382 4922 76388 4924
rect 76444 4922 76468 4924
rect 76524 4922 76548 4924
rect 76604 4922 76628 4924
rect 76684 4922 76690 4924
rect 76444 4870 76446 4922
rect 76626 4870 76628 4922
rect 76382 4868 76388 4870
rect 76444 4868 76468 4870
rect 76524 4868 76548 4870
rect 76604 4868 76628 4870
rect 76684 4868 76690 4870
rect 76382 4859 76690 4868
rect 76980 2400 77008 5070
rect 77624 2400 77652 5104
rect 78900 5070 78952 5076
rect 80188 5128 80240 5134
rect 80188 5070 80240 5076
rect 78912 2400 78940 5070
rect 80200 2400 80228 5070
rect 81488 2400 81516 5138
rect 82132 2400 82160 5682
rect 82408 5678 82436 9814
rect 87098 9820 87406 9829
rect 87098 9818 87104 9820
rect 87160 9818 87184 9820
rect 87240 9818 87264 9820
rect 87320 9818 87344 9820
rect 87400 9818 87406 9820
rect 87160 9766 87162 9818
rect 87342 9766 87344 9818
rect 87098 9764 87104 9766
rect 87160 9764 87184 9766
rect 87240 9764 87264 9766
rect 87320 9764 87344 9766
rect 87400 9764 87406 9766
rect 87098 9755 87406 9764
rect 87834 9276 88142 9285
rect 87834 9274 87840 9276
rect 87896 9274 87920 9276
rect 87976 9274 88000 9276
rect 88056 9274 88080 9276
rect 88136 9274 88142 9276
rect 87896 9222 87898 9274
rect 88078 9222 88080 9274
rect 87834 9220 87840 9222
rect 87896 9220 87920 9222
rect 87976 9220 88000 9222
rect 88056 9220 88080 9222
rect 88136 9220 88142 9222
rect 87834 9211 88142 9220
rect 87098 8732 87406 8741
rect 87098 8730 87104 8732
rect 87160 8730 87184 8732
rect 87240 8730 87264 8732
rect 87320 8730 87344 8732
rect 87400 8730 87406 8732
rect 87160 8678 87162 8730
rect 87342 8678 87344 8730
rect 87098 8676 87104 8678
rect 87160 8676 87184 8678
rect 87240 8676 87264 8678
rect 87320 8676 87344 8678
rect 87400 8676 87406 8678
rect 87098 8667 87406 8676
rect 87834 8188 88142 8197
rect 87834 8186 87840 8188
rect 87896 8186 87920 8188
rect 87976 8186 88000 8188
rect 88056 8186 88080 8188
rect 88136 8186 88142 8188
rect 87896 8134 87898 8186
rect 88078 8134 88080 8186
rect 87834 8132 87840 8134
rect 87896 8132 87920 8134
rect 87976 8132 88000 8134
rect 88056 8132 88080 8134
rect 88136 8132 88142 8134
rect 87834 8123 88142 8132
rect 87098 7644 87406 7653
rect 87098 7642 87104 7644
rect 87160 7642 87184 7644
rect 87240 7642 87264 7644
rect 87320 7642 87344 7644
rect 87400 7642 87406 7644
rect 87160 7590 87162 7642
rect 87342 7590 87344 7642
rect 87098 7588 87104 7590
rect 87160 7588 87184 7590
rect 87240 7588 87264 7590
rect 87320 7588 87344 7590
rect 87400 7588 87406 7590
rect 87098 7579 87406 7588
rect 87834 7100 88142 7109
rect 87834 7098 87840 7100
rect 87896 7098 87920 7100
rect 87976 7098 88000 7100
rect 88056 7098 88080 7100
rect 88136 7098 88142 7100
rect 87896 7046 87898 7098
rect 88078 7046 88080 7098
rect 87834 7044 87840 7046
rect 87896 7044 87920 7046
rect 87976 7044 88000 7046
rect 88056 7044 88080 7046
rect 88136 7044 88142 7046
rect 87834 7035 88142 7044
rect 82396 5672 82448 5678
rect 82396 5614 82448 5620
rect 1618 1600 1674 2400
rect 2262 1600 2318 2400
rect 2906 1600 2962 2400
rect 3550 1600 3606 2400
rect 4194 1600 4250 2400
rect 4838 1600 4894 2400
rect 5482 1600 5538 2400
rect 6126 1600 6182 2400
rect 6770 1600 6826 2400
rect 7414 1600 7470 2400
rect 8058 1600 8114 2400
rect 8702 1600 8758 2400
rect 9346 1600 9402 2400
rect 9990 1600 10046 2400
rect 10634 1600 10690 2400
rect 11278 1600 11334 2400
rect 12566 1600 12622 2400
rect 13854 1600 13910 2400
rect 14498 1600 14554 2400
rect 15786 1600 15842 2400
rect 16430 1600 16486 2400
rect 17718 1600 17774 2400
rect 19006 1600 19062 2400
rect 19650 1600 19706 2400
rect 20938 1600 20994 2400
rect 22226 1600 22282 2400
rect 23514 1600 23570 2400
rect 24158 1600 24214 2400
rect 25446 1600 25502 2400
rect 26734 1600 26790 2400
rect 27378 1600 27434 2400
rect 28666 1600 28722 2400
rect 29954 1600 30010 2400
rect 31242 1600 31298 2400
rect 31886 1600 31942 2400
rect 33174 1600 33230 2400
rect 34462 1600 34518 2400
rect 35106 1600 35162 2400
rect 36394 1600 36450 2400
rect 37682 1600 37738 2400
rect 38970 1600 39026 2400
rect 39614 1600 39670 2400
rect 40902 1600 40958 2400
rect 42190 1600 42246 2400
rect 42834 1600 42890 2400
rect 44122 1600 44178 2400
rect 45410 1600 45466 2400
rect 52494 1600 52550 2400
rect 53782 1600 53838 2400
rect 54426 1600 54482 2400
rect 55714 1600 55770 2400
rect 57002 1600 57058 2400
rect 58290 1600 58346 2400
rect 58934 1600 58990 2400
rect 60222 1600 60278 2400
rect 61510 1600 61566 2400
rect 62154 1600 62210 2400
rect 63442 1600 63498 2400
rect 64730 1600 64786 2400
rect 66018 1600 66074 2400
rect 66662 1600 66718 2400
rect 67950 1600 68006 2400
rect 69238 1600 69294 2400
rect 69882 1600 69938 2400
rect 71170 1600 71226 2400
rect 72458 1600 72514 2400
rect 73746 1600 73802 2400
rect 74390 1600 74446 2400
rect 75678 1600 75734 2400
rect 76966 1600 77022 2400
rect 77610 1600 77666 2400
rect 78898 1600 78954 2400
rect 80186 1600 80242 2400
rect 81474 1600 81530 2400
rect 82118 1600 82174 2400
<< via2 >>
rect 18728 89242 18784 89244
rect 18808 89242 18864 89244
rect 18888 89242 18944 89244
rect 18968 89242 19024 89244
rect 18728 89190 18774 89242
rect 18774 89190 18784 89242
rect 18808 89190 18838 89242
rect 18838 89190 18850 89242
rect 18850 89190 18864 89242
rect 18888 89190 18902 89242
rect 18902 89190 18914 89242
rect 18914 89190 18944 89242
rect 18968 89190 18978 89242
rect 18978 89190 19024 89242
rect 18728 89188 18784 89190
rect 18808 89188 18864 89190
rect 18888 89188 18944 89190
rect 18968 89188 19024 89190
rect 37728 89242 37784 89244
rect 37808 89242 37864 89244
rect 37888 89242 37944 89244
rect 37968 89242 38024 89244
rect 37728 89190 37774 89242
rect 37774 89190 37784 89242
rect 37808 89190 37838 89242
rect 37838 89190 37850 89242
rect 37850 89190 37864 89242
rect 37888 89190 37902 89242
rect 37902 89190 37914 89242
rect 37914 89190 37944 89242
rect 37968 89190 37978 89242
rect 37978 89190 38024 89242
rect 37728 89188 37784 89190
rect 37808 89188 37864 89190
rect 37888 89188 37944 89190
rect 37968 89188 38024 89190
rect 5960 87066 6016 87068
rect 6040 87066 6096 87068
rect 6120 87066 6176 87068
rect 6200 87066 6256 87068
rect 5960 87014 6006 87066
rect 6006 87014 6016 87066
rect 6040 87014 6070 87066
rect 6070 87014 6082 87066
rect 6082 87014 6096 87066
rect 6120 87014 6134 87066
rect 6134 87014 6146 87066
rect 6146 87014 6176 87066
rect 6200 87014 6210 87066
rect 6210 87014 6256 87066
rect 5960 87012 6016 87014
rect 6040 87012 6096 87014
rect 6120 87012 6176 87014
rect 6200 87012 6256 87014
rect 6696 86522 6752 86524
rect 6776 86522 6832 86524
rect 6856 86522 6912 86524
rect 6936 86522 6992 86524
rect 6696 86470 6742 86522
rect 6742 86470 6752 86522
rect 6776 86470 6806 86522
rect 6806 86470 6818 86522
rect 6818 86470 6832 86522
rect 6856 86470 6870 86522
rect 6870 86470 6882 86522
rect 6882 86470 6912 86522
rect 6936 86470 6946 86522
rect 6946 86470 6992 86522
rect 6696 86468 6752 86470
rect 6776 86468 6832 86470
rect 6856 86468 6912 86470
rect 6936 86468 6992 86470
rect 5960 85978 6016 85980
rect 6040 85978 6096 85980
rect 6120 85978 6176 85980
rect 6200 85978 6256 85980
rect 5960 85926 6006 85978
rect 6006 85926 6016 85978
rect 6040 85926 6070 85978
rect 6070 85926 6082 85978
rect 6082 85926 6096 85978
rect 6120 85926 6134 85978
rect 6134 85926 6146 85978
rect 6146 85926 6176 85978
rect 6200 85926 6210 85978
rect 6210 85926 6256 85978
rect 5960 85924 6016 85926
rect 6040 85924 6096 85926
rect 6120 85924 6176 85926
rect 6200 85924 6256 85926
rect 6696 85434 6752 85436
rect 6776 85434 6832 85436
rect 6856 85434 6912 85436
rect 6936 85434 6992 85436
rect 6696 85382 6742 85434
rect 6742 85382 6752 85434
rect 6776 85382 6806 85434
rect 6806 85382 6818 85434
rect 6818 85382 6832 85434
rect 6856 85382 6870 85434
rect 6870 85382 6882 85434
rect 6882 85382 6912 85434
rect 6936 85382 6946 85434
rect 6946 85382 6992 85434
rect 6696 85380 6752 85382
rect 6776 85380 6832 85382
rect 6856 85380 6912 85382
rect 6936 85380 6992 85382
rect 5960 84890 6016 84892
rect 6040 84890 6096 84892
rect 6120 84890 6176 84892
rect 6200 84890 6256 84892
rect 5960 84838 6006 84890
rect 6006 84838 6016 84890
rect 6040 84838 6070 84890
rect 6070 84838 6082 84890
rect 6082 84838 6096 84890
rect 6120 84838 6134 84890
rect 6134 84838 6146 84890
rect 6146 84838 6176 84890
rect 6200 84838 6210 84890
rect 6210 84838 6256 84890
rect 5960 84836 6016 84838
rect 6040 84836 6096 84838
rect 6120 84836 6176 84838
rect 6200 84836 6256 84838
rect 6696 84346 6752 84348
rect 6776 84346 6832 84348
rect 6856 84346 6912 84348
rect 6936 84346 6992 84348
rect 6696 84294 6742 84346
rect 6742 84294 6752 84346
rect 6776 84294 6806 84346
rect 6806 84294 6818 84346
rect 6818 84294 6832 84346
rect 6856 84294 6870 84346
rect 6870 84294 6882 84346
rect 6882 84294 6912 84346
rect 6936 84294 6946 84346
rect 6946 84294 6992 84346
rect 6696 84292 6752 84294
rect 6776 84292 6832 84294
rect 6856 84292 6912 84294
rect 6936 84292 6992 84294
rect 5960 83802 6016 83804
rect 6040 83802 6096 83804
rect 6120 83802 6176 83804
rect 6200 83802 6256 83804
rect 5960 83750 6006 83802
rect 6006 83750 6016 83802
rect 6040 83750 6070 83802
rect 6070 83750 6082 83802
rect 6082 83750 6096 83802
rect 6120 83750 6134 83802
rect 6134 83750 6146 83802
rect 6146 83750 6176 83802
rect 6200 83750 6210 83802
rect 6210 83750 6256 83802
rect 5960 83748 6016 83750
rect 6040 83748 6096 83750
rect 6120 83748 6176 83750
rect 6200 83748 6256 83750
rect 6696 83258 6752 83260
rect 6776 83258 6832 83260
rect 6856 83258 6912 83260
rect 6936 83258 6992 83260
rect 6696 83206 6742 83258
rect 6742 83206 6752 83258
rect 6776 83206 6806 83258
rect 6806 83206 6818 83258
rect 6818 83206 6832 83258
rect 6856 83206 6870 83258
rect 6870 83206 6882 83258
rect 6882 83206 6912 83258
rect 6936 83206 6946 83258
rect 6946 83206 6992 83258
rect 6696 83204 6752 83206
rect 6776 83204 6832 83206
rect 6856 83204 6912 83206
rect 6936 83204 6992 83206
rect 5960 82714 6016 82716
rect 6040 82714 6096 82716
rect 6120 82714 6176 82716
rect 6200 82714 6256 82716
rect 5960 82662 6006 82714
rect 6006 82662 6016 82714
rect 6040 82662 6070 82714
rect 6070 82662 6082 82714
rect 6082 82662 6096 82714
rect 6120 82662 6134 82714
rect 6134 82662 6146 82714
rect 6146 82662 6176 82714
rect 6200 82662 6210 82714
rect 6210 82662 6256 82714
rect 5960 82660 6016 82662
rect 6040 82660 6096 82662
rect 6120 82660 6176 82662
rect 6200 82660 6256 82662
rect 6696 82170 6752 82172
rect 6776 82170 6832 82172
rect 6856 82170 6912 82172
rect 6936 82170 6992 82172
rect 6696 82118 6742 82170
rect 6742 82118 6752 82170
rect 6776 82118 6806 82170
rect 6806 82118 6818 82170
rect 6818 82118 6832 82170
rect 6856 82118 6870 82170
rect 6870 82118 6882 82170
rect 6882 82118 6912 82170
rect 6936 82118 6946 82170
rect 6946 82118 6992 82170
rect 6696 82116 6752 82118
rect 6776 82116 6832 82118
rect 6856 82116 6912 82118
rect 6936 82116 6992 82118
rect 5960 81626 6016 81628
rect 6040 81626 6096 81628
rect 6120 81626 6176 81628
rect 6200 81626 6256 81628
rect 5960 81574 6006 81626
rect 6006 81574 6016 81626
rect 6040 81574 6070 81626
rect 6070 81574 6082 81626
rect 6082 81574 6096 81626
rect 6120 81574 6134 81626
rect 6134 81574 6146 81626
rect 6146 81574 6176 81626
rect 6200 81574 6210 81626
rect 6210 81574 6256 81626
rect 5960 81572 6016 81574
rect 6040 81572 6096 81574
rect 6120 81572 6176 81574
rect 6200 81572 6256 81574
rect 6696 81082 6752 81084
rect 6776 81082 6832 81084
rect 6856 81082 6912 81084
rect 6936 81082 6992 81084
rect 6696 81030 6742 81082
rect 6742 81030 6752 81082
rect 6776 81030 6806 81082
rect 6806 81030 6818 81082
rect 6818 81030 6832 81082
rect 6856 81030 6870 81082
rect 6870 81030 6882 81082
rect 6882 81030 6912 81082
rect 6936 81030 6946 81082
rect 6946 81030 6992 81082
rect 6696 81028 6752 81030
rect 6776 81028 6832 81030
rect 6856 81028 6912 81030
rect 6936 81028 6992 81030
rect 2906 80520 2962 80576
rect 5960 80538 6016 80540
rect 6040 80538 6096 80540
rect 6120 80538 6176 80540
rect 6200 80538 6256 80540
rect 5960 80486 6006 80538
rect 6006 80486 6016 80538
rect 6040 80486 6070 80538
rect 6070 80486 6082 80538
rect 6082 80486 6096 80538
rect 6120 80486 6134 80538
rect 6134 80486 6146 80538
rect 6146 80486 6176 80538
rect 6200 80486 6210 80538
rect 6210 80486 6256 80538
rect 5960 80484 6016 80486
rect 6040 80484 6096 80486
rect 6120 80484 6176 80486
rect 6200 80484 6256 80486
rect 7138 80384 7194 80440
rect 6696 79994 6752 79996
rect 6776 79994 6832 79996
rect 6856 79994 6912 79996
rect 6936 79994 6992 79996
rect 6696 79942 6742 79994
rect 6742 79942 6752 79994
rect 6776 79942 6806 79994
rect 6806 79942 6818 79994
rect 6818 79942 6832 79994
rect 6856 79942 6870 79994
rect 6870 79942 6882 79994
rect 6882 79942 6912 79994
rect 6936 79942 6946 79994
rect 6946 79942 6992 79994
rect 6696 79940 6752 79942
rect 6776 79940 6832 79942
rect 6856 79940 6912 79942
rect 6936 79940 6992 79942
rect 5960 79450 6016 79452
rect 6040 79450 6096 79452
rect 6120 79450 6176 79452
rect 6200 79450 6256 79452
rect 5960 79398 6006 79450
rect 6006 79398 6016 79450
rect 6040 79398 6070 79450
rect 6070 79398 6082 79450
rect 6082 79398 6096 79450
rect 6120 79398 6134 79450
rect 6134 79398 6146 79450
rect 6146 79398 6176 79450
rect 6200 79398 6210 79450
rect 6210 79398 6256 79450
rect 5960 79396 6016 79398
rect 6040 79396 6096 79398
rect 6120 79396 6176 79398
rect 6200 79396 6256 79398
rect 7138 79296 7194 79352
rect 2722 79160 2778 79216
rect 6696 78906 6752 78908
rect 6776 78906 6832 78908
rect 6856 78906 6912 78908
rect 6936 78906 6992 78908
rect 6696 78854 6742 78906
rect 6742 78854 6752 78906
rect 6776 78854 6806 78906
rect 6806 78854 6818 78906
rect 6818 78854 6832 78906
rect 6856 78854 6870 78906
rect 6870 78854 6882 78906
rect 6882 78854 6912 78906
rect 6936 78854 6946 78906
rect 6946 78854 6992 78906
rect 6696 78852 6752 78854
rect 6776 78852 6832 78854
rect 6856 78852 6912 78854
rect 6936 78852 6992 78854
rect 2906 78500 2962 78536
rect 2906 78480 2908 78500
rect 2908 78480 2960 78500
rect 2960 78480 2962 78500
rect 5960 78362 6016 78364
rect 6040 78362 6096 78364
rect 6120 78362 6176 78364
rect 6200 78362 6256 78364
rect 5960 78310 6006 78362
rect 6006 78310 6016 78362
rect 6040 78310 6070 78362
rect 6070 78310 6082 78362
rect 6082 78310 6096 78362
rect 6120 78310 6134 78362
rect 6134 78310 6146 78362
rect 6146 78310 6176 78362
rect 6200 78310 6210 78362
rect 6210 78310 6256 78362
rect 5960 78308 6016 78310
rect 6040 78308 6096 78310
rect 6120 78308 6176 78310
rect 6200 78308 6256 78310
rect 7138 78208 7194 78264
rect 6696 77818 6752 77820
rect 6776 77818 6832 77820
rect 6856 77818 6912 77820
rect 6936 77818 6992 77820
rect 6696 77766 6742 77818
rect 6742 77766 6752 77818
rect 6776 77766 6806 77818
rect 6806 77766 6818 77818
rect 6818 77766 6832 77818
rect 6856 77766 6870 77818
rect 6870 77766 6882 77818
rect 6882 77766 6912 77818
rect 6936 77766 6946 77818
rect 6946 77766 6992 77818
rect 6696 77764 6752 77766
rect 6776 77764 6832 77766
rect 6856 77764 6912 77766
rect 6936 77764 6992 77766
rect 4378 77120 4434 77176
rect 5960 77274 6016 77276
rect 6040 77274 6096 77276
rect 6120 77274 6176 77276
rect 6200 77274 6256 77276
rect 5960 77222 6006 77274
rect 6006 77222 6016 77274
rect 6040 77222 6070 77274
rect 6070 77222 6082 77274
rect 6082 77222 6096 77274
rect 6120 77222 6134 77274
rect 6134 77222 6146 77274
rect 6146 77222 6176 77274
rect 6200 77222 6210 77274
rect 6210 77222 6256 77274
rect 5960 77220 6016 77222
rect 6040 77220 6096 77222
rect 6120 77220 6176 77222
rect 6200 77220 6256 77222
rect 5666 76984 5722 77040
rect 6696 76730 6752 76732
rect 6776 76730 6832 76732
rect 6856 76730 6912 76732
rect 6936 76730 6992 76732
rect 6696 76678 6742 76730
rect 6742 76678 6752 76730
rect 6776 76678 6806 76730
rect 6806 76678 6818 76730
rect 6818 76678 6832 76730
rect 6856 76678 6870 76730
rect 6870 76678 6882 76730
rect 6882 76678 6912 76730
rect 6936 76678 6946 76730
rect 6946 76678 6992 76730
rect 6696 76676 6752 76678
rect 6776 76676 6832 76678
rect 6856 76676 6912 76678
rect 6936 76676 6992 76678
rect 5960 76186 6016 76188
rect 6040 76186 6096 76188
rect 6120 76186 6176 76188
rect 6200 76186 6256 76188
rect 5960 76134 6006 76186
rect 6006 76134 6016 76186
rect 6040 76134 6070 76186
rect 6070 76134 6082 76186
rect 6082 76134 6096 76186
rect 6120 76134 6134 76186
rect 6134 76134 6146 76186
rect 6146 76134 6176 76186
rect 6200 76134 6210 76186
rect 6210 76134 6256 76186
rect 5960 76132 6016 76134
rect 6040 76132 6096 76134
rect 6120 76132 6176 76134
rect 6200 76132 6256 76134
rect 7138 76032 7194 76088
rect 2906 75780 2962 75816
rect 2906 75760 2908 75780
rect 2908 75760 2960 75780
rect 2960 75760 2962 75780
rect 6696 75642 6752 75644
rect 6776 75642 6832 75644
rect 6856 75642 6912 75644
rect 6936 75642 6992 75644
rect 6696 75590 6742 75642
rect 6742 75590 6752 75642
rect 6776 75590 6806 75642
rect 6806 75590 6818 75642
rect 6818 75590 6832 75642
rect 6856 75590 6870 75642
rect 6870 75590 6882 75642
rect 6882 75590 6912 75642
rect 6936 75590 6946 75642
rect 6946 75590 6992 75642
rect 6696 75588 6752 75590
rect 6776 75588 6832 75590
rect 6856 75588 6912 75590
rect 6936 75588 6992 75590
rect 2906 75080 2962 75136
rect 5960 75098 6016 75100
rect 6040 75098 6096 75100
rect 6120 75098 6176 75100
rect 6200 75098 6256 75100
rect 5960 75046 6006 75098
rect 6006 75046 6016 75098
rect 6040 75046 6070 75098
rect 6070 75046 6082 75098
rect 6082 75046 6096 75098
rect 6120 75046 6134 75098
rect 6134 75046 6146 75098
rect 6146 75046 6176 75098
rect 6200 75046 6210 75098
rect 6210 75046 6256 75098
rect 5960 75044 6016 75046
rect 6040 75044 6096 75046
rect 6120 75044 6176 75046
rect 6200 75044 6256 75046
rect 7138 74944 7194 75000
rect 6696 74554 6752 74556
rect 6776 74554 6832 74556
rect 6856 74554 6912 74556
rect 6936 74554 6992 74556
rect 6696 74502 6742 74554
rect 6742 74502 6752 74554
rect 6776 74502 6806 74554
rect 6806 74502 6818 74554
rect 6818 74502 6832 74554
rect 6856 74502 6870 74554
rect 6870 74502 6882 74554
rect 6882 74502 6912 74554
rect 6936 74502 6946 74554
rect 6946 74502 6992 74554
rect 6696 74500 6752 74502
rect 6776 74500 6832 74502
rect 6856 74500 6912 74502
rect 6936 74500 6992 74502
rect 5960 74010 6016 74012
rect 6040 74010 6096 74012
rect 6120 74010 6176 74012
rect 6200 74010 6256 74012
rect 5960 73958 6006 74010
rect 6006 73958 6016 74010
rect 6040 73958 6070 74010
rect 6070 73958 6082 74010
rect 6082 73958 6096 74010
rect 6120 73958 6134 74010
rect 6134 73958 6146 74010
rect 6146 73958 6176 74010
rect 6200 73958 6210 74010
rect 6210 73958 6256 74010
rect 5960 73956 6016 73958
rect 6040 73956 6096 73958
rect 6120 73956 6176 73958
rect 6200 73956 6256 73958
rect 7138 73856 7194 73912
rect 2906 73720 2962 73776
rect 6696 73466 6752 73468
rect 6776 73466 6832 73468
rect 6856 73466 6912 73468
rect 6936 73466 6992 73468
rect 6696 73414 6742 73466
rect 6742 73414 6752 73466
rect 6776 73414 6806 73466
rect 6806 73414 6818 73466
rect 6818 73414 6832 73466
rect 6856 73414 6870 73466
rect 6870 73414 6882 73466
rect 6882 73414 6912 73466
rect 6936 73414 6946 73466
rect 6946 73414 6992 73466
rect 6696 73412 6752 73414
rect 6776 73412 6832 73414
rect 6856 73412 6912 73414
rect 6936 73412 6992 73414
rect 2906 73060 2962 73096
rect 2906 73040 2908 73060
rect 2908 73040 2960 73060
rect 2960 73040 2962 73060
rect 5960 72922 6016 72924
rect 6040 72922 6096 72924
rect 6120 72922 6176 72924
rect 6200 72922 6256 72924
rect 5960 72870 6006 72922
rect 6006 72870 6016 72922
rect 6040 72870 6070 72922
rect 6070 72870 6082 72922
rect 6082 72870 6096 72922
rect 6120 72870 6134 72922
rect 6134 72870 6146 72922
rect 6146 72870 6176 72922
rect 6200 72870 6210 72922
rect 6210 72870 6256 72922
rect 5960 72868 6016 72870
rect 6040 72868 6096 72870
rect 6120 72868 6176 72870
rect 6200 72868 6256 72870
rect 7138 72768 7194 72824
rect 6696 72378 6752 72380
rect 6776 72378 6832 72380
rect 6856 72378 6912 72380
rect 6936 72378 6992 72380
rect 6696 72326 6742 72378
rect 6742 72326 6752 72378
rect 6776 72326 6806 72378
rect 6806 72326 6818 72378
rect 6818 72326 6832 72378
rect 6856 72326 6870 72378
rect 6870 72326 6882 72378
rect 6882 72326 6912 72378
rect 6936 72326 6946 72378
rect 6946 72326 6992 72378
rect 6696 72324 6752 72326
rect 6776 72324 6832 72326
rect 6856 72324 6912 72326
rect 6936 72324 6992 72326
rect 4378 71680 4434 71736
rect 5960 71834 6016 71836
rect 6040 71834 6096 71836
rect 6120 71834 6176 71836
rect 6200 71834 6256 71836
rect 5960 71782 6006 71834
rect 6006 71782 6016 71834
rect 6040 71782 6070 71834
rect 6070 71782 6082 71834
rect 6082 71782 6096 71834
rect 6120 71782 6134 71834
rect 6134 71782 6146 71834
rect 6146 71782 6176 71834
rect 6200 71782 6210 71834
rect 6210 71782 6256 71834
rect 5960 71780 6016 71782
rect 6040 71780 6096 71782
rect 6120 71780 6176 71782
rect 6200 71780 6256 71782
rect 5666 71544 5722 71600
rect 6696 71290 6752 71292
rect 6776 71290 6832 71292
rect 6856 71290 6912 71292
rect 6936 71290 6992 71292
rect 6696 71238 6742 71290
rect 6742 71238 6752 71290
rect 6776 71238 6806 71290
rect 6806 71238 6818 71290
rect 6818 71238 6832 71290
rect 6856 71238 6870 71290
rect 6870 71238 6882 71290
rect 6882 71238 6912 71290
rect 6936 71238 6946 71290
rect 6946 71238 6992 71290
rect 6696 71236 6752 71238
rect 6776 71236 6832 71238
rect 6856 71236 6912 71238
rect 6936 71236 6992 71238
rect 5666 70864 5722 70920
rect 5960 70746 6016 70748
rect 6040 70746 6096 70748
rect 6120 70746 6176 70748
rect 6200 70746 6256 70748
rect 5960 70694 6006 70746
rect 6006 70694 6016 70746
rect 6040 70694 6070 70746
rect 6070 70694 6082 70746
rect 6082 70694 6096 70746
rect 6120 70694 6134 70746
rect 6134 70694 6146 70746
rect 6146 70694 6176 70746
rect 6200 70694 6210 70746
rect 6210 70694 6256 70746
rect 5960 70692 6016 70694
rect 6040 70692 6096 70694
rect 6120 70692 6176 70694
rect 6200 70692 6256 70694
rect 2906 70340 2962 70376
rect 2906 70320 2908 70340
rect 2908 70320 2960 70340
rect 2960 70320 2962 70340
rect 6696 70202 6752 70204
rect 6776 70202 6832 70204
rect 6856 70202 6912 70204
rect 6936 70202 6992 70204
rect 6696 70150 6742 70202
rect 6742 70150 6752 70202
rect 6776 70150 6806 70202
rect 6806 70150 6818 70202
rect 6818 70150 6832 70202
rect 6856 70150 6870 70202
rect 6870 70150 6882 70202
rect 6882 70150 6912 70202
rect 6936 70150 6946 70202
rect 6946 70150 6992 70202
rect 6696 70148 6752 70150
rect 6776 70148 6832 70150
rect 6856 70148 6912 70150
rect 6936 70148 6992 70150
rect 2906 69640 2962 69696
rect 5960 69658 6016 69660
rect 6040 69658 6096 69660
rect 6120 69658 6176 69660
rect 6200 69658 6256 69660
rect 5960 69606 6006 69658
rect 6006 69606 6016 69658
rect 6040 69606 6070 69658
rect 6070 69606 6082 69658
rect 6082 69606 6096 69658
rect 6120 69606 6134 69658
rect 6134 69606 6146 69658
rect 6146 69606 6176 69658
rect 6200 69606 6210 69658
rect 6210 69606 6256 69658
rect 5960 69604 6016 69606
rect 6040 69604 6096 69606
rect 6120 69604 6176 69606
rect 6200 69604 6256 69606
rect 7138 69504 7194 69560
rect 6696 69114 6752 69116
rect 6776 69114 6832 69116
rect 6856 69114 6912 69116
rect 6936 69114 6992 69116
rect 6696 69062 6742 69114
rect 6742 69062 6752 69114
rect 6776 69062 6806 69114
rect 6806 69062 6818 69114
rect 6818 69062 6832 69114
rect 6856 69062 6870 69114
rect 6870 69062 6882 69114
rect 6882 69062 6912 69114
rect 6936 69062 6946 69114
rect 6946 69062 6992 69114
rect 6696 69060 6752 69062
rect 6776 69060 6832 69062
rect 6856 69060 6912 69062
rect 6936 69060 6992 69062
rect 5960 68570 6016 68572
rect 6040 68570 6096 68572
rect 6120 68570 6176 68572
rect 6200 68570 6256 68572
rect 5960 68518 6006 68570
rect 6006 68518 6016 68570
rect 6040 68518 6070 68570
rect 6070 68518 6082 68570
rect 6082 68518 6096 68570
rect 6120 68518 6134 68570
rect 6134 68518 6146 68570
rect 6146 68518 6176 68570
rect 6200 68518 6210 68570
rect 6210 68518 6256 68570
rect 5960 68516 6016 68518
rect 6040 68516 6096 68518
rect 6120 68516 6176 68518
rect 6200 68516 6256 68518
rect 7138 68416 7194 68472
rect 2906 68280 2962 68336
rect 6696 68026 6752 68028
rect 6776 68026 6832 68028
rect 6856 68026 6912 68028
rect 6936 68026 6992 68028
rect 6696 67974 6742 68026
rect 6742 67974 6752 68026
rect 6776 67974 6806 68026
rect 6806 67974 6818 68026
rect 6818 67974 6832 68026
rect 6856 67974 6870 68026
rect 6870 67974 6882 68026
rect 6882 67974 6912 68026
rect 6936 67974 6946 68026
rect 6946 67974 6992 68026
rect 6696 67972 6752 67974
rect 6776 67972 6832 67974
rect 6856 67972 6912 67974
rect 6936 67972 6992 67974
rect 2906 67620 2962 67656
rect 2906 67600 2908 67620
rect 2908 67600 2960 67620
rect 2960 67600 2962 67620
rect 5960 67482 6016 67484
rect 6040 67482 6096 67484
rect 6120 67482 6176 67484
rect 6200 67482 6256 67484
rect 5960 67430 6006 67482
rect 6006 67430 6016 67482
rect 6040 67430 6070 67482
rect 6070 67430 6082 67482
rect 6082 67430 6096 67482
rect 6120 67430 6134 67482
rect 6134 67430 6146 67482
rect 6146 67430 6176 67482
rect 6200 67430 6210 67482
rect 6210 67430 6256 67482
rect 5960 67428 6016 67430
rect 6040 67428 6096 67430
rect 6120 67428 6176 67430
rect 6200 67428 6256 67430
rect 7138 67328 7194 67384
rect 6696 66938 6752 66940
rect 6776 66938 6832 66940
rect 6856 66938 6912 66940
rect 6936 66938 6992 66940
rect 6696 66886 6742 66938
rect 6742 66886 6752 66938
rect 6776 66886 6806 66938
rect 6806 66886 6818 66938
rect 6818 66886 6832 66938
rect 6856 66886 6870 66938
rect 6870 66886 6882 66938
rect 6882 66886 6912 66938
rect 6936 66886 6946 66938
rect 6946 66886 6992 66938
rect 6696 66884 6752 66886
rect 6776 66884 6832 66886
rect 6856 66884 6912 66886
rect 6936 66884 6992 66886
rect 4378 66240 4434 66296
rect 5960 66394 6016 66396
rect 6040 66394 6096 66396
rect 6120 66394 6176 66396
rect 6200 66394 6256 66396
rect 5960 66342 6006 66394
rect 6006 66342 6016 66394
rect 6040 66342 6070 66394
rect 6070 66342 6082 66394
rect 6082 66342 6096 66394
rect 6120 66342 6134 66394
rect 6134 66342 6146 66394
rect 6146 66342 6176 66394
rect 6200 66342 6210 66394
rect 6210 66342 6256 66394
rect 5960 66340 6016 66342
rect 6040 66340 6096 66342
rect 6120 66340 6176 66342
rect 6200 66340 6256 66342
rect 5482 66104 5538 66160
rect 6696 65850 6752 65852
rect 6776 65850 6832 65852
rect 6856 65850 6912 65852
rect 6936 65850 6992 65852
rect 6696 65798 6742 65850
rect 6742 65798 6752 65850
rect 6776 65798 6806 65850
rect 6806 65798 6818 65850
rect 6818 65798 6832 65850
rect 6856 65798 6870 65850
rect 6870 65798 6882 65850
rect 6882 65798 6912 65850
rect 6936 65798 6946 65850
rect 6946 65798 6992 65850
rect 6696 65796 6752 65798
rect 6776 65796 6832 65798
rect 6856 65796 6912 65798
rect 6936 65796 6992 65798
rect 5390 65424 5446 65480
rect 5960 65306 6016 65308
rect 6040 65306 6096 65308
rect 6120 65306 6176 65308
rect 6200 65306 6256 65308
rect 5960 65254 6006 65306
rect 6006 65254 6016 65306
rect 6040 65254 6070 65306
rect 6070 65254 6082 65306
rect 6082 65254 6096 65306
rect 6120 65254 6134 65306
rect 6134 65254 6146 65306
rect 6146 65254 6176 65306
rect 6200 65254 6210 65306
rect 6210 65254 6256 65306
rect 5960 65252 6016 65254
rect 6040 65252 6096 65254
rect 6120 65252 6176 65254
rect 6200 65252 6256 65254
rect 2906 64916 2908 64936
rect 2908 64916 2960 64936
rect 2960 64916 2962 64936
rect 2906 64880 2962 64916
rect 6696 64762 6752 64764
rect 6776 64762 6832 64764
rect 6856 64762 6912 64764
rect 6936 64762 6992 64764
rect 6696 64710 6742 64762
rect 6742 64710 6752 64762
rect 6776 64710 6806 64762
rect 6806 64710 6818 64762
rect 6818 64710 6832 64762
rect 6856 64710 6870 64762
rect 6870 64710 6882 64762
rect 6882 64710 6912 64762
rect 6936 64710 6946 64762
rect 6946 64710 6992 64762
rect 6696 64708 6752 64710
rect 6776 64708 6832 64710
rect 6856 64708 6912 64710
rect 6936 64708 6992 64710
rect 2906 64200 2962 64256
rect 5960 64218 6016 64220
rect 6040 64218 6096 64220
rect 6120 64218 6176 64220
rect 6200 64218 6256 64220
rect 5960 64166 6006 64218
rect 6006 64166 6016 64218
rect 6040 64166 6070 64218
rect 6070 64166 6082 64218
rect 6082 64166 6096 64218
rect 6120 64166 6134 64218
rect 6134 64166 6146 64218
rect 6146 64166 6176 64218
rect 6200 64166 6210 64218
rect 6210 64166 6256 64218
rect 5960 64164 6016 64166
rect 6040 64164 6096 64166
rect 6120 64164 6176 64166
rect 6200 64164 6256 64166
rect 7230 64064 7286 64120
rect 6696 63674 6752 63676
rect 6776 63674 6832 63676
rect 6856 63674 6912 63676
rect 6936 63674 6992 63676
rect 6696 63622 6742 63674
rect 6742 63622 6752 63674
rect 6776 63622 6806 63674
rect 6806 63622 6818 63674
rect 6818 63622 6832 63674
rect 6856 63622 6870 63674
rect 6870 63622 6882 63674
rect 6882 63622 6912 63674
rect 6936 63622 6946 63674
rect 6946 63622 6992 63674
rect 6696 63620 6752 63622
rect 6776 63620 6832 63622
rect 6856 63620 6912 63622
rect 6936 63620 6992 63622
rect 5960 63130 6016 63132
rect 6040 63130 6096 63132
rect 6120 63130 6176 63132
rect 6200 63130 6256 63132
rect 5960 63078 6006 63130
rect 6006 63078 6016 63130
rect 6040 63078 6070 63130
rect 6070 63078 6082 63130
rect 6082 63078 6096 63130
rect 6120 63078 6134 63130
rect 6134 63078 6146 63130
rect 6146 63078 6176 63130
rect 6200 63078 6210 63130
rect 6210 63078 6256 63130
rect 5960 63076 6016 63078
rect 6040 63076 6096 63078
rect 6120 63076 6176 63078
rect 6200 63076 6256 63078
rect 7230 62976 7286 63032
rect 2906 62840 2962 62896
rect 6696 62586 6752 62588
rect 6776 62586 6832 62588
rect 6856 62586 6912 62588
rect 6936 62586 6992 62588
rect 6696 62534 6742 62586
rect 6742 62534 6752 62586
rect 6776 62534 6806 62586
rect 6806 62534 6818 62586
rect 6818 62534 6832 62586
rect 6856 62534 6870 62586
rect 6870 62534 6882 62586
rect 6882 62534 6912 62586
rect 6936 62534 6946 62586
rect 6946 62534 6992 62586
rect 6696 62532 6752 62534
rect 6776 62532 6832 62534
rect 6856 62532 6912 62534
rect 6936 62532 6992 62534
rect 5206 62160 5262 62216
rect 5960 62042 6016 62044
rect 6040 62042 6096 62044
rect 6120 62042 6176 62044
rect 6200 62042 6256 62044
rect 5960 61990 6006 62042
rect 6006 61990 6016 62042
rect 6040 61990 6070 62042
rect 6070 61990 6082 62042
rect 6082 61990 6096 62042
rect 6120 61990 6134 62042
rect 6134 61990 6146 62042
rect 6146 61990 6176 62042
rect 6200 61990 6210 62042
rect 6210 61990 6256 62042
rect 5960 61988 6016 61990
rect 6040 61988 6096 61990
rect 6120 61988 6176 61990
rect 6200 61988 6256 61990
rect 6696 61498 6752 61500
rect 6776 61498 6832 61500
rect 6856 61498 6912 61500
rect 6936 61498 6992 61500
rect 6696 61446 6742 61498
rect 6742 61446 6752 61498
rect 6776 61446 6806 61498
rect 6806 61446 6818 61498
rect 6818 61446 6832 61498
rect 6856 61446 6870 61498
rect 6870 61446 6882 61498
rect 6882 61446 6912 61498
rect 6936 61446 6946 61498
rect 6946 61446 6992 61498
rect 6696 61444 6752 61446
rect 6776 61444 6832 61446
rect 6856 61444 6912 61446
rect 6936 61444 6992 61446
rect 5960 60954 6016 60956
rect 6040 60954 6096 60956
rect 6120 60954 6176 60956
rect 6200 60954 6256 60956
rect 5960 60902 6006 60954
rect 6006 60902 6016 60954
rect 6040 60902 6070 60954
rect 6070 60902 6082 60954
rect 6082 60902 6096 60954
rect 6120 60902 6134 60954
rect 6134 60902 6146 60954
rect 6146 60902 6176 60954
rect 6200 60902 6210 60954
rect 6210 60902 6256 60954
rect 5960 60900 6016 60902
rect 6040 60900 6096 60902
rect 6120 60900 6176 60902
rect 6200 60900 6256 60902
rect 5206 60800 5262 60856
rect 6696 60410 6752 60412
rect 6776 60410 6832 60412
rect 6856 60410 6912 60412
rect 6936 60410 6992 60412
rect 6696 60358 6742 60410
rect 6742 60358 6752 60410
rect 6776 60358 6806 60410
rect 6806 60358 6818 60410
rect 6818 60358 6832 60410
rect 6856 60358 6870 60410
rect 6870 60358 6882 60410
rect 6882 60358 6912 60410
rect 6936 60358 6946 60410
rect 6946 60358 6992 60410
rect 6696 60356 6752 60358
rect 6776 60356 6832 60358
rect 6856 60356 6912 60358
rect 6936 60356 6992 60358
rect 5960 59866 6016 59868
rect 6040 59866 6096 59868
rect 6120 59866 6176 59868
rect 6200 59866 6256 59868
rect 5960 59814 6006 59866
rect 6006 59814 6016 59866
rect 6040 59814 6070 59866
rect 6070 59814 6082 59866
rect 6082 59814 6096 59866
rect 6120 59814 6134 59866
rect 6134 59814 6146 59866
rect 6146 59814 6176 59866
rect 6200 59814 6210 59866
rect 6210 59814 6256 59866
rect 5960 59812 6016 59814
rect 6040 59812 6096 59814
rect 6120 59812 6176 59814
rect 6200 59812 6256 59814
rect 5666 59576 5722 59632
rect 2906 59476 2908 59496
rect 2908 59476 2960 59496
rect 2960 59476 2962 59496
rect 2906 59440 2962 59476
rect 6696 59322 6752 59324
rect 6776 59322 6832 59324
rect 6856 59322 6912 59324
rect 6936 59322 6992 59324
rect 6696 59270 6742 59322
rect 6742 59270 6752 59322
rect 6776 59270 6806 59322
rect 6806 59270 6818 59322
rect 6818 59270 6832 59322
rect 6856 59270 6870 59322
rect 6870 59270 6882 59322
rect 6882 59270 6912 59322
rect 6936 59270 6946 59322
rect 6946 59270 6992 59322
rect 6696 59268 6752 59270
rect 6776 59268 6832 59270
rect 6856 59268 6912 59270
rect 6936 59268 6992 59270
rect 2906 58760 2962 58816
rect 5960 58778 6016 58780
rect 6040 58778 6096 58780
rect 6120 58778 6176 58780
rect 6200 58778 6256 58780
rect 5960 58726 6006 58778
rect 6006 58726 6016 58778
rect 6040 58726 6070 58778
rect 6070 58726 6082 58778
rect 6082 58726 6096 58778
rect 6120 58726 6134 58778
rect 6134 58726 6146 58778
rect 6146 58726 6176 58778
rect 6200 58726 6210 58778
rect 6210 58726 6256 58778
rect 5960 58724 6016 58726
rect 6040 58724 6096 58726
rect 6120 58724 6176 58726
rect 6200 58724 6256 58726
rect 7230 58624 7286 58680
rect 6696 58234 6752 58236
rect 6776 58234 6832 58236
rect 6856 58234 6912 58236
rect 6936 58234 6992 58236
rect 6696 58182 6742 58234
rect 6742 58182 6752 58234
rect 6776 58182 6806 58234
rect 6806 58182 6818 58234
rect 6818 58182 6832 58234
rect 6856 58182 6870 58234
rect 6870 58182 6882 58234
rect 6882 58182 6912 58234
rect 6936 58182 6946 58234
rect 6946 58182 6992 58234
rect 6696 58180 6752 58182
rect 6776 58180 6832 58182
rect 6856 58180 6912 58182
rect 6936 58180 6992 58182
rect 5960 57690 6016 57692
rect 6040 57690 6096 57692
rect 6120 57690 6176 57692
rect 6200 57690 6256 57692
rect 5960 57638 6006 57690
rect 6006 57638 6016 57690
rect 6040 57638 6070 57690
rect 6070 57638 6082 57690
rect 6082 57638 6096 57690
rect 6120 57638 6134 57690
rect 6134 57638 6146 57690
rect 6146 57638 6176 57690
rect 6200 57638 6210 57690
rect 6210 57638 6256 57690
rect 5960 57636 6016 57638
rect 6040 57636 6096 57638
rect 6120 57636 6176 57638
rect 6200 57636 6256 57638
rect 7230 57536 7286 57592
rect 2906 57400 2962 57456
rect 6696 57146 6752 57148
rect 6776 57146 6832 57148
rect 6856 57146 6912 57148
rect 6936 57146 6992 57148
rect 6696 57094 6742 57146
rect 6742 57094 6752 57146
rect 6776 57094 6806 57146
rect 6806 57094 6818 57146
rect 6818 57094 6832 57146
rect 6856 57094 6870 57146
rect 6870 57094 6882 57146
rect 6882 57094 6912 57146
rect 6936 57094 6946 57146
rect 6946 57094 6992 57146
rect 6696 57092 6752 57094
rect 6776 57092 6832 57094
rect 6856 57092 6912 57094
rect 6936 57092 6992 57094
rect 4930 56720 4986 56776
rect 5960 56602 6016 56604
rect 6040 56602 6096 56604
rect 6120 56602 6176 56604
rect 6200 56602 6256 56604
rect 5960 56550 6006 56602
rect 6006 56550 6016 56602
rect 6040 56550 6070 56602
rect 6070 56550 6082 56602
rect 6082 56550 6096 56602
rect 6120 56550 6134 56602
rect 6134 56550 6146 56602
rect 6146 56550 6176 56602
rect 6200 56550 6210 56602
rect 6210 56550 6256 56602
rect 5960 56548 6016 56550
rect 6040 56548 6096 56550
rect 6120 56548 6176 56550
rect 6200 56548 6256 56550
rect 5390 56312 5446 56368
rect 6696 56058 6752 56060
rect 6776 56058 6832 56060
rect 6856 56058 6912 56060
rect 6936 56058 6992 56060
rect 6696 56006 6742 56058
rect 6742 56006 6752 56058
rect 6776 56006 6806 56058
rect 6806 56006 6818 56058
rect 6818 56006 6832 56058
rect 6856 56006 6870 56058
rect 6870 56006 6882 56058
rect 6882 56006 6912 56058
rect 6936 56006 6946 56058
rect 6946 56006 6992 56058
rect 6696 56004 6752 56006
rect 6776 56004 6832 56006
rect 6856 56004 6912 56006
rect 6936 56004 6992 56006
rect 5022 55360 5078 55416
rect 5960 55514 6016 55516
rect 6040 55514 6096 55516
rect 6120 55514 6176 55516
rect 6200 55514 6256 55516
rect 5960 55462 6006 55514
rect 6006 55462 6016 55514
rect 6040 55462 6070 55514
rect 6070 55462 6082 55514
rect 6082 55462 6096 55514
rect 6120 55462 6134 55514
rect 6134 55462 6146 55514
rect 6146 55462 6176 55514
rect 6200 55462 6210 55514
rect 6210 55462 6256 55514
rect 5960 55460 6016 55462
rect 6040 55460 6096 55462
rect 6120 55460 6176 55462
rect 6200 55460 6256 55462
rect 5666 55224 5722 55280
rect 6696 54970 6752 54972
rect 6776 54970 6832 54972
rect 6856 54970 6912 54972
rect 6936 54970 6992 54972
rect 6696 54918 6742 54970
rect 6742 54918 6752 54970
rect 6776 54918 6806 54970
rect 6806 54918 6818 54970
rect 6818 54918 6832 54970
rect 6856 54918 6870 54970
rect 6870 54918 6882 54970
rect 6882 54918 6912 54970
rect 6936 54918 6946 54970
rect 6946 54918 6992 54970
rect 6696 54916 6752 54918
rect 6776 54916 6832 54918
rect 6856 54916 6912 54918
rect 6936 54916 6992 54918
rect 8426 84328 8482 84384
rect 14406 84328 14462 84384
rect 19388 88698 19444 88700
rect 19468 88698 19524 88700
rect 19548 88698 19604 88700
rect 19628 88698 19684 88700
rect 19388 88646 19434 88698
rect 19434 88646 19444 88698
rect 19468 88646 19498 88698
rect 19498 88646 19510 88698
rect 19510 88646 19524 88698
rect 19548 88646 19562 88698
rect 19562 88646 19574 88698
rect 19574 88646 19604 88698
rect 19628 88646 19638 88698
rect 19638 88646 19684 88698
rect 19388 88644 19444 88646
rect 19468 88644 19524 88646
rect 19548 88644 19604 88646
rect 19628 88644 19684 88646
rect 18728 88154 18784 88156
rect 18808 88154 18864 88156
rect 18888 88154 18944 88156
rect 18968 88154 19024 88156
rect 18728 88102 18774 88154
rect 18774 88102 18784 88154
rect 18808 88102 18838 88154
rect 18838 88102 18850 88154
rect 18850 88102 18864 88154
rect 18888 88102 18902 88154
rect 18902 88102 18914 88154
rect 18914 88102 18944 88154
rect 18968 88102 18978 88154
rect 18978 88102 19024 88154
rect 18728 88100 18784 88102
rect 18808 88100 18864 88102
rect 18888 88100 18944 88102
rect 18968 88100 19024 88102
rect 19388 87610 19444 87612
rect 19468 87610 19524 87612
rect 19548 87610 19604 87612
rect 19628 87610 19684 87612
rect 19388 87558 19434 87610
rect 19434 87558 19444 87610
rect 19468 87558 19498 87610
rect 19498 87558 19510 87610
rect 19510 87558 19524 87610
rect 19548 87558 19562 87610
rect 19562 87558 19574 87610
rect 19574 87558 19604 87610
rect 19628 87558 19638 87610
rect 19638 87558 19684 87610
rect 19388 87556 19444 87558
rect 19468 87556 19524 87558
rect 19548 87556 19604 87558
rect 19628 87556 19684 87558
rect 18728 87066 18784 87068
rect 18808 87066 18864 87068
rect 18888 87066 18944 87068
rect 18968 87066 19024 87068
rect 18728 87014 18774 87066
rect 18774 87014 18784 87066
rect 18808 87014 18838 87066
rect 18838 87014 18850 87066
rect 18850 87014 18864 87066
rect 18888 87014 18902 87066
rect 18902 87014 18914 87066
rect 18914 87014 18944 87066
rect 18968 87014 18978 87066
rect 18978 87014 19024 87066
rect 18728 87012 18784 87014
rect 18808 87012 18864 87014
rect 18888 87012 18944 87014
rect 18968 87012 19024 87014
rect 19388 86522 19444 86524
rect 19468 86522 19524 86524
rect 19548 86522 19604 86524
rect 19628 86522 19684 86524
rect 19388 86470 19434 86522
rect 19434 86470 19444 86522
rect 19468 86470 19498 86522
rect 19498 86470 19510 86522
rect 19510 86470 19524 86522
rect 19548 86470 19562 86522
rect 19562 86470 19574 86522
rect 19574 86470 19604 86522
rect 19628 86470 19638 86522
rect 19638 86470 19684 86522
rect 19388 86468 19444 86470
rect 19468 86468 19524 86470
rect 19548 86468 19604 86470
rect 19628 86468 19684 86470
rect 2538 54680 2594 54736
rect 5960 54426 6016 54428
rect 6040 54426 6096 54428
rect 6120 54426 6176 54428
rect 6200 54426 6256 54428
rect 5960 54374 6006 54426
rect 6006 54374 6016 54426
rect 6040 54374 6070 54426
rect 6070 54374 6082 54426
rect 6082 54374 6096 54426
rect 6120 54374 6134 54426
rect 6134 54374 6146 54426
rect 6146 54374 6176 54426
rect 6200 54374 6210 54426
rect 6210 54374 6256 54426
rect 5960 54372 6016 54374
rect 6040 54372 6096 54374
rect 6120 54372 6176 54374
rect 6200 54372 6256 54374
rect 5666 54136 5722 54192
rect 5206 54036 5208 54056
rect 5208 54036 5260 54056
rect 5260 54036 5262 54056
rect 5206 54000 5262 54036
rect 6696 53882 6752 53884
rect 6776 53882 6832 53884
rect 6856 53882 6912 53884
rect 6936 53882 6992 53884
rect 6696 53830 6742 53882
rect 6742 53830 6752 53882
rect 6776 53830 6806 53882
rect 6806 53830 6818 53882
rect 6818 53830 6832 53882
rect 6856 53830 6870 53882
rect 6870 53830 6882 53882
rect 6882 53830 6912 53882
rect 6936 53830 6946 53882
rect 6946 53830 6992 53882
rect 6696 53828 6752 53830
rect 6776 53828 6832 53830
rect 6856 53828 6912 53830
rect 6936 53828 6992 53830
rect 2906 53320 2962 53376
rect 5960 53338 6016 53340
rect 6040 53338 6096 53340
rect 6120 53338 6176 53340
rect 6200 53338 6256 53340
rect 5960 53286 6006 53338
rect 6006 53286 6016 53338
rect 6040 53286 6070 53338
rect 6070 53286 6082 53338
rect 6082 53286 6096 53338
rect 6120 53286 6134 53338
rect 6134 53286 6146 53338
rect 6146 53286 6176 53338
rect 6200 53286 6210 53338
rect 6210 53286 6256 53338
rect 5960 53284 6016 53286
rect 6040 53284 6096 53286
rect 6120 53284 6176 53286
rect 6200 53284 6256 53286
rect 6696 52794 6752 52796
rect 6776 52794 6832 52796
rect 6856 52794 6912 52796
rect 6936 52794 6992 52796
rect 6696 52742 6742 52794
rect 6742 52742 6752 52794
rect 6776 52742 6806 52794
rect 6806 52742 6818 52794
rect 6818 52742 6832 52794
rect 6856 52742 6870 52794
rect 6870 52742 6882 52794
rect 6882 52742 6912 52794
rect 6936 52742 6946 52794
rect 6946 52742 6992 52794
rect 6696 52740 6752 52742
rect 6776 52740 6832 52742
rect 6856 52740 6912 52742
rect 6936 52740 6992 52742
rect 2906 52640 2962 52696
rect 5960 52250 6016 52252
rect 6040 52250 6096 52252
rect 6120 52250 6176 52252
rect 6200 52250 6256 52252
rect 5960 52198 6006 52250
rect 6006 52198 6016 52250
rect 6040 52198 6070 52250
rect 6070 52198 6082 52250
rect 6082 52198 6096 52250
rect 6120 52198 6134 52250
rect 6134 52198 6146 52250
rect 6146 52198 6176 52250
rect 6200 52198 6210 52250
rect 6210 52198 6256 52250
rect 5960 52196 6016 52198
rect 6040 52196 6096 52198
rect 6120 52196 6176 52198
rect 6200 52196 6256 52198
rect 2906 51960 2962 52016
rect 6696 51706 6752 51708
rect 6776 51706 6832 51708
rect 6856 51706 6912 51708
rect 6936 51706 6992 51708
rect 6696 51654 6742 51706
rect 6742 51654 6752 51706
rect 6776 51654 6806 51706
rect 6806 51654 6818 51706
rect 6818 51654 6832 51706
rect 6856 51654 6870 51706
rect 6870 51654 6882 51706
rect 6882 51654 6912 51706
rect 6936 51654 6946 51706
rect 6946 51654 6992 51706
rect 6696 51652 6752 51654
rect 6776 51652 6832 51654
rect 6856 51652 6912 51654
rect 6936 51652 6992 51654
rect 2906 51280 2962 51336
rect 5960 51162 6016 51164
rect 6040 51162 6096 51164
rect 6120 51162 6176 51164
rect 6200 51162 6256 51164
rect 5960 51110 6006 51162
rect 6006 51110 6016 51162
rect 6040 51110 6070 51162
rect 6070 51110 6082 51162
rect 6082 51110 6096 51162
rect 6120 51110 6134 51162
rect 6134 51110 6146 51162
rect 6146 51110 6176 51162
rect 6200 51110 6210 51162
rect 6210 51110 6256 51162
rect 5960 51108 6016 51110
rect 6040 51108 6096 51110
rect 6120 51108 6176 51110
rect 6200 51108 6256 51110
rect 5666 50872 5722 50928
rect 6696 50618 6752 50620
rect 6776 50618 6832 50620
rect 6856 50618 6912 50620
rect 6936 50618 6992 50620
rect 6696 50566 6742 50618
rect 6742 50566 6752 50618
rect 6776 50566 6806 50618
rect 6806 50566 6818 50618
rect 6818 50566 6832 50618
rect 6856 50566 6870 50618
rect 6870 50566 6882 50618
rect 6882 50566 6912 50618
rect 6936 50566 6946 50618
rect 6946 50566 6992 50618
rect 6696 50564 6752 50566
rect 6776 50564 6832 50566
rect 6856 50564 6912 50566
rect 6936 50564 6992 50566
rect 5960 50074 6016 50076
rect 6040 50074 6096 50076
rect 6120 50074 6176 50076
rect 6200 50074 6256 50076
rect 5960 50022 6006 50074
rect 6006 50022 6016 50074
rect 6040 50022 6070 50074
rect 6070 50022 6082 50074
rect 6082 50022 6096 50074
rect 6120 50022 6134 50074
rect 6134 50022 6146 50074
rect 6146 50022 6176 50074
rect 6200 50022 6210 50074
rect 6210 50022 6256 50074
rect 5960 50020 6016 50022
rect 6040 50020 6096 50022
rect 6120 50020 6176 50022
rect 6200 50020 6256 50022
rect 6696 49530 6752 49532
rect 6776 49530 6832 49532
rect 6856 49530 6912 49532
rect 6936 49530 6992 49532
rect 6696 49478 6742 49530
rect 6742 49478 6752 49530
rect 6776 49478 6806 49530
rect 6806 49478 6818 49530
rect 6818 49478 6832 49530
rect 6856 49478 6870 49530
rect 6870 49478 6882 49530
rect 6882 49478 6912 49530
rect 6936 49478 6946 49530
rect 6946 49478 6992 49530
rect 6696 49476 6752 49478
rect 6776 49476 6832 49478
rect 6856 49476 6912 49478
rect 6936 49476 6992 49478
rect 2906 49240 2962 49296
rect 5960 48986 6016 48988
rect 6040 48986 6096 48988
rect 6120 48986 6176 48988
rect 6200 48986 6256 48988
rect 5960 48934 6006 48986
rect 6006 48934 6016 48986
rect 6040 48934 6070 48986
rect 6070 48934 6082 48986
rect 6082 48934 6096 48986
rect 6120 48934 6134 48986
rect 6134 48934 6146 48986
rect 6146 48934 6176 48986
rect 6200 48934 6210 48986
rect 6210 48934 6256 48986
rect 5960 48932 6016 48934
rect 6040 48932 6096 48934
rect 6120 48932 6176 48934
rect 6200 48932 6256 48934
rect 6696 48442 6752 48444
rect 6776 48442 6832 48444
rect 6856 48442 6912 48444
rect 6936 48442 6992 48444
rect 6696 48390 6742 48442
rect 6742 48390 6752 48442
rect 6776 48390 6806 48442
rect 6806 48390 6818 48442
rect 6818 48390 6832 48442
rect 6856 48390 6870 48442
rect 6870 48390 6882 48442
rect 6882 48390 6912 48442
rect 6936 48390 6946 48442
rect 6946 48390 6992 48442
rect 6696 48388 6752 48390
rect 6776 48388 6832 48390
rect 6856 48388 6912 48390
rect 6936 48388 6992 48390
rect 5960 47898 6016 47900
rect 6040 47898 6096 47900
rect 6120 47898 6176 47900
rect 6200 47898 6256 47900
rect 5960 47846 6006 47898
rect 6006 47846 6016 47898
rect 6040 47846 6070 47898
rect 6070 47846 6082 47898
rect 6082 47846 6096 47898
rect 6120 47846 6134 47898
rect 6134 47846 6146 47898
rect 6146 47846 6176 47898
rect 6200 47846 6210 47898
rect 6210 47846 6256 47898
rect 5960 47844 6016 47846
rect 6040 47844 6096 47846
rect 6120 47844 6176 47846
rect 6200 47844 6256 47846
rect 6696 47354 6752 47356
rect 6776 47354 6832 47356
rect 6856 47354 6912 47356
rect 6936 47354 6992 47356
rect 6696 47302 6742 47354
rect 6742 47302 6752 47354
rect 6776 47302 6806 47354
rect 6806 47302 6818 47354
rect 6818 47302 6832 47354
rect 6856 47302 6870 47354
rect 6870 47302 6882 47354
rect 6882 47302 6912 47354
rect 6936 47302 6946 47354
rect 6946 47302 6992 47354
rect 6696 47300 6752 47302
rect 6776 47300 6832 47302
rect 6856 47300 6912 47302
rect 6936 47300 6992 47302
rect 7138 53204 7194 53240
rect 7138 53184 7140 53204
rect 7140 53184 7192 53204
rect 7192 53184 7194 53204
rect 7138 52096 7194 52152
rect 5960 46810 6016 46812
rect 6040 46810 6096 46812
rect 6120 46810 6176 46812
rect 6200 46810 6256 46812
rect 5960 46758 6006 46810
rect 6006 46758 6016 46810
rect 6040 46758 6070 46810
rect 6070 46758 6082 46810
rect 6082 46758 6096 46810
rect 6120 46758 6134 46810
rect 6134 46758 6146 46810
rect 6146 46758 6176 46810
rect 6200 46758 6210 46810
rect 6210 46758 6256 46810
rect 5960 46756 6016 46758
rect 6040 46756 6096 46758
rect 6120 46756 6176 46758
rect 6200 46756 6256 46758
rect 2906 46520 2962 46576
rect 6696 46266 6752 46268
rect 6776 46266 6832 46268
rect 6856 46266 6912 46268
rect 6936 46266 6992 46268
rect 6696 46214 6742 46266
rect 6742 46214 6752 46266
rect 6776 46214 6806 46266
rect 6806 46214 6818 46266
rect 6818 46214 6832 46266
rect 6856 46214 6870 46266
rect 6870 46214 6882 46266
rect 6882 46214 6912 46266
rect 6936 46214 6946 46266
rect 6946 46214 6992 46266
rect 6696 46212 6752 46214
rect 6776 46212 6832 46214
rect 6856 46212 6912 46214
rect 6936 46212 6992 46214
rect 2906 45860 2962 45896
rect 2906 45840 2908 45860
rect 2908 45840 2960 45860
rect 2960 45840 2962 45860
rect 5960 45722 6016 45724
rect 6040 45722 6096 45724
rect 6120 45722 6176 45724
rect 6200 45722 6256 45724
rect 5960 45670 6006 45722
rect 6006 45670 6016 45722
rect 6040 45670 6070 45722
rect 6070 45670 6082 45722
rect 6082 45670 6096 45722
rect 6120 45670 6134 45722
rect 6134 45670 6146 45722
rect 6146 45670 6176 45722
rect 6200 45670 6210 45722
rect 6210 45670 6256 45722
rect 5960 45668 6016 45670
rect 6040 45668 6096 45670
rect 6120 45668 6176 45670
rect 6200 45668 6256 45670
rect 6696 45178 6752 45180
rect 6776 45178 6832 45180
rect 6856 45178 6912 45180
rect 6936 45178 6992 45180
rect 6696 45126 6742 45178
rect 6742 45126 6752 45178
rect 6776 45126 6806 45178
rect 6806 45126 6818 45178
rect 6818 45126 6832 45178
rect 6856 45126 6870 45178
rect 6870 45126 6882 45178
rect 6882 45126 6912 45178
rect 6936 45126 6946 45178
rect 6946 45126 6992 45178
rect 6696 45124 6752 45126
rect 6776 45124 6832 45126
rect 6856 45124 6912 45126
rect 6936 45124 6992 45126
rect 5960 44634 6016 44636
rect 6040 44634 6096 44636
rect 6120 44634 6176 44636
rect 6200 44634 6256 44636
rect 5960 44582 6006 44634
rect 6006 44582 6016 44634
rect 6040 44582 6070 44634
rect 6070 44582 6082 44634
rect 6082 44582 6096 44634
rect 6120 44582 6134 44634
rect 6134 44582 6146 44634
rect 6146 44582 6176 44634
rect 6200 44582 6210 44634
rect 6210 44582 6256 44634
rect 5960 44580 6016 44582
rect 6040 44580 6096 44582
rect 6120 44580 6176 44582
rect 6200 44580 6256 44582
rect 2538 44480 2594 44536
rect 6696 44090 6752 44092
rect 6776 44090 6832 44092
rect 6856 44090 6912 44092
rect 6936 44090 6992 44092
rect 6696 44038 6742 44090
rect 6742 44038 6752 44090
rect 6776 44038 6806 44090
rect 6806 44038 6818 44090
rect 6818 44038 6832 44090
rect 6856 44038 6870 44090
rect 6870 44038 6882 44090
rect 6882 44038 6912 44090
rect 6936 44038 6946 44090
rect 6946 44038 6992 44090
rect 6696 44036 6752 44038
rect 6776 44036 6832 44038
rect 6856 44036 6912 44038
rect 6936 44036 6992 44038
rect 5206 43800 5262 43856
rect 5960 43546 6016 43548
rect 6040 43546 6096 43548
rect 6120 43546 6176 43548
rect 6200 43546 6256 43548
rect 5960 43494 6006 43546
rect 6006 43494 6016 43546
rect 6040 43494 6070 43546
rect 6070 43494 6082 43546
rect 6082 43494 6096 43546
rect 6120 43494 6134 43546
rect 6134 43494 6146 43546
rect 6146 43494 6176 43546
rect 6200 43494 6210 43546
rect 6210 43494 6256 43546
rect 5960 43492 6016 43494
rect 6040 43492 6096 43494
rect 6120 43492 6176 43494
rect 6200 43492 6256 43494
rect 2906 43140 2962 43176
rect 2906 43120 2908 43140
rect 2908 43120 2960 43140
rect 2960 43120 2962 43140
rect 6696 43002 6752 43004
rect 6776 43002 6832 43004
rect 6856 43002 6912 43004
rect 6936 43002 6992 43004
rect 6696 42950 6742 43002
rect 6742 42950 6752 43002
rect 6776 42950 6806 43002
rect 6806 42950 6818 43002
rect 6818 42950 6832 43002
rect 6856 42950 6870 43002
rect 6870 42950 6882 43002
rect 6882 42950 6912 43002
rect 6936 42950 6946 43002
rect 6946 42950 6992 43002
rect 7138 42984 7194 43040
rect 6696 42948 6752 42950
rect 6776 42948 6832 42950
rect 6856 42948 6912 42950
rect 6936 42948 6992 42950
rect 2906 42440 2962 42496
rect 5960 42458 6016 42460
rect 6040 42458 6096 42460
rect 6120 42458 6176 42460
rect 6200 42458 6256 42460
rect 5960 42406 6006 42458
rect 6006 42406 6016 42458
rect 6040 42406 6070 42458
rect 6070 42406 6082 42458
rect 6082 42406 6096 42458
rect 6120 42406 6134 42458
rect 6134 42406 6146 42458
rect 6146 42406 6176 42458
rect 6200 42406 6210 42458
rect 6210 42406 6256 42458
rect 5960 42404 6016 42406
rect 6040 42404 6096 42406
rect 6120 42404 6176 42406
rect 6200 42404 6256 42406
rect 6696 41914 6752 41916
rect 6776 41914 6832 41916
rect 6856 41914 6912 41916
rect 6936 41914 6992 41916
rect 6696 41862 6742 41914
rect 6742 41862 6752 41914
rect 6776 41862 6806 41914
rect 6806 41862 6818 41914
rect 6818 41862 6832 41914
rect 6856 41862 6870 41914
rect 6870 41862 6882 41914
rect 6882 41862 6912 41914
rect 6936 41862 6946 41914
rect 6946 41862 6992 41914
rect 7138 41896 7194 41952
rect 6696 41860 6752 41862
rect 6776 41860 6832 41862
rect 6856 41860 6912 41862
rect 6936 41860 6992 41862
rect 2906 41760 2962 41816
rect 4378 41080 4434 41136
rect 5960 41370 6016 41372
rect 6040 41370 6096 41372
rect 6120 41370 6176 41372
rect 6200 41370 6256 41372
rect 5960 41318 6006 41370
rect 6006 41318 6016 41370
rect 6040 41318 6070 41370
rect 6070 41318 6082 41370
rect 6082 41318 6096 41370
rect 6120 41318 6134 41370
rect 6134 41318 6146 41370
rect 6146 41318 6176 41370
rect 6200 41318 6210 41370
rect 6210 41318 6256 41370
rect 5960 41316 6016 41318
rect 6040 41316 6096 41318
rect 6120 41316 6176 41318
rect 6200 41316 6256 41318
rect 5666 40944 5722 41000
rect 6696 40826 6752 40828
rect 6776 40826 6832 40828
rect 6856 40826 6912 40828
rect 6936 40826 6992 40828
rect 6696 40774 6742 40826
rect 6742 40774 6752 40826
rect 6776 40774 6806 40826
rect 6806 40774 6818 40826
rect 6818 40774 6832 40826
rect 6856 40774 6870 40826
rect 6870 40774 6882 40826
rect 6882 40774 6912 40826
rect 6936 40774 6946 40826
rect 6946 40774 6992 40826
rect 6696 40772 6752 40774
rect 6776 40772 6832 40774
rect 6856 40772 6912 40774
rect 6936 40772 6992 40774
rect 5960 40282 6016 40284
rect 6040 40282 6096 40284
rect 6120 40282 6176 40284
rect 6200 40282 6256 40284
rect 5960 40230 6006 40282
rect 6006 40230 6016 40282
rect 6040 40230 6070 40282
rect 6070 40230 6082 40282
rect 6082 40230 6096 40282
rect 6120 40230 6134 40282
rect 6134 40230 6146 40282
rect 6146 40230 6176 40282
rect 6200 40230 6210 40282
rect 6210 40230 6256 40282
rect 5960 40228 6016 40230
rect 6040 40228 6096 40230
rect 6120 40228 6176 40230
rect 6200 40228 6256 40230
rect 2906 39720 2962 39776
rect 6696 39738 6752 39740
rect 6776 39738 6832 39740
rect 6856 39738 6912 39740
rect 6936 39738 6992 39740
rect 6696 39686 6742 39738
rect 6742 39686 6752 39738
rect 6776 39686 6806 39738
rect 6806 39686 6818 39738
rect 6818 39686 6832 39738
rect 6856 39686 6870 39738
rect 6870 39686 6882 39738
rect 6882 39686 6912 39738
rect 6936 39686 6946 39738
rect 6946 39686 6992 39738
rect 7138 39720 7194 39776
rect 6696 39684 6752 39686
rect 6776 39684 6832 39686
rect 6856 39684 6912 39686
rect 6936 39684 6992 39686
rect 5960 39194 6016 39196
rect 6040 39194 6096 39196
rect 6120 39194 6176 39196
rect 6200 39194 6256 39196
rect 5960 39142 6006 39194
rect 6006 39142 6016 39194
rect 6040 39142 6070 39194
rect 6070 39142 6082 39194
rect 6082 39142 6096 39194
rect 6120 39142 6134 39194
rect 6134 39142 6146 39194
rect 6146 39142 6176 39194
rect 6200 39142 6210 39194
rect 6210 39142 6256 39194
rect 5960 39140 6016 39142
rect 6040 39140 6096 39142
rect 6120 39140 6176 39142
rect 6200 39140 6256 39142
rect 6696 38650 6752 38652
rect 6776 38650 6832 38652
rect 6856 38650 6912 38652
rect 6936 38650 6992 38652
rect 6696 38598 6742 38650
rect 6742 38598 6752 38650
rect 6776 38598 6806 38650
rect 6806 38598 6818 38650
rect 6818 38598 6832 38650
rect 6856 38598 6870 38650
rect 6870 38598 6882 38650
rect 6882 38598 6912 38650
rect 6936 38598 6946 38650
rect 6946 38598 6992 38650
rect 7414 38632 7470 38688
rect 6696 38596 6752 38598
rect 6776 38596 6832 38598
rect 6856 38596 6912 38598
rect 6936 38596 6992 38598
rect 4378 38360 4434 38416
rect 5960 38106 6016 38108
rect 6040 38106 6096 38108
rect 6120 38106 6176 38108
rect 6200 38106 6256 38108
rect 5960 38054 6006 38106
rect 6006 38054 6016 38106
rect 6040 38054 6070 38106
rect 6070 38054 6082 38106
rect 6082 38054 6096 38106
rect 6120 38054 6134 38106
rect 6134 38054 6146 38106
rect 6146 38054 6176 38106
rect 6200 38054 6210 38106
rect 6210 38054 6256 38106
rect 5960 38052 6016 38054
rect 6040 38052 6096 38054
rect 6120 38052 6176 38054
rect 6200 38052 6256 38054
rect 2906 37700 2962 37736
rect 2906 37680 2908 37700
rect 2908 37680 2960 37700
rect 2960 37680 2962 37700
rect 6696 37562 6752 37564
rect 6776 37562 6832 37564
rect 6856 37562 6912 37564
rect 6936 37562 6992 37564
rect 6696 37510 6742 37562
rect 6742 37510 6752 37562
rect 6776 37510 6806 37562
rect 6806 37510 6818 37562
rect 6818 37510 6832 37562
rect 6856 37510 6870 37562
rect 6870 37510 6882 37562
rect 6882 37510 6912 37562
rect 6936 37510 6946 37562
rect 6946 37510 6992 37562
rect 7138 37544 7194 37600
rect 6696 37508 6752 37510
rect 6776 37508 6832 37510
rect 6856 37508 6912 37510
rect 6936 37508 6992 37510
rect 5960 37018 6016 37020
rect 6040 37018 6096 37020
rect 6120 37018 6176 37020
rect 6200 37018 6256 37020
rect 5960 36966 6006 37018
rect 6006 36966 6016 37018
rect 6040 36966 6070 37018
rect 6070 36966 6082 37018
rect 6082 36966 6096 37018
rect 6120 36966 6134 37018
rect 6134 36966 6146 37018
rect 6146 36966 6176 37018
rect 6200 36966 6210 37018
rect 6210 36966 6256 37018
rect 5960 36964 6016 36966
rect 6040 36964 6096 36966
rect 6120 36964 6176 36966
rect 6200 36964 6256 36966
rect 6696 36474 6752 36476
rect 6776 36474 6832 36476
rect 6856 36474 6912 36476
rect 6936 36474 6992 36476
rect 6696 36422 6742 36474
rect 6742 36422 6752 36474
rect 6776 36422 6806 36474
rect 6806 36422 6818 36474
rect 6818 36422 6832 36474
rect 6856 36422 6870 36474
rect 6870 36422 6882 36474
rect 6882 36422 6912 36474
rect 6936 36422 6946 36474
rect 6946 36422 6992 36474
rect 7138 36456 7194 36512
rect 6696 36420 6752 36422
rect 6776 36420 6832 36422
rect 6856 36420 6912 36422
rect 6936 36420 6992 36422
rect 2906 36320 2962 36376
rect 4378 35640 4434 35696
rect 5960 35930 6016 35932
rect 6040 35930 6096 35932
rect 6120 35930 6176 35932
rect 6200 35930 6256 35932
rect 5960 35878 6006 35930
rect 6006 35878 6016 35930
rect 6040 35878 6070 35930
rect 6070 35878 6082 35930
rect 6082 35878 6096 35930
rect 6120 35878 6134 35930
rect 6134 35878 6146 35930
rect 6146 35878 6176 35930
rect 6200 35878 6210 35930
rect 6210 35878 6256 35930
rect 5960 35876 6016 35878
rect 6040 35876 6096 35878
rect 6120 35876 6176 35878
rect 6200 35876 6256 35878
rect 5666 35504 5722 35560
rect 6696 35386 6752 35388
rect 6776 35386 6832 35388
rect 6856 35386 6912 35388
rect 6936 35386 6992 35388
rect 6696 35334 6742 35386
rect 6742 35334 6752 35386
rect 6776 35334 6806 35386
rect 6806 35334 6818 35386
rect 6818 35334 6832 35386
rect 6856 35334 6870 35386
rect 6870 35334 6882 35386
rect 6882 35334 6912 35386
rect 6936 35334 6946 35386
rect 6946 35334 6992 35386
rect 6696 35332 6752 35334
rect 6776 35332 6832 35334
rect 6856 35332 6912 35334
rect 6936 35332 6992 35334
rect 5960 34842 6016 34844
rect 6040 34842 6096 34844
rect 6120 34842 6176 34844
rect 6200 34842 6256 34844
rect 5960 34790 6006 34842
rect 6006 34790 6016 34842
rect 6040 34790 6070 34842
rect 6070 34790 6082 34842
rect 6082 34790 6096 34842
rect 6120 34790 6134 34842
rect 6134 34790 6146 34842
rect 6146 34790 6176 34842
rect 6200 34790 6210 34842
rect 6210 34790 6256 34842
rect 5960 34788 6016 34790
rect 6040 34788 6096 34790
rect 6120 34788 6176 34790
rect 6200 34788 6256 34790
rect 2906 34280 2962 34336
rect 6696 34298 6752 34300
rect 6776 34298 6832 34300
rect 6856 34298 6912 34300
rect 6936 34298 6992 34300
rect 6696 34246 6742 34298
rect 6742 34246 6752 34298
rect 6776 34246 6806 34298
rect 6806 34246 6818 34298
rect 6818 34246 6832 34298
rect 6856 34246 6870 34298
rect 6870 34246 6882 34298
rect 6882 34246 6912 34298
rect 6936 34246 6946 34298
rect 6946 34246 6992 34298
rect 7138 34280 7194 34336
rect 6696 34244 6752 34246
rect 6776 34244 6832 34246
rect 6856 34244 6912 34246
rect 6936 34244 6992 34246
rect 5960 33754 6016 33756
rect 6040 33754 6096 33756
rect 6120 33754 6176 33756
rect 6200 33754 6256 33756
rect 5960 33702 6006 33754
rect 6006 33702 6016 33754
rect 6040 33702 6070 33754
rect 6070 33702 6082 33754
rect 6082 33702 6096 33754
rect 6120 33702 6134 33754
rect 6134 33702 6146 33754
rect 6146 33702 6176 33754
rect 6200 33702 6210 33754
rect 6210 33702 6256 33754
rect 5960 33700 6016 33702
rect 6040 33700 6096 33702
rect 6120 33700 6176 33702
rect 6200 33700 6256 33702
rect 2906 33600 2962 33656
rect 6696 33210 6752 33212
rect 6776 33210 6832 33212
rect 6856 33210 6912 33212
rect 6936 33210 6992 33212
rect 6696 33158 6742 33210
rect 6742 33158 6752 33210
rect 6776 33158 6806 33210
rect 6806 33158 6818 33210
rect 6818 33158 6832 33210
rect 6856 33158 6870 33210
rect 6870 33158 6882 33210
rect 6882 33158 6912 33210
rect 6936 33158 6946 33210
rect 6946 33158 6992 33210
rect 6696 33156 6752 33158
rect 6776 33156 6832 33158
rect 6856 33156 6912 33158
rect 6936 33156 6992 33158
rect 4378 32920 4434 32976
rect 5666 32920 5722 32976
rect 5960 32666 6016 32668
rect 6040 32666 6096 32668
rect 6120 32666 6176 32668
rect 6200 32666 6256 32668
rect 5960 32614 6006 32666
rect 6006 32614 6016 32666
rect 6040 32614 6070 32666
rect 6070 32614 6082 32666
rect 6082 32614 6096 32666
rect 6120 32614 6134 32666
rect 6134 32614 6146 32666
rect 6146 32614 6176 32666
rect 6200 32614 6210 32666
rect 6210 32614 6256 32666
rect 5960 32612 6016 32614
rect 6040 32612 6096 32614
rect 6120 32612 6176 32614
rect 6200 32612 6256 32614
rect 2906 32260 2962 32296
rect 2906 32240 2908 32260
rect 2908 32240 2960 32260
rect 2960 32240 2962 32260
rect 6696 32122 6752 32124
rect 6776 32122 6832 32124
rect 6856 32122 6912 32124
rect 6936 32122 6992 32124
rect 6696 32070 6742 32122
rect 6742 32070 6752 32122
rect 6776 32070 6806 32122
rect 6806 32070 6818 32122
rect 6818 32070 6832 32122
rect 6856 32070 6870 32122
rect 6870 32070 6882 32122
rect 6882 32070 6912 32122
rect 6936 32070 6946 32122
rect 6946 32070 6992 32122
rect 7138 32104 7194 32160
rect 6696 32068 6752 32070
rect 6776 32068 6832 32070
rect 6856 32068 6912 32070
rect 6936 32068 6992 32070
rect 5960 31578 6016 31580
rect 6040 31578 6096 31580
rect 6120 31578 6176 31580
rect 6200 31578 6256 31580
rect 5960 31526 6006 31578
rect 6006 31526 6016 31578
rect 6040 31526 6070 31578
rect 6070 31526 6082 31578
rect 6082 31526 6096 31578
rect 6120 31526 6134 31578
rect 6134 31526 6146 31578
rect 6146 31526 6176 31578
rect 6200 31526 6210 31578
rect 6210 31526 6256 31578
rect 5960 31524 6016 31526
rect 6040 31524 6096 31526
rect 6120 31524 6176 31526
rect 6200 31524 6256 31526
rect 6696 31034 6752 31036
rect 6776 31034 6832 31036
rect 6856 31034 6912 31036
rect 6936 31034 6992 31036
rect 6696 30982 6742 31034
rect 6742 30982 6752 31034
rect 6776 30982 6806 31034
rect 6806 30982 6818 31034
rect 6818 30982 6832 31034
rect 6856 30982 6870 31034
rect 6870 30982 6882 31034
rect 6882 30982 6912 31034
rect 6936 30982 6946 31034
rect 6946 30982 6992 31034
rect 7138 31016 7194 31072
rect 6696 30980 6752 30982
rect 6776 30980 6832 30982
rect 6856 30980 6912 30982
rect 6936 30980 6992 30982
rect 2906 30880 2962 30936
rect 4378 30200 4434 30256
rect 5960 30490 6016 30492
rect 6040 30490 6096 30492
rect 6120 30490 6176 30492
rect 6200 30490 6256 30492
rect 5960 30438 6006 30490
rect 6006 30438 6016 30490
rect 6040 30438 6070 30490
rect 6070 30438 6082 30490
rect 6082 30438 6096 30490
rect 6120 30438 6134 30490
rect 6134 30438 6146 30490
rect 6146 30438 6176 30490
rect 6200 30438 6210 30490
rect 6210 30438 6256 30490
rect 5960 30436 6016 30438
rect 6040 30436 6096 30438
rect 6120 30436 6176 30438
rect 6200 30436 6256 30438
rect 5666 30064 5722 30120
rect 6696 29946 6752 29948
rect 6776 29946 6832 29948
rect 6856 29946 6912 29948
rect 6936 29946 6992 29948
rect 6696 29894 6742 29946
rect 6742 29894 6752 29946
rect 6776 29894 6806 29946
rect 6806 29894 6818 29946
rect 6818 29894 6832 29946
rect 6856 29894 6870 29946
rect 6870 29894 6882 29946
rect 6882 29894 6912 29946
rect 6936 29894 6946 29946
rect 6946 29894 6992 29946
rect 6696 29892 6752 29894
rect 6776 29892 6832 29894
rect 6856 29892 6912 29894
rect 6936 29892 6992 29894
rect 5960 29402 6016 29404
rect 6040 29402 6096 29404
rect 6120 29402 6176 29404
rect 6200 29402 6256 29404
rect 5960 29350 6006 29402
rect 6006 29350 6016 29402
rect 6040 29350 6070 29402
rect 6070 29350 6082 29402
rect 6082 29350 6096 29402
rect 6120 29350 6134 29402
rect 6134 29350 6146 29402
rect 6146 29350 6176 29402
rect 6200 29350 6210 29402
rect 6210 29350 6256 29402
rect 5960 29348 6016 29350
rect 6040 29348 6096 29350
rect 6120 29348 6176 29350
rect 6200 29348 6256 29350
rect 2906 28840 2962 28896
rect 6696 28858 6752 28860
rect 6776 28858 6832 28860
rect 6856 28858 6912 28860
rect 6936 28858 6992 28860
rect 6696 28806 6742 28858
rect 6742 28806 6752 28858
rect 6776 28806 6806 28858
rect 6806 28806 6818 28858
rect 6818 28806 6832 28858
rect 6856 28806 6870 28858
rect 6870 28806 6882 28858
rect 6882 28806 6912 28858
rect 6936 28806 6946 28858
rect 6946 28806 6992 28858
rect 7138 28840 7194 28896
rect 6696 28804 6752 28806
rect 6776 28804 6832 28806
rect 6856 28804 6912 28806
rect 6936 28804 6992 28806
rect 5960 28314 6016 28316
rect 6040 28314 6096 28316
rect 6120 28314 6176 28316
rect 6200 28314 6256 28316
rect 5960 28262 6006 28314
rect 6006 28262 6016 28314
rect 6040 28262 6070 28314
rect 6070 28262 6082 28314
rect 6082 28262 6096 28314
rect 6120 28262 6134 28314
rect 6134 28262 6146 28314
rect 6146 28262 6176 28314
rect 6200 28262 6210 28314
rect 6210 28262 6256 28314
rect 5960 28260 6016 28262
rect 6040 28260 6096 28262
rect 6120 28260 6176 28262
rect 6200 28260 6256 28262
rect 6696 27770 6752 27772
rect 6776 27770 6832 27772
rect 6856 27770 6912 27772
rect 6936 27770 6992 27772
rect 6696 27718 6742 27770
rect 6742 27718 6752 27770
rect 6776 27718 6806 27770
rect 6806 27718 6818 27770
rect 6818 27718 6832 27770
rect 6856 27718 6870 27770
rect 6870 27718 6882 27770
rect 6882 27718 6912 27770
rect 6936 27718 6946 27770
rect 6946 27718 6992 27770
rect 6696 27716 6752 27718
rect 6776 27716 6832 27718
rect 6856 27716 6912 27718
rect 6936 27716 6992 27718
rect 5114 27480 5170 27536
rect 5390 27480 5446 27536
rect 5960 27226 6016 27228
rect 6040 27226 6096 27228
rect 6120 27226 6176 27228
rect 6200 27226 6256 27228
rect 5960 27174 6006 27226
rect 6006 27174 6016 27226
rect 6040 27174 6070 27226
rect 6070 27174 6082 27226
rect 6082 27174 6096 27226
rect 6120 27174 6134 27226
rect 6134 27174 6146 27226
rect 6146 27174 6176 27226
rect 6200 27174 6210 27226
rect 6210 27174 6256 27226
rect 5960 27172 6016 27174
rect 6040 27172 6096 27174
rect 6120 27172 6176 27174
rect 6200 27172 6256 27174
rect 2906 26836 2908 26856
rect 2908 26836 2960 26856
rect 2960 26836 2962 26856
rect 2906 26800 2962 26836
rect 6696 26682 6752 26684
rect 6776 26682 6832 26684
rect 6856 26682 6912 26684
rect 6936 26682 6992 26684
rect 6696 26630 6742 26682
rect 6742 26630 6752 26682
rect 6776 26630 6806 26682
rect 6806 26630 6818 26682
rect 6818 26630 6832 26682
rect 6856 26630 6870 26682
rect 6870 26630 6882 26682
rect 6882 26630 6912 26682
rect 6936 26630 6946 26682
rect 6946 26630 6992 26682
rect 7138 26664 7194 26720
rect 6696 26628 6752 26630
rect 6776 26628 6832 26630
rect 6856 26628 6912 26630
rect 6936 26628 6992 26630
rect 5960 26138 6016 26140
rect 6040 26138 6096 26140
rect 6120 26138 6176 26140
rect 6200 26138 6256 26140
rect 5960 26086 6006 26138
rect 6006 26086 6016 26138
rect 6040 26086 6070 26138
rect 6070 26086 6082 26138
rect 6082 26086 6096 26138
rect 6120 26086 6134 26138
rect 6134 26086 6146 26138
rect 6146 26086 6176 26138
rect 6200 26086 6210 26138
rect 6210 26086 6256 26138
rect 5960 26084 6016 26086
rect 6040 26084 6096 26086
rect 6120 26084 6176 26086
rect 6200 26084 6256 26086
rect 6696 25594 6752 25596
rect 6776 25594 6832 25596
rect 6856 25594 6912 25596
rect 6936 25594 6992 25596
rect 6696 25542 6742 25594
rect 6742 25542 6752 25594
rect 6776 25542 6806 25594
rect 6806 25542 6818 25594
rect 6818 25542 6832 25594
rect 6856 25542 6870 25594
rect 6870 25542 6882 25594
rect 6882 25542 6912 25594
rect 6936 25542 6946 25594
rect 6946 25542 6992 25594
rect 7138 25576 7194 25632
rect 6696 25540 6752 25542
rect 6776 25540 6832 25542
rect 6856 25540 6912 25542
rect 6936 25540 6992 25542
rect 2906 25440 2962 25496
rect 4930 24760 4986 24816
rect 5960 25050 6016 25052
rect 6040 25050 6096 25052
rect 6120 25050 6176 25052
rect 6200 25050 6256 25052
rect 5960 24998 6006 25050
rect 6006 24998 6016 25050
rect 6040 24998 6070 25050
rect 6070 24998 6082 25050
rect 6082 24998 6096 25050
rect 6120 24998 6134 25050
rect 6134 24998 6146 25050
rect 6146 24998 6176 25050
rect 6200 24998 6210 25050
rect 6210 24998 6256 25050
rect 5960 24996 6016 24998
rect 6040 24996 6096 24998
rect 6120 24996 6176 24998
rect 6200 24996 6256 24998
rect 5666 24624 5722 24680
rect 6696 24506 6752 24508
rect 6776 24506 6832 24508
rect 6856 24506 6912 24508
rect 6936 24506 6992 24508
rect 6696 24454 6742 24506
rect 6742 24454 6752 24506
rect 6776 24454 6806 24506
rect 6806 24454 6818 24506
rect 6818 24454 6832 24506
rect 6856 24454 6870 24506
rect 6870 24454 6882 24506
rect 6882 24454 6912 24506
rect 6936 24454 6946 24506
rect 6946 24454 6992 24506
rect 6696 24452 6752 24454
rect 6776 24452 6832 24454
rect 6856 24452 6912 24454
rect 6936 24452 6992 24454
rect 5960 23962 6016 23964
rect 6040 23962 6096 23964
rect 6120 23962 6176 23964
rect 6200 23962 6256 23964
rect 5960 23910 6006 23962
rect 6006 23910 6016 23962
rect 6040 23910 6070 23962
rect 6070 23910 6082 23962
rect 6082 23910 6096 23962
rect 6120 23910 6134 23962
rect 6134 23910 6146 23962
rect 6146 23910 6176 23962
rect 6200 23910 6210 23962
rect 6210 23910 6256 23962
rect 5960 23908 6016 23910
rect 6040 23908 6096 23910
rect 6120 23908 6176 23910
rect 6200 23908 6256 23910
rect 2906 23400 2962 23456
rect 6696 23418 6752 23420
rect 6776 23418 6832 23420
rect 6856 23418 6912 23420
rect 6936 23418 6992 23420
rect 6696 23366 6742 23418
rect 6742 23366 6752 23418
rect 6776 23366 6806 23418
rect 6806 23366 6818 23418
rect 6818 23366 6832 23418
rect 6856 23366 6870 23418
rect 6870 23366 6882 23418
rect 6882 23366 6912 23418
rect 6936 23366 6946 23418
rect 6946 23366 6992 23418
rect 7138 23400 7194 23456
rect 6696 23364 6752 23366
rect 6776 23364 6832 23366
rect 6856 23364 6912 23366
rect 6936 23364 6992 23366
rect 5960 22874 6016 22876
rect 6040 22874 6096 22876
rect 6120 22874 6176 22876
rect 6200 22874 6256 22876
rect 5960 22822 6006 22874
rect 6006 22822 6016 22874
rect 6040 22822 6070 22874
rect 6070 22822 6082 22874
rect 6082 22822 6096 22874
rect 6120 22822 6134 22874
rect 6134 22822 6146 22874
rect 6146 22822 6176 22874
rect 6200 22822 6210 22874
rect 6210 22822 6256 22874
rect 5960 22820 6016 22822
rect 6040 22820 6096 22822
rect 6120 22820 6176 22822
rect 6200 22820 6256 22822
rect 6696 22330 6752 22332
rect 6776 22330 6832 22332
rect 6856 22330 6912 22332
rect 6936 22330 6992 22332
rect 6696 22278 6742 22330
rect 6742 22278 6752 22330
rect 6776 22278 6806 22330
rect 6806 22278 6818 22330
rect 6818 22278 6832 22330
rect 6856 22278 6870 22330
rect 6870 22278 6882 22330
rect 6882 22278 6912 22330
rect 6936 22278 6946 22330
rect 6946 22278 6992 22330
rect 7138 22312 7194 22368
rect 6696 22276 6752 22278
rect 6776 22276 6832 22278
rect 6856 22276 6912 22278
rect 6936 22276 6992 22278
rect 5206 22040 5262 22096
rect 5960 21786 6016 21788
rect 6040 21786 6096 21788
rect 6120 21786 6176 21788
rect 6200 21786 6256 21788
rect 5960 21734 6006 21786
rect 6006 21734 6016 21786
rect 6040 21734 6070 21786
rect 6070 21734 6082 21786
rect 6082 21734 6096 21786
rect 6120 21734 6134 21786
rect 6134 21734 6146 21786
rect 6146 21734 6176 21786
rect 6200 21734 6210 21786
rect 6210 21734 6256 21786
rect 5960 21732 6016 21734
rect 6040 21732 6096 21734
rect 6120 21732 6176 21734
rect 6200 21732 6256 21734
rect 2906 21396 2908 21416
rect 2908 21396 2960 21416
rect 2960 21396 2962 21416
rect 2906 21360 2962 21396
rect 6696 21242 6752 21244
rect 6776 21242 6832 21244
rect 6856 21242 6912 21244
rect 6936 21242 6992 21244
rect 6696 21190 6742 21242
rect 6742 21190 6752 21242
rect 6776 21190 6806 21242
rect 6806 21190 6818 21242
rect 6818 21190 6832 21242
rect 6856 21190 6870 21242
rect 6870 21190 6882 21242
rect 6882 21190 6912 21242
rect 6936 21190 6946 21242
rect 6946 21190 6992 21242
rect 7138 21224 7194 21280
rect 6696 21188 6752 21190
rect 6776 21188 6832 21190
rect 6856 21188 6912 21190
rect 6936 21188 6992 21190
rect 5960 20698 6016 20700
rect 6040 20698 6096 20700
rect 6120 20698 6176 20700
rect 6200 20698 6256 20700
rect 5960 20646 6006 20698
rect 6006 20646 6016 20698
rect 6040 20646 6070 20698
rect 6070 20646 6082 20698
rect 6082 20646 6096 20698
rect 6120 20646 6134 20698
rect 6134 20646 6146 20698
rect 6146 20646 6176 20698
rect 6200 20646 6210 20698
rect 6210 20646 6256 20698
rect 5960 20644 6016 20646
rect 6040 20644 6096 20646
rect 6120 20644 6176 20646
rect 6200 20644 6256 20646
rect 6696 20154 6752 20156
rect 6776 20154 6832 20156
rect 6856 20154 6912 20156
rect 6936 20154 6992 20156
rect 6696 20102 6742 20154
rect 6742 20102 6752 20154
rect 6776 20102 6806 20154
rect 6806 20102 6818 20154
rect 6818 20102 6832 20154
rect 6856 20102 6870 20154
rect 6870 20102 6882 20154
rect 6882 20102 6912 20154
rect 6936 20102 6946 20154
rect 6946 20102 6992 20154
rect 7138 20136 7194 20192
rect 6696 20100 6752 20102
rect 6776 20100 6832 20102
rect 6856 20100 6912 20102
rect 6936 20100 6992 20102
rect 2906 20000 2962 20056
rect 5960 19610 6016 19612
rect 6040 19610 6096 19612
rect 6120 19610 6176 19612
rect 6200 19610 6256 19612
rect 5960 19558 6006 19610
rect 6006 19558 6016 19610
rect 6040 19558 6070 19610
rect 6070 19558 6082 19610
rect 6082 19558 6096 19610
rect 6120 19558 6134 19610
rect 6134 19558 6146 19610
rect 6146 19558 6176 19610
rect 6200 19558 6210 19610
rect 6210 19558 6256 19610
rect 5960 19556 6016 19558
rect 6040 19556 6096 19558
rect 6120 19556 6176 19558
rect 6200 19556 6256 19558
rect 4930 19320 4986 19376
rect 6696 19066 6752 19068
rect 6776 19066 6832 19068
rect 6856 19066 6912 19068
rect 6936 19066 6992 19068
rect 6696 19014 6742 19066
rect 6742 19014 6752 19066
rect 6776 19014 6806 19066
rect 6806 19014 6818 19066
rect 6818 19014 6832 19066
rect 6856 19014 6870 19066
rect 6870 19014 6882 19066
rect 6882 19014 6912 19066
rect 6936 19014 6946 19066
rect 6946 19014 6992 19066
rect 6696 19012 6752 19014
rect 6776 19012 6832 19014
rect 6856 19012 6912 19014
rect 6936 19012 6992 19014
rect 5960 18522 6016 18524
rect 6040 18522 6096 18524
rect 6120 18522 6176 18524
rect 6200 18522 6256 18524
rect 5960 18470 6006 18522
rect 6006 18470 6016 18522
rect 6040 18470 6070 18522
rect 6070 18470 6082 18522
rect 6082 18470 6096 18522
rect 6120 18470 6134 18522
rect 6134 18470 6146 18522
rect 6146 18470 6176 18522
rect 6200 18470 6210 18522
rect 6210 18470 6256 18522
rect 5960 18468 6016 18470
rect 6040 18468 6096 18470
rect 6120 18468 6176 18470
rect 6200 18468 6256 18470
rect 5114 17960 5170 18016
rect 6696 17978 6752 17980
rect 6776 17978 6832 17980
rect 6856 17978 6912 17980
rect 6936 17978 6992 17980
rect 6696 17926 6742 17978
rect 6742 17926 6752 17978
rect 6776 17926 6806 17978
rect 6806 17926 6818 17978
rect 6818 17926 6832 17978
rect 6856 17926 6870 17978
rect 6870 17926 6882 17978
rect 6882 17926 6912 17978
rect 6936 17926 6946 17978
rect 6946 17926 6992 17978
rect 6696 17924 6752 17926
rect 6776 17924 6832 17926
rect 6856 17924 6912 17926
rect 6936 17924 6992 17926
rect 5960 17434 6016 17436
rect 6040 17434 6096 17436
rect 6120 17434 6176 17436
rect 6200 17434 6256 17436
rect 5960 17382 6006 17434
rect 6006 17382 6016 17434
rect 6040 17382 6070 17434
rect 6070 17382 6082 17434
rect 6082 17382 6096 17434
rect 6120 17382 6134 17434
rect 6134 17382 6146 17434
rect 6146 17382 6176 17434
rect 6200 17382 6210 17434
rect 6210 17382 6256 17434
rect 5960 17380 6016 17382
rect 6040 17380 6096 17382
rect 6120 17380 6176 17382
rect 6200 17380 6256 17382
rect 6696 16890 6752 16892
rect 6776 16890 6832 16892
rect 6856 16890 6912 16892
rect 6936 16890 6992 16892
rect 6696 16838 6742 16890
rect 6742 16838 6752 16890
rect 6776 16838 6806 16890
rect 6806 16838 6818 16890
rect 6818 16838 6832 16890
rect 6856 16838 6870 16890
rect 6870 16838 6882 16890
rect 6882 16838 6912 16890
rect 6936 16838 6946 16890
rect 6946 16838 6992 16890
rect 7138 16872 7194 16928
rect 6696 16836 6752 16838
rect 6776 16836 6832 16838
rect 6856 16836 6912 16838
rect 6936 16836 6992 16838
rect 5206 16600 5262 16656
rect 5960 16346 6016 16348
rect 6040 16346 6096 16348
rect 6120 16346 6176 16348
rect 6200 16346 6256 16348
rect 5960 16294 6006 16346
rect 6006 16294 6016 16346
rect 6040 16294 6070 16346
rect 6070 16294 6082 16346
rect 6082 16294 6096 16346
rect 6120 16294 6134 16346
rect 6134 16294 6146 16346
rect 6146 16294 6176 16346
rect 6200 16294 6210 16346
rect 6210 16294 6256 16346
rect 5960 16292 6016 16294
rect 6040 16292 6096 16294
rect 6120 16292 6176 16294
rect 6200 16292 6256 16294
rect 2906 15956 2908 15976
rect 2908 15956 2960 15976
rect 2960 15956 2962 15976
rect 2906 15920 2962 15956
rect 6696 15802 6752 15804
rect 6776 15802 6832 15804
rect 6856 15802 6912 15804
rect 6936 15802 6992 15804
rect 6696 15750 6742 15802
rect 6742 15750 6752 15802
rect 6776 15750 6806 15802
rect 6806 15750 6818 15802
rect 6818 15750 6832 15802
rect 6856 15750 6870 15802
rect 6870 15750 6882 15802
rect 6882 15750 6912 15802
rect 6936 15750 6946 15802
rect 6946 15750 6992 15802
rect 7598 15784 7654 15840
rect 6696 15748 6752 15750
rect 6776 15748 6832 15750
rect 6856 15748 6912 15750
rect 6936 15748 6992 15750
rect 5960 15258 6016 15260
rect 6040 15258 6096 15260
rect 6120 15258 6176 15260
rect 6200 15258 6256 15260
rect 5960 15206 6006 15258
rect 6006 15206 6016 15258
rect 6040 15206 6070 15258
rect 6070 15206 6082 15258
rect 6082 15206 6096 15258
rect 6120 15206 6134 15258
rect 6134 15206 6146 15258
rect 6146 15206 6176 15258
rect 6200 15206 6210 15258
rect 6210 15206 6256 15258
rect 5960 15204 6016 15206
rect 6040 15204 6096 15206
rect 6120 15204 6176 15206
rect 6200 15204 6256 15206
rect 6696 14714 6752 14716
rect 6776 14714 6832 14716
rect 6856 14714 6912 14716
rect 6936 14714 6992 14716
rect 6696 14662 6742 14714
rect 6742 14662 6752 14714
rect 6776 14662 6806 14714
rect 6806 14662 6818 14714
rect 6818 14662 6832 14714
rect 6856 14662 6870 14714
rect 6870 14662 6882 14714
rect 6882 14662 6912 14714
rect 6936 14662 6946 14714
rect 6946 14662 6992 14714
rect 7598 14696 7654 14752
rect 6696 14660 6752 14662
rect 6776 14660 6832 14662
rect 6856 14660 6912 14662
rect 6936 14660 6992 14662
rect 2906 14560 2962 14616
rect 4930 13880 4986 13936
rect 5960 14170 6016 14172
rect 6040 14170 6096 14172
rect 6120 14170 6176 14172
rect 6200 14170 6256 14172
rect 5960 14118 6006 14170
rect 6006 14118 6016 14170
rect 6040 14118 6070 14170
rect 6070 14118 6082 14170
rect 6082 14118 6096 14170
rect 6120 14118 6134 14170
rect 6134 14118 6146 14170
rect 6146 14118 6176 14170
rect 6200 14118 6210 14170
rect 6210 14118 6256 14170
rect 5960 14116 6016 14118
rect 6040 14116 6096 14118
rect 6120 14116 6176 14118
rect 6200 14116 6256 14118
rect 5666 13744 5722 13800
rect 6696 13626 6752 13628
rect 6776 13626 6832 13628
rect 6856 13626 6912 13628
rect 6936 13626 6992 13628
rect 6696 13574 6742 13626
rect 6742 13574 6752 13626
rect 6776 13574 6806 13626
rect 6806 13574 6818 13626
rect 6818 13574 6832 13626
rect 6856 13574 6870 13626
rect 6870 13574 6882 13626
rect 6882 13574 6912 13626
rect 6936 13574 6946 13626
rect 6946 13574 6992 13626
rect 6696 13572 6752 13574
rect 6776 13572 6832 13574
rect 6856 13572 6912 13574
rect 6936 13572 6992 13574
rect 5960 13082 6016 13084
rect 6040 13082 6096 13084
rect 6120 13082 6176 13084
rect 6200 13082 6256 13084
rect 5960 13030 6006 13082
rect 6006 13030 6016 13082
rect 6040 13030 6070 13082
rect 6070 13030 6082 13082
rect 6082 13030 6096 13082
rect 6120 13030 6134 13082
rect 6134 13030 6146 13082
rect 6146 13030 6176 13082
rect 6200 13030 6210 13082
rect 6210 13030 6256 13082
rect 5960 13028 6016 13030
rect 6040 13028 6096 13030
rect 6120 13028 6176 13030
rect 6200 13028 6256 13030
rect 6696 12538 6752 12540
rect 6776 12538 6832 12540
rect 6856 12538 6912 12540
rect 6936 12538 6992 12540
rect 6696 12486 6742 12538
rect 6742 12486 6752 12538
rect 6776 12486 6806 12538
rect 6806 12486 6818 12538
rect 6818 12486 6832 12538
rect 6856 12486 6870 12538
rect 6870 12486 6882 12538
rect 6882 12486 6912 12538
rect 6936 12486 6946 12538
rect 6946 12486 6992 12538
rect 6696 12484 6752 12486
rect 6776 12484 6832 12486
rect 6856 12484 6912 12486
rect 6936 12484 6992 12486
rect 5960 11994 6016 11996
rect 6040 11994 6096 11996
rect 6120 11994 6176 11996
rect 6200 11994 6256 11996
rect 5960 11942 6006 11994
rect 6006 11942 6016 11994
rect 6040 11942 6070 11994
rect 6070 11942 6082 11994
rect 6082 11942 6096 11994
rect 6120 11942 6134 11994
rect 6134 11942 6146 11994
rect 6146 11942 6176 11994
rect 6200 11942 6210 11994
rect 6210 11942 6256 11994
rect 5960 11940 6016 11942
rect 6040 11940 6096 11942
rect 6120 11940 6176 11942
rect 6200 11940 6256 11942
rect 6696 11450 6752 11452
rect 6776 11450 6832 11452
rect 6856 11450 6912 11452
rect 6936 11450 6992 11452
rect 6696 11398 6742 11450
rect 6742 11398 6752 11450
rect 6776 11398 6806 11450
rect 6806 11398 6818 11450
rect 6818 11398 6832 11450
rect 6856 11398 6870 11450
rect 6870 11398 6882 11450
rect 6882 11398 6912 11450
rect 6936 11398 6946 11450
rect 6946 11398 6992 11450
rect 6696 11396 6752 11398
rect 6776 11396 6832 11398
rect 6856 11396 6912 11398
rect 6936 11396 6992 11398
rect 5960 10906 6016 10908
rect 6040 10906 6096 10908
rect 6120 10906 6176 10908
rect 6200 10906 6256 10908
rect 5960 10854 6006 10906
rect 6006 10854 6016 10906
rect 6040 10854 6070 10906
rect 6070 10854 6082 10906
rect 6082 10854 6096 10906
rect 6120 10854 6134 10906
rect 6134 10854 6146 10906
rect 6146 10854 6176 10906
rect 6200 10854 6210 10906
rect 6210 10854 6256 10906
rect 5960 10852 6016 10854
rect 6040 10852 6096 10854
rect 6120 10852 6176 10854
rect 6200 10852 6256 10854
rect 7874 10480 7930 10536
rect 6696 10362 6752 10364
rect 6776 10362 6832 10364
rect 6856 10362 6912 10364
rect 6936 10362 6992 10364
rect 6696 10310 6742 10362
rect 6742 10310 6752 10362
rect 6776 10310 6806 10362
rect 6806 10310 6818 10362
rect 6818 10310 6832 10362
rect 6856 10310 6870 10362
rect 6870 10310 6882 10362
rect 6882 10310 6912 10362
rect 6936 10310 6946 10362
rect 6946 10310 6992 10362
rect 6696 10308 6752 10310
rect 6776 10308 6832 10310
rect 6856 10308 6912 10310
rect 6936 10308 6992 10310
rect 8334 47200 8390 47256
rect 8334 10344 8390 10400
rect 8150 10208 8206 10264
rect 5960 9818 6016 9820
rect 6040 9818 6096 9820
rect 6120 9818 6176 9820
rect 6200 9818 6256 9820
rect 5960 9766 6006 9818
rect 6006 9766 6016 9818
rect 6040 9766 6070 9818
rect 6070 9766 6082 9818
rect 6082 9766 6096 9818
rect 6120 9766 6134 9818
rect 6134 9766 6146 9818
rect 6146 9766 6176 9818
rect 6200 9766 6210 9818
rect 6210 9766 6256 9818
rect 5960 9764 6016 9766
rect 6040 9764 6096 9766
rect 6120 9764 6176 9766
rect 6200 9764 6256 9766
rect 6696 9274 6752 9276
rect 6776 9274 6832 9276
rect 6856 9274 6912 9276
rect 6936 9274 6992 9276
rect 6696 9222 6742 9274
rect 6742 9222 6752 9274
rect 6776 9222 6806 9274
rect 6806 9222 6818 9274
rect 6818 9222 6832 9274
rect 6856 9222 6870 9274
rect 6870 9222 6882 9274
rect 6882 9222 6912 9274
rect 6936 9222 6946 9274
rect 6946 9222 6992 9274
rect 6696 9220 6752 9222
rect 6776 9220 6832 9222
rect 6856 9220 6912 9222
rect 6936 9220 6992 9222
rect 5960 8730 6016 8732
rect 6040 8730 6096 8732
rect 6120 8730 6176 8732
rect 6200 8730 6256 8732
rect 5960 8678 6006 8730
rect 6006 8678 6016 8730
rect 6040 8678 6070 8730
rect 6070 8678 6082 8730
rect 6082 8678 6096 8730
rect 6120 8678 6134 8730
rect 6134 8678 6146 8730
rect 6146 8678 6176 8730
rect 6200 8678 6210 8730
rect 6210 8678 6256 8730
rect 5960 8676 6016 8678
rect 6040 8676 6096 8678
rect 6120 8676 6176 8678
rect 6200 8676 6256 8678
rect 9806 84192 9862 84248
rect 9622 61856 9678 61912
rect 9622 60768 9678 60824
rect 38388 88698 38444 88700
rect 38468 88698 38524 88700
rect 38548 88698 38604 88700
rect 38628 88698 38684 88700
rect 38388 88646 38434 88698
rect 38434 88646 38444 88698
rect 38468 88646 38498 88698
rect 38498 88646 38510 88698
rect 38510 88646 38524 88698
rect 38548 88646 38562 88698
rect 38562 88646 38574 88698
rect 38574 88646 38604 88698
rect 38628 88646 38638 88698
rect 38638 88646 38684 88698
rect 38388 88644 38444 88646
rect 38468 88644 38524 88646
rect 38548 88644 38604 88646
rect 38628 88644 38684 88646
rect 37728 88154 37784 88156
rect 37808 88154 37864 88156
rect 37888 88154 37944 88156
rect 37968 88154 38024 88156
rect 37728 88102 37774 88154
rect 37774 88102 37784 88154
rect 37808 88102 37838 88154
rect 37838 88102 37850 88154
rect 37850 88102 37864 88154
rect 37888 88102 37902 88154
rect 37902 88102 37914 88154
rect 37914 88102 37944 88154
rect 37968 88102 37978 88154
rect 37978 88102 38024 88154
rect 37728 88100 37784 88102
rect 37808 88100 37864 88102
rect 37888 88100 37944 88102
rect 37968 88100 38024 88102
rect 38388 87610 38444 87612
rect 38468 87610 38524 87612
rect 38548 87610 38604 87612
rect 38628 87610 38684 87612
rect 38388 87558 38434 87610
rect 38434 87558 38444 87610
rect 38468 87558 38498 87610
rect 38498 87558 38510 87610
rect 38510 87558 38524 87610
rect 38548 87558 38562 87610
rect 38562 87558 38574 87610
rect 38574 87558 38604 87610
rect 38628 87558 38638 87610
rect 38638 87558 38684 87610
rect 38388 87556 38444 87558
rect 38468 87556 38524 87558
rect 38548 87556 38604 87558
rect 38628 87556 38684 87558
rect 37728 87066 37784 87068
rect 37808 87066 37864 87068
rect 37888 87066 37944 87068
rect 37968 87066 38024 87068
rect 37728 87014 37774 87066
rect 37774 87014 37784 87066
rect 37808 87014 37838 87066
rect 37838 87014 37850 87066
rect 37850 87014 37864 87066
rect 37888 87014 37902 87066
rect 37902 87014 37914 87066
rect 37914 87014 37944 87066
rect 37968 87014 37978 87066
rect 37978 87014 38024 87066
rect 37728 87012 37784 87014
rect 37808 87012 37864 87014
rect 37888 87012 37944 87014
rect 37968 87012 38024 87014
rect 38388 86522 38444 86524
rect 38468 86522 38524 86524
rect 38548 86522 38604 86524
rect 38628 86522 38684 86524
rect 38388 86470 38434 86522
rect 38434 86470 38444 86522
rect 38468 86470 38498 86522
rect 38498 86470 38510 86522
rect 38510 86470 38524 86522
rect 38548 86470 38562 86522
rect 38562 86470 38574 86522
rect 38574 86470 38604 86522
rect 38628 86470 38638 86522
rect 38638 86470 38684 86522
rect 38388 86468 38444 86470
rect 38468 86468 38524 86470
rect 38548 86468 38604 86470
rect 38628 86468 38684 86470
rect 56728 89242 56784 89244
rect 56808 89242 56864 89244
rect 56888 89242 56944 89244
rect 56968 89242 57024 89244
rect 56728 89190 56774 89242
rect 56774 89190 56784 89242
rect 56808 89190 56838 89242
rect 56838 89190 56850 89242
rect 56850 89190 56864 89242
rect 56888 89190 56902 89242
rect 56902 89190 56914 89242
rect 56914 89190 56944 89242
rect 56968 89190 56978 89242
rect 56978 89190 57024 89242
rect 56728 89188 56784 89190
rect 56808 89188 56864 89190
rect 56888 89188 56944 89190
rect 56968 89188 57024 89190
rect 75728 89242 75784 89244
rect 75808 89242 75864 89244
rect 75888 89242 75944 89244
rect 75968 89242 76024 89244
rect 75728 89190 75774 89242
rect 75774 89190 75784 89242
rect 75808 89190 75838 89242
rect 75838 89190 75850 89242
rect 75850 89190 75864 89242
rect 75888 89190 75902 89242
rect 75902 89190 75914 89242
rect 75914 89190 75944 89242
rect 75968 89190 75978 89242
rect 75978 89190 76024 89242
rect 75728 89188 75784 89190
rect 75808 89188 75864 89190
rect 75888 89188 75944 89190
rect 75968 89188 76024 89190
rect 56728 88154 56784 88156
rect 56808 88154 56864 88156
rect 56888 88154 56944 88156
rect 56968 88154 57024 88156
rect 56728 88102 56774 88154
rect 56774 88102 56784 88154
rect 56808 88102 56838 88154
rect 56838 88102 56850 88154
rect 56850 88102 56864 88154
rect 56888 88102 56902 88154
rect 56902 88102 56914 88154
rect 56914 88102 56944 88154
rect 56968 88102 56978 88154
rect 56978 88102 57024 88154
rect 56728 88100 56784 88102
rect 56808 88100 56864 88102
rect 56888 88100 56944 88102
rect 56968 88100 57024 88102
rect 56728 87066 56784 87068
rect 56808 87066 56864 87068
rect 56888 87066 56944 87068
rect 56968 87066 57024 87068
rect 56728 87014 56774 87066
rect 56774 87014 56784 87066
rect 56808 87014 56838 87066
rect 56838 87014 56850 87066
rect 56850 87014 56864 87066
rect 56888 87014 56902 87066
rect 56902 87014 56914 87066
rect 56914 87014 56944 87066
rect 56968 87014 56978 87066
rect 56978 87014 57024 87066
rect 56728 87012 56784 87014
rect 56808 87012 56864 87014
rect 56888 87012 56944 87014
rect 56968 87012 57024 87014
rect 57388 88698 57444 88700
rect 57468 88698 57524 88700
rect 57548 88698 57604 88700
rect 57628 88698 57684 88700
rect 57388 88646 57434 88698
rect 57434 88646 57444 88698
rect 57468 88646 57498 88698
rect 57498 88646 57510 88698
rect 57510 88646 57524 88698
rect 57548 88646 57562 88698
rect 57562 88646 57574 88698
rect 57574 88646 57604 88698
rect 57628 88646 57638 88698
rect 57638 88646 57684 88698
rect 57388 88644 57444 88646
rect 57468 88644 57524 88646
rect 57548 88644 57604 88646
rect 57628 88644 57684 88646
rect 57388 87610 57444 87612
rect 57468 87610 57524 87612
rect 57548 87610 57604 87612
rect 57628 87610 57684 87612
rect 57388 87558 57434 87610
rect 57434 87558 57444 87610
rect 57468 87558 57498 87610
rect 57498 87558 57510 87610
rect 57510 87558 57524 87610
rect 57548 87558 57562 87610
rect 57562 87558 57574 87610
rect 57574 87558 57604 87610
rect 57628 87558 57638 87610
rect 57638 87558 57684 87610
rect 57388 87556 57444 87558
rect 57468 87556 57524 87558
rect 57548 87556 57604 87558
rect 57628 87556 57684 87558
rect 57388 86522 57444 86524
rect 57468 86522 57524 86524
rect 57548 86522 57604 86524
rect 57628 86522 57684 86524
rect 57388 86470 57434 86522
rect 57434 86470 57444 86522
rect 57468 86470 57498 86522
rect 57498 86470 57510 86522
rect 57510 86470 57524 86522
rect 57548 86470 57562 86522
rect 57562 86470 57574 86522
rect 57574 86470 57604 86522
rect 57628 86470 57638 86522
rect 57638 86470 57684 86522
rect 57388 86468 57444 86470
rect 57468 86468 57524 86470
rect 57548 86468 57604 86470
rect 57628 86468 57684 86470
rect 76388 88698 76444 88700
rect 76468 88698 76524 88700
rect 76548 88698 76604 88700
rect 76628 88698 76684 88700
rect 76388 88646 76434 88698
rect 76434 88646 76444 88698
rect 76468 88646 76498 88698
rect 76498 88646 76510 88698
rect 76510 88646 76524 88698
rect 76548 88646 76562 88698
rect 76562 88646 76574 88698
rect 76574 88646 76604 88698
rect 76628 88646 76638 88698
rect 76638 88646 76684 88698
rect 76388 88644 76444 88646
rect 76468 88644 76524 88646
rect 76548 88644 76604 88646
rect 76628 88644 76684 88646
rect 75728 88154 75784 88156
rect 75808 88154 75864 88156
rect 75888 88154 75944 88156
rect 75968 88154 76024 88156
rect 75728 88102 75774 88154
rect 75774 88102 75784 88154
rect 75808 88102 75838 88154
rect 75838 88102 75850 88154
rect 75850 88102 75864 88154
rect 75888 88102 75902 88154
rect 75902 88102 75914 88154
rect 75914 88102 75944 88154
rect 75968 88102 75978 88154
rect 75978 88102 76024 88154
rect 75728 88100 75784 88102
rect 75808 88100 75864 88102
rect 75888 88100 75944 88102
rect 75968 88100 76024 88102
rect 76388 87610 76444 87612
rect 76468 87610 76524 87612
rect 76548 87610 76604 87612
rect 76628 87610 76684 87612
rect 76388 87558 76434 87610
rect 76434 87558 76444 87610
rect 76468 87558 76498 87610
rect 76498 87558 76510 87610
rect 76510 87558 76524 87610
rect 76548 87558 76562 87610
rect 76562 87558 76574 87610
rect 76574 87558 76604 87610
rect 76628 87558 76638 87610
rect 76638 87558 76684 87610
rect 76388 87556 76444 87558
rect 76468 87556 76524 87558
rect 76548 87556 76604 87558
rect 76628 87556 76684 87558
rect 75728 87066 75784 87068
rect 75808 87066 75864 87068
rect 75888 87066 75944 87068
rect 75968 87066 76024 87068
rect 75728 87014 75774 87066
rect 75774 87014 75784 87066
rect 75808 87014 75838 87066
rect 75838 87014 75850 87066
rect 75850 87014 75864 87066
rect 75888 87014 75902 87066
rect 75902 87014 75914 87066
rect 75914 87014 75944 87066
rect 75968 87014 75978 87066
rect 75978 87014 76024 87066
rect 75728 87012 75784 87014
rect 75808 87012 75864 87014
rect 75888 87012 75944 87014
rect 75968 87012 76024 87014
rect 76388 86522 76444 86524
rect 76468 86522 76524 86524
rect 76548 86522 76604 86524
rect 76628 86522 76684 86524
rect 76388 86470 76434 86522
rect 76434 86470 76444 86522
rect 76468 86470 76498 86522
rect 76498 86470 76510 86522
rect 76510 86470 76524 86522
rect 76548 86470 76562 86522
rect 76562 86470 76574 86522
rect 76574 86470 76604 86522
rect 76628 86470 76638 86522
rect 76638 86470 76684 86522
rect 76388 86468 76444 86470
rect 76468 86468 76524 86470
rect 76548 86468 76604 86470
rect 76628 86468 76684 86470
rect 51436 84192 51492 84248
rect 9806 48016 9862 48072
rect 11122 48016 11178 48072
rect 13330 47200 13386 47256
rect 9806 46792 9862 46848
rect 9622 19016 9678 19072
rect 9622 17928 9678 17984
rect 50332 47200 50388 47256
rect 51436 46792 51492 46848
rect 87104 87066 87160 87068
rect 87184 87066 87240 87068
rect 87264 87066 87320 87068
rect 87344 87066 87400 87068
rect 87104 87014 87150 87066
rect 87150 87014 87160 87066
rect 87184 87014 87214 87066
rect 87214 87014 87226 87066
rect 87226 87014 87240 87066
rect 87264 87014 87278 87066
rect 87278 87014 87290 87066
rect 87290 87014 87320 87066
rect 87344 87014 87354 87066
rect 87354 87014 87400 87066
rect 87104 87012 87160 87014
rect 87184 87012 87240 87014
rect 87264 87012 87320 87014
rect 87344 87012 87400 87014
rect 87840 86522 87896 86524
rect 87920 86522 87976 86524
rect 88000 86522 88056 86524
rect 88080 86522 88136 86524
rect 87840 86470 87886 86522
rect 87886 86470 87896 86522
rect 87920 86470 87950 86522
rect 87950 86470 87962 86522
rect 87962 86470 87976 86522
rect 88000 86470 88014 86522
rect 88014 86470 88026 86522
rect 88026 86470 88056 86522
rect 88080 86470 88090 86522
rect 88090 86470 88136 86522
rect 87840 86468 87896 86470
rect 87920 86468 87976 86470
rect 88000 86468 88056 86470
rect 88080 86468 88136 86470
rect 87104 85978 87160 85980
rect 87184 85978 87240 85980
rect 87264 85978 87320 85980
rect 87344 85978 87400 85980
rect 87104 85926 87150 85978
rect 87150 85926 87160 85978
rect 87184 85926 87214 85978
rect 87214 85926 87226 85978
rect 87226 85926 87240 85978
rect 87264 85926 87278 85978
rect 87278 85926 87290 85978
rect 87290 85926 87320 85978
rect 87344 85926 87354 85978
rect 87354 85926 87400 85978
rect 87104 85924 87160 85926
rect 87184 85924 87240 85926
rect 87264 85924 87320 85926
rect 87344 85924 87400 85926
rect 87840 85434 87896 85436
rect 87920 85434 87976 85436
rect 88000 85434 88056 85436
rect 88080 85434 88136 85436
rect 87840 85382 87886 85434
rect 87886 85382 87896 85434
rect 87920 85382 87950 85434
rect 87950 85382 87962 85434
rect 87962 85382 87976 85434
rect 88000 85382 88014 85434
rect 88014 85382 88026 85434
rect 88026 85382 88056 85434
rect 88080 85382 88090 85434
rect 88090 85382 88136 85434
rect 87840 85380 87896 85382
rect 87920 85380 87976 85382
rect 88000 85380 88056 85382
rect 88080 85380 88136 85382
rect 87104 84890 87160 84892
rect 87184 84890 87240 84892
rect 87264 84890 87320 84892
rect 87344 84890 87400 84892
rect 87104 84838 87150 84890
rect 87150 84838 87160 84890
rect 87184 84838 87214 84890
rect 87214 84838 87226 84890
rect 87226 84838 87240 84890
rect 87264 84838 87278 84890
rect 87278 84838 87290 84890
rect 87290 84838 87320 84890
rect 87344 84838 87354 84890
rect 87354 84838 87400 84890
rect 87104 84836 87160 84838
rect 87184 84836 87240 84838
rect 87264 84836 87320 84838
rect 87344 84836 87400 84838
rect 87840 84346 87896 84348
rect 87920 84346 87976 84348
rect 88000 84346 88056 84348
rect 88080 84346 88136 84348
rect 87840 84294 87886 84346
rect 87886 84294 87896 84346
rect 87920 84294 87950 84346
rect 87950 84294 87962 84346
rect 87962 84294 87976 84346
rect 88000 84294 88014 84346
rect 88014 84294 88026 84346
rect 88026 84294 88056 84346
rect 88080 84294 88090 84346
rect 88090 84294 88136 84346
rect 87840 84292 87896 84294
rect 87920 84292 87976 84294
rect 88000 84292 88056 84294
rect 88080 84292 88136 84294
rect 87104 83802 87160 83804
rect 87184 83802 87240 83804
rect 87264 83802 87320 83804
rect 87344 83802 87400 83804
rect 87104 83750 87150 83802
rect 87150 83750 87160 83802
rect 87184 83750 87214 83802
rect 87214 83750 87226 83802
rect 87226 83750 87240 83802
rect 87264 83750 87278 83802
rect 87278 83750 87290 83802
rect 87290 83750 87320 83802
rect 87344 83750 87354 83802
rect 87354 83750 87400 83802
rect 87104 83748 87160 83750
rect 87184 83748 87240 83750
rect 87264 83748 87320 83750
rect 87344 83748 87400 83750
rect 87840 83258 87896 83260
rect 87920 83258 87976 83260
rect 88000 83258 88056 83260
rect 88080 83258 88136 83260
rect 87840 83206 87886 83258
rect 87886 83206 87896 83258
rect 87920 83206 87950 83258
rect 87950 83206 87962 83258
rect 87962 83206 87976 83258
rect 88000 83206 88014 83258
rect 88014 83206 88026 83258
rect 88026 83206 88056 83258
rect 88080 83206 88090 83258
rect 88090 83206 88136 83258
rect 87840 83204 87896 83206
rect 87920 83204 87976 83206
rect 88000 83204 88056 83206
rect 88080 83204 88136 83206
rect 87104 82714 87160 82716
rect 87184 82714 87240 82716
rect 87264 82714 87320 82716
rect 87344 82714 87400 82716
rect 87104 82662 87150 82714
rect 87150 82662 87160 82714
rect 87184 82662 87214 82714
rect 87214 82662 87226 82714
rect 87226 82662 87240 82714
rect 87264 82662 87278 82714
rect 87278 82662 87290 82714
rect 87290 82662 87320 82714
rect 87344 82662 87354 82714
rect 87354 82662 87400 82714
rect 87104 82660 87160 82662
rect 87184 82660 87240 82662
rect 87264 82660 87320 82662
rect 87344 82660 87400 82662
rect 87840 82170 87896 82172
rect 87920 82170 87976 82172
rect 88000 82170 88056 82172
rect 88080 82170 88136 82172
rect 87840 82118 87886 82170
rect 87886 82118 87896 82170
rect 87920 82118 87950 82170
rect 87950 82118 87962 82170
rect 87962 82118 87976 82170
rect 88000 82118 88014 82170
rect 88014 82118 88026 82170
rect 88026 82118 88056 82170
rect 88080 82118 88090 82170
rect 88090 82118 88136 82170
rect 87840 82116 87896 82118
rect 87920 82116 87976 82118
rect 88000 82116 88056 82118
rect 88080 82116 88136 82118
rect 87104 81626 87160 81628
rect 87184 81626 87240 81628
rect 87264 81626 87320 81628
rect 87344 81626 87400 81628
rect 87104 81574 87150 81626
rect 87150 81574 87160 81626
rect 87184 81574 87214 81626
rect 87214 81574 87226 81626
rect 87226 81574 87240 81626
rect 87264 81574 87278 81626
rect 87278 81574 87290 81626
rect 87290 81574 87320 81626
rect 87344 81574 87354 81626
rect 87354 81574 87400 81626
rect 87104 81572 87160 81574
rect 87184 81572 87240 81574
rect 87264 81572 87320 81574
rect 87344 81572 87400 81574
rect 87840 81082 87896 81084
rect 87920 81082 87976 81084
rect 88000 81082 88056 81084
rect 88080 81082 88136 81084
rect 87840 81030 87886 81082
rect 87886 81030 87896 81082
rect 87920 81030 87950 81082
rect 87950 81030 87962 81082
rect 87962 81030 87976 81082
rect 88000 81030 88014 81082
rect 88014 81030 88026 81082
rect 88026 81030 88056 81082
rect 88080 81030 88090 81082
rect 88090 81030 88136 81082
rect 87840 81028 87896 81030
rect 87920 81028 87976 81030
rect 88000 81028 88056 81030
rect 88080 81028 88136 81030
rect 87104 80538 87160 80540
rect 87184 80538 87240 80540
rect 87264 80538 87320 80540
rect 87344 80538 87400 80540
rect 87104 80486 87150 80538
rect 87150 80486 87160 80538
rect 87184 80486 87214 80538
rect 87214 80486 87226 80538
rect 87226 80486 87240 80538
rect 87264 80486 87278 80538
rect 87278 80486 87290 80538
rect 87290 80486 87320 80538
rect 87344 80486 87354 80538
rect 87354 80486 87400 80538
rect 88650 80520 88706 80576
rect 87104 80484 87160 80486
rect 87184 80484 87240 80486
rect 87264 80484 87320 80486
rect 87344 80484 87400 80486
rect 84326 80384 84382 80440
rect 87840 79994 87896 79996
rect 87920 79994 87976 79996
rect 88000 79994 88056 79996
rect 88080 79994 88136 79996
rect 87840 79942 87886 79994
rect 87886 79942 87896 79994
rect 87920 79942 87950 79994
rect 87950 79942 87962 79994
rect 87962 79942 87976 79994
rect 88000 79942 88014 79994
rect 88014 79942 88026 79994
rect 88026 79942 88056 79994
rect 88080 79942 88090 79994
rect 88090 79942 88136 79994
rect 87840 79940 87896 79942
rect 87920 79940 87976 79942
rect 88000 79940 88056 79942
rect 88080 79940 88136 79942
rect 87104 79450 87160 79452
rect 87184 79450 87240 79452
rect 87264 79450 87320 79452
rect 87344 79450 87400 79452
rect 87104 79398 87150 79450
rect 87150 79398 87160 79450
rect 87184 79398 87214 79450
rect 87214 79398 87226 79450
rect 87226 79398 87240 79450
rect 87264 79398 87278 79450
rect 87278 79398 87290 79450
rect 87290 79398 87320 79450
rect 87344 79398 87354 79450
rect 87354 79398 87400 79450
rect 87104 79396 87160 79398
rect 87184 79396 87240 79398
rect 87264 79396 87320 79398
rect 87344 79396 87400 79398
rect 84326 79296 84382 79352
rect 88650 79160 88706 79216
rect 87840 78906 87896 78908
rect 87920 78906 87976 78908
rect 88000 78906 88056 78908
rect 88080 78906 88136 78908
rect 87840 78854 87886 78906
rect 87886 78854 87896 78906
rect 87920 78854 87950 78906
rect 87950 78854 87962 78906
rect 87962 78854 87976 78906
rect 88000 78854 88014 78906
rect 88014 78854 88026 78906
rect 88026 78854 88056 78906
rect 88080 78854 88090 78906
rect 88090 78854 88136 78906
rect 87840 78852 87896 78854
rect 87920 78852 87976 78854
rect 88000 78852 88056 78854
rect 88080 78852 88136 78854
rect 88650 78480 88706 78536
rect 87104 78362 87160 78364
rect 87184 78362 87240 78364
rect 87264 78362 87320 78364
rect 87344 78362 87400 78364
rect 87104 78310 87150 78362
rect 87150 78310 87160 78362
rect 87184 78310 87214 78362
rect 87214 78310 87226 78362
rect 87226 78310 87240 78362
rect 87264 78310 87278 78362
rect 87278 78310 87290 78362
rect 87290 78310 87320 78362
rect 87344 78310 87354 78362
rect 87354 78310 87400 78362
rect 87104 78308 87160 78310
rect 87184 78308 87240 78310
rect 87264 78308 87320 78310
rect 87344 78308 87400 78310
rect 84326 78208 84382 78264
rect 87840 77818 87896 77820
rect 87920 77818 87976 77820
rect 88000 77818 88056 77820
rect 88080 77818 88136 77820
rect 87840 77766 87886 77818
rect 87886 77766 87896 77818
rect 87920 77766 87950 77818
rect 87950 77766 87962 77818
rect 87962 77766 87976 77818
rect 88000 77766 88014 77818
rect 88014 77766 88026 77818
rect 88026 77766 88056 77818
rect 88080 77766 88090 77818
rect 88090 77766 88136 77818
rect 87840 77764 87896 77766
rect 87920 77764 87976 77766
rect 88000 77764 88056 77766
rect 88080 77764 88136 77766
rect 87104 77274 87160 77276
rect 87184 77274 87240 77276
rect 87264 77274 87320 77276
rect 87344 77274 87400 77276
rect 87104 77222 87150 77274
rect 87150 77222 87160 77274
rect 87184 77222 87214 77274
rect 87214 77222 87226 77274
rect 87226 77222 87240 77274
rect 87264 77222 87278 77274
rect 87278 77222 87290 77274
rect 87290 77222 87320 77274
rect 87344 77222 87354 77274
rect 87354 77222 87400 77274
rect 87104 77220 87160 77222
rect 87184 77220 87240 77222
rect 87264 77220 87320 77222
rect 87344 77220 87400 77222
rect 84326 77120 84382 77176
rect 90030 77120 90086 77176
rect 87840 76730 87896 76732
rect 87920 76730 87976 76732
rect 88000 76730 88056 76732
rect 88080 76730 88136 76732
rect 87840 76678 87886 76730
rect 87886 76678 87896 76730
rect 87920 76678 87950 76730
rect 87950 76678 87962 76730
rect 87962 76678 87976 76730
rect 88000 76678 88014 76730
rect 88014 76678 88026 76730
rect 88026 76678 88056 76730
rect 88080 76678 88090 76730
rect 88090 76678 88136 76730
rect 87840 76676 87896 76678
rect 87920 76676 87976 76678
rect 88000 76676 88056 76678
rect 88080 76676 88136 76678
rect 87104 76186 87160 76188
rect 87184 76186 87240 76188
rect 87264 76186 87320 76188
rect 87344 76186 87400 76188
rect 87104 76134 87150 76186
rect 87150 76134 87160 76186
rect 87184 76134 87214 76186
rect 87214 76134 87226 76186
rect 87226 76134 87240 76186
rect 87264 76134 87278 76186
rect 87278 76134 87290 76186
rect 87290 76134 87320 76186
rect 87344 76134 87354 76186
rect 87354 76134 87400 76186
rect 87104 76132 87160 76134
rect 87184 76132 87240 76134
rect 87264 76132 87320 76134
rect 87344 76132 87400 76134
rect 84326 75984 84382 76020
rect 84326 75964 84328 75984
rect 84328 75964 84380 75984
rect 84380 75964 84382 75984
rect 88742 75796 88744 75816
rect 88744 75796 88796 75816
rect 88796 75796 88798 75816
rect 88742 75760 88798 75796
rect 87840 75642 87896 75644
rect 87920 75642 87976 75644
rect 88000 75642 88056 75644
rect 88080 75642 88136 75644
rect 87840 75590 87886 75642
rect 87886 75590 87896 75642
rect 87920 75590 87950 75642
rect 87950 75590 87962 75642
rect 87962 75590 87976 75642
rect 88000 75590 88014 75642
rect 88014 75590 88026 75642
rect 88026 75590 88056 75642
rect 88080 75590 88090 75642
rect 88090 75590 88136 75642
rect 87840 75588 87896 75590
rect 87920 75588 87976 75590
rect 88000 75588 88056 75590
rect 88080 75588 88136 75590
rect 87104 75098 87160 75100
rect 87184 75098 87240 75100
rect 87264 75098 87320 75100
rect 87344 75098 87400 75100
rect 87104 75046 87150 75098
rect 87150 75046 87160 75098
rect 87184 75046 87214 75098
rect 87214 75046 87226 75098
rect 87226 75046 87240 75098
rect 87264 75046 87278 75098
rect 87278 75046 87290 75098
rect 87290 75046 87320 75098
rect 87344 75046 87354 75098
rect 87354 75046 87400 75098
rect 88558 75080 88614 75136
rect 87104 75044 87160 75046
rect 87184 75044 87240 75046
rect 87264 75044 87320 75046
rect 87344 75044 87400 75046
rect 84326 74944 84382 75000
rect 87840 74554 87896 74556
rect 87920 74554 87976 74556
rect 88000 74554 88056 74556
rect 88080 74554 88136 74556
rect 87840 74502 87886 74554
rect 87886 74502 87896 74554
rect 87920 74502 87950 74554
rect 87950 74502 87962 74554
rect 87962 74502 87976 74554
rect 88000 74502 88014 74554
rect 88014 74502 88026 74554
rect 88026 74502 88056 74554
rect 88080 74502 88090 74554
rect 88090 74502 88136 74554
rect 87840 74500 87896 74502
rect 87920 74500 87976 74502
rect 88000 74500 88056 74502
rect 88080 74500 88136 74502
rect 87104 74010 87160 74012
rect 87184 74010 87240 74012
rect 87264 74010 87320 74012
rect 87344 74010 87400 74012
rect 87104 73958 87150 74010
rect 87150 73958 87160 74010
rect 87184 73958 87214 74010
rect 87214 73958 87226 74010
rect 87226 73958 87240 74010
rect 87264 73958 87278 74010
rect 87278 73958 87290 74010
rect 87290 73958 87320 74010
rect 87344 73958 87354 74010
rect 87354 73958 87400 74010
rect 87104 73956 87160 73958
rect 87184 73956 87240 73958
rect 87264 73956 87320 73958
rect 87344 73956 87400 73958
rect 84326 73856 84382 73912
rect 88558 73720 88614 73776
rect 87840 73466 87896 73468
rect 87920 73466 87976 73468
rect 88000 73466 88056 73468
rect 88080 73466 88136 73468
rect 87840 73414 87886 73466
rect 87886 73414 87896 73466
rect 87920 73414 87950 73466
rect 87950 73414 87962 73466
rect 87962 73414 87976 73466
rect 88000 73414 88014 73466
rect 88014 73414 88026 73466
rect 88026 73414 88056 73466
rect 88080 73414 88090 73466
rect 88090 73414 88136 73466
rect 87840 73412 87896 73414
rect 87920 73412 87976 73414
rect 88000 73412 88056 73414
rect 88080 73412 88136 73414
rect 88650 73040 88706 73096
rect 87104 72922 87160 72924
rect 87184 72922 87240 72924
rect 87264 72922 87320 72924
rect 87344 72922 87400 72924
rect 87104 72870 87150 72922
rect 87150 72870 87160 72922
rect 87184 72870 87214 72922
rect 87214 72870 87226 72922
rect 87226 72870 87240 72922
rect 87264 72870 87278 72922
rect 87278 72870 87290 72922
rect 87290 72870 87320 72922
rect 87344 72870 87354 72922
rect 87354 72870 87400 72922
rect 87104 72868 87160 72870
rect 87184 72868 87240 72870
rect 87264 72868 87320 72870
rect 87344 72868 87400 72870
rect 84326 72768 84382 72824
rect 87840 72378 87896 72380
rect 87920 72378 87976 72380
rect 88000 72378 88056 72380
rect 88080 72378 88136 72380
rect 87840 72326 87886 72378
rect 87886 72326 87896 72378
rect 87920 72326 87950 72378
rect 87950 72326 87962 72378
rect 87962 72326 87976 72378
rect 88000 72326 88014 72378
rect 88014 72326 88026 72378
rect 88026 72326 88056 72378
rect 88080 72326 88090 72378
rect 88090 72326 88136 72378
rect 87840 72324 87896 72326
rect 87920 72324 87976 72326
rect 88000 72324 88056 72326
rect 88080 72324 88136 72326
rect 87178 71988 87180 72008
rect 87180 71988 87232 72008
rect 87232 71988 87234 72008
rect 87178 71952 87234 71988
rect 87104 71834 87160 71836
rect 87184 71834 87240 71836
rect 87264 71834 87320 71836
rect 87344 71834 87400 71836
rect 87104 71782 87150 71834
rect 87150 71782 87160 71834
rect 87184 71782 87214 71834
rect 87214 71782 87226 71834
rect 87226 71782 87240 71834
rect 87264 71782 87278 71834
rect 87278 71782 87290 71834
rect 87290 71782 87320 71834
rect 87344 71782 87354 71834
rect 87354 71782 87400 71834
rect 87104 71780 87160 71782
rect 87184 71780 87240 71782
rect 87264 71780 87320 71782
rect 87344 71780 87400 71782
rect 90122 71680 90178 71736
rect 87840 71290 87896 71292
rect 87920 71290 87976 71292
rect 88000 71290 88056 71292
rect 88080 71290 88136 71292
rect 87840 71238 87886 71290
rect 87886 71238 87896 71290
rect 87920 71238 87950 71290
rect 87950 71238 87962 71290
rect 87962 71238 87976 71290
rect 88000 71238 88014 71290
rect 88014 71238 88026 71290
rect 88026 71238 88056 71290
rect 88080 71238 88090 71290
rect 88090 71238 88136 71290
rect 87840 71236 87896 71238
rect 87920 71236 87976 71238
rect 88000 71236 88056 71238
rect 88080 71236 88136 71238
rect 87104 70746 87160 70748
rect 87184 70746 87240 70748
rect 87264 70746 87320 70748
rect 87344 70746 87400 70748
rect 87104 70694 87150 70746
rect 87150 70694 87160 70746
rect 87184 70694 87214 70746
rect 87214 70694 87226 70746
rect 87226 70694 87240 70746
rect 87264 70694 87278 70746
rect 87278 70694 87290 70746
rect 87290 70694 87320 70746
rect 87344 70694 87354 70746
rect 87354 70694 87400 70746
rect 87104 70692 87160 70694
rect 87184 70692 87240 70694
rect 87264 70692 87320 70694
rect 87344 70692 87400 70694
rect 84326 70592 84382 70648
rect 89938 70356 89940 70376
rect 89940 70356 89992 70376
rect 89992 70356 89994 70376
rect 89938 70320 89994 70356
rect 87840 70202 87896 70204
rect 87920 70202 87976 70204
rect 88000 70202 88056 70204
rect 88080 70202 88136 70204
rect 87840 70150 87886 70202
rect 87886 70150 87896 70202
rect 87920 70150 87950 70202
rect 87950 70150 87962 70202
rect 87962 70150 87976 70202
rect 88000 70150 88014 70202
rect 88014 70150 88026 70202
rect 88026 70150 88056 70202
rect 88080 70150 88090 70202
rect 88090 70150 88136 70202
rect 87840 70148 87896 70150
rect 87920 70148 87976 70150
rect 88000 70148 88056 70150
rect 88080 70148 88136 70150
rect 87104 69658 87160 69660
rect 87184 69658 87240 69660
rect 87264 69658 87320 69660
rect 87344 69658 87400 69660
rect 87104 69606 87150 69658
rect 87150 69606 87160 69658
rect 87184 69606 87214 69658
rect 87214 69606 87226 69658
rect 87226 69606 87240 69658
rect 87264 69606 87278 69658
rect 87278 69606 87290 69658
rect 87290 69606 87320 69658
rect 87344 69606 87354 69658
rect 87354 69606 87400 69658
rect 88558 69640 88614 69696
rect 87104 69604 87160 69606
rect 87184 69604 87240 69606
rect 87264 69604 87320 69606
rect 87344 69604 87400 69606
rect 84326 69504 84382 69560
rect 87840 69114 87896 69116
rect 87920 69114 87976 69116
rect 88000 69114 88056 69116
rect 88080 69114 88136 69116
rect 87840 69062 87886 69114
rect 87886 69062 87896 69114
rect 87920 69062 87950 69114
rect 87950 69062 87962 69114
rect 87962 69062 87976 69114
rect 88000 69062 88014 69114
rect 88014 69062 88026 69114
rect 88026 69062 88056 69114
rect 88080 69062 88090 69114
rect 88090 69062 88136 69114
rect 87840 69060 87896 69062
rect 87920 69060 87976 69062
rect 88000 69060 88056 69062
rect 88080 69060 88136 69062
rect 89938 68960 89994 69016
rect 87104 68570 87160 68572
rect 87184 68570 87240 68572
rect 87264 68570 87320 68572
rect 87344 68570 87400 68572
rect 87104 68518 87150 68570
rect 87150 68518 87160 68570
rect 87184 68518 87214 68570
rect 87214 68518 87226 68570
rect 87226 68518 87240 68570
rect 87264 68518 87278 68570
rect 87278 68518 87290 68570
rect 87290 68518 87320 68570
rect 87344 68518 87354 68570
rect 87354 68518 87400 68570
rect 87104 68516 87160 68518
rect 87184 68516 87240 68518
rect 87264 68516 87320 68518
rect 87344 68516 87400 68518
rect 84326 68416 84382 68472
rect 88650 68280 88706 68336
rect 87840 68026 87896 68028
rect 87920 68026 87976 68028
rect 88000 68026 88056 68028
rect 88080 68026 88136 68028
rect 87840 67974 87886 68026
rect 87886 67974 87896 68026
rect 87920 67974 87950 68026
rect 87950 67974 87962 68026
rect 87962 67974 87976 68026
rect 88000 67974 88014 68026
rect 88014 67974 88026 68026
rect 88026 67974 88056 68026
rect 88080 67974 88090 68026
rect 88090 67974 88136 68026
rect 87840 67972 87896 67974
rect 87920 67972 87976 67974
rect 88000 67972 88056 67974
rect 88080 67972 88136 67974
rect 88650 67600 88706 67656
rect 87104 67482 87160 67484
rect 87184 67482 87240 67484
rect 87264 67482 87320 67484
rect 87344 67482 87400 67484
rect 87104 67430 87150 67482
rect 87150 67430 87160 67482
rect 87184 67430 87214 67482
rect 87214 67430 87226 67482
rect 87226 67430 87240 67482
rect 87264 67430 87278 67482
rect 87278 67430 87290 67482
rect 87290 67430 87320 67482
rect 87344 67430 87354 67482
rect 87354 67430 87400 67482
rect 87104 67428 87160 67430
rect 87184 67428 87240 67430
rect 87264 67428 87320 67430
rect 87344 67428 87400 67430
rect 84326 67328 84382 67384
rect 87840 66938 87896 66940
rect 87920 66938 87976 66940
rect 88000 66938 88056 66940
rect 88080 66938 88136 66940
rect 87840 66886 87886 66938
rect 87886 66886 87896 66938
rect 87920 66886 87950 66938
rect 87950 66886 87962 66938
rect 87962 66886 87976 66938
rect 88000 66886 88014 66938
rect 88014 66886 88026 66938
rect 88026 66886 88056 66938
rect 88080 66886 88090 66938
rect 88090 66886 88136 66938
rect 87840 66884 87896 66886
rect 87920 66884 87976 66886
rect 88000 66884 88056 66886
rect 88080 66884 88136 66886
rect 87104 66394 87160 66396
rect 87184 66394 87240 66396
rect 87264 66394 87320 66396
rect 87344 66394 87400 66396
rect 87104 66342 87150 66394
rect 87150 66342 87160 66394
rect 87184 66342 87214 66394
rect 87214 66342 87226 66394
rect 87226 66342 87240 66394
rect 87264 66342 87278 66394
rect 87278 66342 87290 66394
rect 87290 66342 87320 66394
rect 87344 66342 87354 66394
rect 87354 66342 87400 66394
rect 87104 66340 87160 66342
rect 87184 66340 87240 66342
rect 87264 66340 87320 66342
rect 87344 66340 87400 66342
rect 90122 66240 90178 66296
rect 87454 66104 87510 66160
rect 87840 65850 87896 65852
rect 87920 65850 87976 65852
rect 88000 65850 88056 65852
rect 88080 65850 88136 65852
rect 87840 65798 87886 65850
rect 87886 65798 87896 65850
rect 87920 65798 87950 65850
rect 87950 65798 87962 65850
rect 87962 65798 87976 65850
rect 88000 65798 88014 65850
rect 88014 65798 88026 65850
rect 88026 65798 88056 65850
rect 88080 65798 88090 65850
rect 88090 65798 88136 65850
rect 87840 65796 87896 65798
rect 87920 65796 87976 65798
rect 88000 65796 88056 65798
rect 88080 65796 88136 65798
rect 87104 65306 87160 65308
rect 87184 65306 87240 65308
rect 87264 65306 87320 65308
rect 87344 65306 87400 65308
rect 87104 65254 87150 65306
rect 87150 65254 87160 65306
rect 87184 65254 87214 65306
rect 87214 65254 87226 65306
rect 87226 65254 87240 65306
rect 87264 65254 87278 65306
rect 87278 65254 87290 65306
rect 87290 65254 87320 65306
rect 87344 65254 87354 65306
rect 87354 65254 87400 65306
rect 87104 65252 87160 65254
rect 87184 65252 87240 65254
rect 87264 65252 87320 65254
rect 87344 65252 87400 65254
rect 84326 65084 84382 65140
rect 89938 64900 89994 64936
rect 89938 64880 89940 64900
rect 89940 64880 89992 64900
rect 89992 64880 89994 64900
rect 87840 64762 87896 64764
rect 87920 64762 87976 64764
rect 88000 64762 88056 64764
rect 88080 64762 88136 64764
rect 87840 64710 87886 64762
rect 87886 64710 87896 64762
rect 87920 64710 87950 64762
rect 87950 64710 87962 64762
rect 87962 64710 87976 64762
rect 88000 64710 88014 64762
rect 88014 64710 88026 64762
rect 88026 64710 88056 64762
rect 88080 64710 88090 64762
rect 88090 64710 88136 64762
rect 87840 64708 87896 64710
rect 87920 64708 87976 64710
rect 88000 64708 88056 64710
rect 88080 64708 88136 64710
rect 87104 64218 87160 64220
rect 87184 64218 87240 64220
rect 87264 64218 87320 64220
rect 87344 64218 87400 64220
rect 87104 64166 87150 64218
rect 87150 64166 87160 64218
rect 87184 64166 87214 64218
rect 87214 64166 87226 64218
rect 87226 64166 87240 64218
rect 87264 64166 87278 64218
rect 87278 64166 87290 64218
rect 87290 64166 87320 64218
rect 87344 64166 87354 64218
rect 87354 64166 87400 64218
rect 88558 64200 88614 64256
rect 87104 64164 87160 64166
rect 87184 64164 87240 64166
rect 87264 64164 87320 64166
rect 87344 64164 87400 64166
rect 84326 64064 84382 64120
rect 87840 63674 87896 63676
rect 87920 63674 87976 63676
rect 88000 63674 88056 63676
rect 88080 63674 88136 63676
rect 87840 63622 87886 63674
rect 87886 63622 87896 63674
rect 87920 63622 87950 63674
rect 87950 63622 87962 63674
rect 87962 63622 87976 63674
rect 88000 63622 88014 63674
rect 88014 63622 88026 63674
rect 88026 63622 88056 63674
rect 88080 63622 88090 63674
rect 88090 63622 88136 63674
rect 87840 63620 87896 63622
rect 87920 63620 87976 63622
rect 88000 63620 88056 63622
rect 88080 63620 88136 63622
rect 87104 63130 87160 63132
rect 87184 63130 87240 63132
rect 87264 63130 87320 63132
rect 87344 63130 87400 63132
rect 87104 63078 87150 63130
rect 87150 63078 87160 63130
rect 87184 63078 87214 63130
rect 87214 63078 87226 63130
rect 87226 63078 87240 63130
rect 87264 63078 87278 63130
rect 87278 63078 87290 63130
rect 87290 63078 87320 63130
rect 87344 63078 87354 63130
rect 87354 63078 87400 63130
rect 87104 63076 87160 63078
rect 87184 63076 87240 63078
rect 87264 63076 87320 63078
rect 87344 63076 87400 63078
rect 84326 62976 84382 63032
rect 88558 62840 88614 62896
rect 87840 62586 87896 62588
rect 87920 62586 87976 62588
rect 88000 62586 88056 62588
rect 88080 62586 88136 62588
rect 87840 62534 87886 62586
rect 87886 62534 87896 62586
rect 87920 62534 87950 62586
rect 87950 62534 87962 62586
rect 87962 62534 87976 62586
rect 88000 62534 88014 62586
rect 88014 62534 88026 62586
rect 88026 62534 88056 62586
rect 88080 62534 88090 62586
rect 88090 62534 88136 62586
rect 87840 62532 87896 62534
rect 87920 62532 87976 62534
rect 88000 62532 88056 62534
rect 88080 62532 88136 62534
rect 88374 62160 88430 62216
rect 89938 62160 89994 62216
rect 87104 62042 87160 62044
rect 87184 62042 87240 62044
rect 87264 62042 87320 62044
rect 87344 62042 87400 62044
rect 87104 61990 87150 62042
rect 87150 61990 87160 62042
rect 87184 61990 87214 62042
rect 87214 61990 87226 62042
rect 87226 61990 87240 62042
rect 87264 61990 87278 62042
rect 87278 61990 87290 62042
rect 87290 61990 87320 62042
rect 87344 61990 87354 62042
rect 87354 61990 87400 62042
rect 87104 61988 87160 61990
rect 87184 61988 87240 61990
rect 87264 61988 87320 61990
rect 87344 61988 87400 61990
rect 87840 61498 87896 61500
rect 87920 61498 87976 61500
rect 88000 61498 88056 61500
rect 88080 61498 88136 61500
rect 87840 61446 87886 61498
rect 87886 61446 87896 61498
rect 87920 61446 87950 61498
rect 87950 61446 87962 61498
rect 87962 61446 87976 61498
rect 88000 61446 88014 61498
rect 88014 61446 88026 61498
rect 88026 61446 88056 61498
rect 88080 61446 88090 61498
rect 88090 61446 88136 61498
rect 87840 61444 87896 61446
rect 87920 61444 87976 61446
rect 88000 61444 88056 61446
rect 88080 61444 88136 61446
rect 87104 60954 87160 60956
rect 87184 60954 87240 60956
rect 87264 60954 87320 60956
rect 87344 60954 87400 60956
rect 87104 60902 87150 60954
rect 87150 60902 87160 60954
rect 87184 60902 87214 60954
rect 87214 60902 87226 60954
rect 87226 60902 87240 60954
rect 87264 60902 87278 60954
rect 87278 60902 87290 60954
rect 87290 60902 87320 60954
rect 87344 60902 87354 60954
rect 87354 60902 87400 60954
rect 87104 60900 87160 60902
rect 87184 60900 87240 60902
rect 87264 60900 87320 60902
rect 87344 60900 87400 60902
rect 89938 60800 89994 60856
rect 88374 60664 88430 60720
rect 87840 60410 87896 60412
rect 87920 60410 87976 60412
rect 88000 60410 88056 60412
rect 88080 60410 88136 60412
rect 87840 60358 87886 60410
rect 87886 60358 87896 60410
rect 87920 60358 87950 60410
rect 87950 60358 87962 60410
rect 87962 60358 87976 60410
rect 88000 60358 88014 60410
rect 88014 60358 88026 60410
rect 88026 60358 88056 60410
rect 88080 60358 88090 60410
rect 88090 60358 88136 60410
rect 87840 60356 87896 60358
rect 87920 60356 87976 60358
rect 88000 60356 88056 60358
rect 88080 60356 88136 60358
rect 87104 59866 87160 59868
rect 87184 59866 87240 59868
rect 87264 59866 87320 59868
rect 87344 59866 87400 59868
rect 87104 59814 87150 59866
rect 87150 59814 87160 59866
rect 87184 59814 87214 59866
rect 87214 59814 87226 59866
rect 87226 59814 87240 59866
rect 87264 59814 87278 59866
rect 87278 59814 87290 59866
rect 87290 59814 87320 59866
rect 87344 59814 87354 59866
rect 87354 59814 87400 59866
rect 87104 59812 87160 59814
rect 87184 59812 87240 59814
rect 87264 59812 87320 59814
rect 87344 59812 87400 59814
rect 84326 59644 84382 59700
rect 89938 59460 89994 59496
rect 89938 59440 89940 59460
rect 89940 59440 89992 59460
rect 89992 59440 89994 59460
rect 87840 59322 87896 59324
rect 87920 59322 87976 59324
rect 88000 59322 88056 59324
rect 88080 59322 88136 59324
rect 87840 59270 87886 59322
rect 87886 59270 87896 59322
rect 87920 59270 87950 59322
rect 87950 59270 87962 59322
rect 87962 59270 87976 59322
rect 88000 59270 88014 59322
rect 88014 59270 88026 59322
rect 88026 59270 88056 59322
rect 88080 59270 88090 59322
rect 88090 59270 88136 59322
rect 87840 59268 87896 59270
rect 87920 59268 87976 59270
rect 88000 59268 88056 59270
rect 88080 59268 88136 59270
rect 87104 58778 87160 58780
rect 87184 58778 87240 58780
rect 87264 58778 87320 58780
rect 87344 58778 87400 58780
rect 87104 58726 87150 58778
rect 87150 58726 87160 58778
rect 87184 58726 87214 58778
rect 87214 58726 87226 58778
rect 87226 58726 87240 58778
rect 87264 58726 87278 58778
rect 87278 58726 87290 58778
rect 87290 58726 87320 58778
rect 87344 58726 87354 58778
rect 87354 58726 87400 58778
rect 88558 58760 88614 58816
rect 87104 58724 87160 58726
rect 87184 58724 87240 58726
rect 87264 58724 87320 58726
rect 87344 58724 87400 58726
rect 84326 58624 84382 58680
rect 87840 58234 87896 58236
rect 87920 58234 87976 58236
rect 88000 58234 88056 58236
rect 88080 58234 88136 58236
rect 87840 58182 87886 58234
rect 87886 58182 87896 58234
rect 87920 58182 87950 58234
rect 87950 58182 87962 58234
rect 87962 58182 87976 58234
rect 88000 58182 88014 58234
rect 88014 58182 88026 58234
rect 88026 58182 88056 58234
rect 88080 58182 88090 58234
rect 88090 58182 88136 58234
rect 87840 58180 87896 58182
rect 87920 58180 87976 58182
rect 88000 58180 88056 58182
rect 88080 58180 88136 58182
rect 87104 57690 87160 57692
rect 87184 57690 87240 57692
rect 87264 57690 87320 57692
rect 87344 57690 87400 57692
rect 87104 57638 87150 57690
rect 87150 57638 87160 57690
rect 87184 57638 87214 57690
rect 87214 57638 87226 57690
rect 87226 57638 87240 57690
rect 87264 57638 87278 57690
rect 87278 57638 87290 57690
rect 87290 57638 87320 57690
rect 87344 57638 87354 57690
rect 87354 57638 87400 57690
rect 87104 57636 87160 57638
rect 87184 57636 87240 57638
rect 87264 57636 87320 57638
rect 87344 57636 87400 57638
rect 84326 57536 84382 57592
rect 88558 57400 88614 57456
rect 87840 57146 87896 57148
rect 87920 57146 87976 57148
rect 88000 57146 88056 57148
rect 88080 57146 88136 57148
rect 87840 57094 87886 57146
rect 87886 57094 87896 57146
rect 87920 57094 87950 57146
rect 87950 57094 87962 57146
rect 87962 57094 87976 57146
rect 88000 57094 88014 57146
rect 88014 57094 88026 57146
rect 88026 57094 88056 57146
rect 88080 57094 88090 57146
rect 88090 57094 88136 57146
rect 87840 57092 87896 57094
rect 87920 57092 87976 57094
rect 88000 57092 88056 57094
rect 88080 57092 88136 57094
rect 88282 56720 88338 56776
rect 89938 56720 89994 56776
rect 87104 56602 87160 56604
rect 87184 56602 87240 56604
rect 87264 56602 87320 56604
rect 87344 56602 87400 56604
rect 87104 56550 87150 56602
rect 87150 56550 87160 56602
rect 87184 56550 87214 56602
rect 87214 56550 87226 56602
rect 87226 56550 87240 56602
rect 87264 56550 87278 56602
rect 87278 56550 87290 56602
rect 87290 56550 87320 56602
rect 87344 56550 87354 56602
rect 87354 56550 87400 56602
rect 87104 56548 87160 56550
rect 87184 56548 87240 56550
rect 87264 56548 87320 56550
rect 87344 56548 87400 56550
rect 87840 56058 87896 56060
rect 87920 56058 87976 56060
rect 88000 56058 88056 56060
rect 88080 56058 88136 56060
rect 87840 56006 87886 56058
rect 87886 56006 87896 56058
rect 87920 56006 87950 56058
rect 87950 56006 87962 56058
rect 87962 56006 87976 56058
rect 88000 56006 88014 56058
rect 88014 56006 88026 56058
rect 88026 56006 88056 56058
rect 88080 56006 88090 56058
rect 88090 56006 88136 56058
rect 87840 56004 87896 56006
rect 87920 56004 87976 56006
rect 88000 56004 88056 56006
rect 88080 56004 88136 56006
rect 87104 55514 87160 55516
rect 87184 55514 87240 55516
rect 87264 55514 87320 55516
rect 87344 55514 87400 55516
rect 87104 55462 87150 55514
rect 87150 55462 87160 55514
rect 87184 55462 87214 55514
rect 87214 55462 87226 55514
rect 87226 55462 87240 55514
rect 87264 55462 87278 55514
rect 87278 55462 87290 55514
rect 87290 55462 87320 55514
rect 87344 55462 87354 55514
rect 87354 55462 87400 55514
rect 87104 55460 87160 55462
rect 87184 55460 87240 55462
rect 87264 55460 87320 55462
rect 87344 55460 87400 55462
rect 89938 55360 89994 55416
rect 88374 55224 88430 55280
rect 87840 54970 87896 54972
rect 87920 54970 87976 54972
rect 88000 54970 88056 54972
rect 88080 54970 88136 54972
rect 87840 54918 87886 54970
rect 87886 54918 87896 54970
rect 87920 54918 87950 54970
rect 87950 54918 87962 54970
rect 87962 54918 87976 54970
rect 88000 54918 88014 54970
rect 88014 54918 88026 54970
rect 88026 54918 88056 54970
rect 88080 54918 88090 54970
rect 88090 54918 88136 54970
rect 87840 54916 87896 54918
rect 87920 54916 87976 54918
rect 88000 54916 88056 54918
rect 88080 54916 88136 54918
rect 87104 54426 87160 54428
rect 87184 54426 87240 54428
rect 87264 54426 87320 54428
rect 87344 54426 87400 54428
rect 87104 54374 87150 54426
rect 87150 54374 87160 54426
rect 87184 54374 87214 54426
rect 87214 54374 87226 54426
rect 87226 54374 87240 54426
rect 87264 54374 87278 54426
rect 87278 54374 87290 54426
rect 87290 54374 87320 54426
rect 87344 54374 87354 54426
rect 87354 54374 87400 54426
rect 87104 54372 87160 54374
rect 87184 54372 87240 54374
rect 87264 54372 87320 54374
rect 87344 54372 87400 54374
rect 84326 54204 84382 54260
rect 89938 54036 89940 54056
rect 89940 54036 89992 54056
rect 89992 54036 89994 54056
rect 89938 54000 89994 54036
rect 87840 53882 87896 53884
rect 87920 53882 87976 53884
rect 88000 53882 88056 53884
rect 88080 53882 88136 53884
rect 87840 53830 87886 53882
rect 87886 53830 87896 53882
rect 87920 53830 87950 53882
rect 87950 53830 87962 53882
rect 87962 53830 87976 53882
rect 88000 53830 88014 53882
rect 88014 53830 88026 53882
rect 88026 53830 88056 53882
rect 88080 53830 88090 53882
rect 88090 53830 88136 53882
rect 87840 53828 87896 53830
rect 87920 53828 87976 53830
rect 88000 53828 88056 53830
rect 88080 53828 88136 53830
rect 87104 53338 87160 53340
rect 87184 53338 87240 53340
rect 87264 53338 87320 53340
rect 87344 53338 87400 53340
rect 87104 53286 87150 53338
rect 87150 53286 87160 53338
rect 87184 53286 87214 53338
rect 87214 53286 87226 53338
rect 87226 53286 87240 53338
rect 87264 53286 87278 53338
rect 87278 53286 87290 53338
rect 87290 53286 87320 53338
rect 87344 53286 87354 53338
rect 87354 53286 87400 53338
rect 88558 53320 88614 53376
rect 87104 53284 87160 53286
rect 87184 53284 87240 53286
rect 87264 53284 87320 53286
rect 87344 53284 87400 53286
rect 84326 53184 84382 53240
rect 87840 52794 87896 52796
rect 87920 52794 87976 52796
rect 88000 52794 88056 52796
rect 88080 52794 88136 52796
rect 87840 52742 87886 52794
rect 87886 52742 87896 52794
rect 87920 52742 87950 52794
rect 87950 52742 87962 52794
rect 87962 52742 87976 52794
rect 88000 52742 88014 52794
rect 88014 52742 88026 52794
rect 88026 52742 88056 52794
rect 88080 52742 88090 52794
rect 88090 52742 88136 52794
rect 87840 52740 87896 52742
rect 87920 52740 87976 52742
rect 88000 52740 88056 52742
rect 88080 52740 88136 52742
rect 89938 52640 89994 52696
rect 87104 52250 87160 52252
rect 87184 52250 87240 52252
rect 87264 52250 87320 52252
rect 87344 52250 87400 52252
rect 87104 52198 87150 52250
rect 87150 52198 87160 52250
rect 87184 52198 87214 52250
rect 87214 52198 87226 52250
rect 87226 52198 87240 52250
rect 87264 52198 87278 52250
rect 87278 52198 87290 52250
rect 87290 52198 87320 52250
rect 87344 52198 87354 52250
rect 87354 52198 87400 52250
rect 87104 52196 87160 52198
rect 87184 52196 87240 52198
rect 87264 52196 87320 52198
rect 87344 52196 87400 52198
rect 84326 52096 84382 52152
rect 88558 51960 88614 52016
rect 87840 51706 87896 51708
rect 87920 51706 87976 51708
rect 88000 51706 88056 51708
rect 88080 51706 88136 51708
rect 87840 51654 87886 51706
rect 87886 51654 87896 51706
rect 87920 51654 87950 51706
rect 87950 51654 87962 51706
rect 87962 51654 87976 51706
rect 88000 51654 88014 51706
rect 88014 51654 88026 51706
rect 88026 51654 88056 51706
rect 88080 51654 88090 51706
rect 88090 51654 88136 51706
rect 87840 51652 87896 51654
rect 87920 51652 87976 51654
rect 88000 51652 88056 51654
rect 88080 51652 88136 51654
rect 87104 51162 87160 51164
rect 87184 51162 87240 51164
rect 87264 51162 87320 51164
rect 87344 51162 87400 51164
rect 87104 51110 87150 51162
rect 87150 51110 87160 51162
rect 87184 51110 87214 51162
rect 87214 51110 87226 51162
rect 87226 51110 87240 51162
rect 87264 51110 87278 51162
rect 87278 51110 87290 51162
rect 87290 51110 87320 51162
rect 87344 51110 87354 51162
rect 87354 51110 87400 51162
rect 87104 51108 87160 51110
rect 87184 51108 87240 51110
rect 87264 51108 87320 51110
rect 87344 51108 87400 51110
rect 88558 51316 88560 51336
rect 88560 51316 88612 51336
rect 88612 51316 88614 51336
rect 88558 51280 88614 51316
rect 88374 50872 88430 50928
rect 87840 50618 87896 50620
rect 87920 50618 87976 50620
rect 88000 50618 88056 50620
rect 88080 50618 88136 50620
rect 87840 50566 87886 50618
rect 87886 50566 87896 50618
rect 87920 50566 87950 50618
rect 87950 50566 87962 50618
rect 87962 50566 87976 50618
rect 88000 50566 88014 50618
rect 88014 50566 88026 50618
rect 88026 50566 88056 50618
rect 88080 50566 88090 50618
rect 88090 50566 88136 50618
rect 87840 50564 87896 50566
rect 87920 50564 87976 50566
rect 88000 50564 88056 50566
rect 88080 50564 88136 50566
rect 87104 50074 87160 50076
rect 87184 50074 87240 50076
rect 87264 50074 87320 50076
rect 87344 50074 87400 50076
rect 87104 50022 87150 50074
rect 87150 50022 87160 50074
rect 87184 50022 87214 50074
rect 87214 50022 87226 50074
rect 87226 50022 87240 50074
rect 87264 50022 87278 50074
rect 87278 50022 87290 50074
rect 87290 50022 87320 50074
rect 87344 50022 87354 50074
rect 87354 50022 87400 50074
rect 87104 50020 87160 50022
rect 87184 50020 87240 50022
rect 87264 50020 87320 50022
rect 87344 50020 87400 50022
rect 87840 49530 87896 49532
rect 87920 49530 87976 49532
rect 88000 49530 88056 49532
rect 88080 49530 88136 49532
rect 87840 49478 87886 49530
rect 87886 49478 87896 49530
rect 87920 49478 87950 49530
rect 87950 49478 87962 49530
rect 87962 49478 87976 49530
rect 88000 49478 88014 49530
rect 88014 49478 88026 49530
rect 88026 49478 88056 49530
rect 88080 49478 88090 49530
rect 88090 49478 88136 49530
rect 87840 49476 87896 49478
rect 87920 49476 87976 49478
rect 88000 49476 88056 49478
rect 88080 49476 88136 49478
rect 89938 49240 89994 49296
rect 87104 48986 87160 48988
rect 87184 48986 87240 48988
rect 87264 48986 87320 48988
rect 87344 48986 87400 48988
rect 87104 48934 87150 48986
rect 87150 48934 87160 48986
rect 87184 48934 87214 48986
rect 87214 48934 87226 48986
rect 87226 48934 87240 48986
rect 87264 48934 87278 48986
rect 87278 48934 87290 48986
rect 87290 48934 87320 48986
rect 87344 48934 87354 48986
rect 87354 48934 87400 48986
rect 87104 48932 87160 48934
rect 87184 48932 87240 48934
rect 87264 48932 87320 48934
rect 87344 48932 87400 48934
rect 89938 48596 89940 48616
rect 89940 48596 89992 48616
rect 89992 48596 89994 48616
rect 89938 48560 89994 48596
rect 87840 48442 87896 48444
rect 87920 48442 87976 48444
rect 88000 48442 88056 48444
rect 88080 48442 88136 48444
rect 87840 48390 87886 48442
rect 87886 48390 87896 48442
rect 87920 48390 87950 48442
rect 87950 48390 87962 48442
rect 87962 48390 87976 48442
rect 88000 48390 88014 48442
rect 88014 48390 88026 48442
rect 88026 48390 88056 48442
rect 88080 48390 88090 48442
rect 88090 48390 88136 48442
rect 87840 48388 87896 48390
rect 87920 48388 87976 48390
rect 88000 48388 88056 48390
rect 88080 48388 88136 48390
rect 87104 47898 87160 47900
rect 87184 47898 87240 47900
rect 87264 47898 87320 47900
rect 87344 47898 87400 47900
rect 87104 47846 87150 47898
rect 87150 47846 87160 47898
rect 87184 47846 87214 47898
rect 87214 47846 87226 47898
rect 87226 47846 87240 47898
rect 87264 47846 87278 47898
rect 87278 47846 87290 47898
rect 87290 47846 87320 47898
rect 87344 47846 87354 47898
rect 87354 47846 87400 47898
rect 88558 47880 88614 47936
rect 87104 47844 87160 47846
rect 87184 47844 87240 47846
rect 87264 47844 87320 47846
rect 87344 47844 87400 47846
rect 87840 47354 87896 47356
rect 87920 47354 87976 47356
rect 88000 47354 88056 47356
rect 88080 47354 88136 47356
rect 87840 47302 87886 47354
rect 87886 47302 87896 47354
rect 87920 47302 87950 47354
rect 87950 47302 87962 47354
rect 87962 47302 87976 47354
rect 88000 47302 88014 47354
rect 88014 47302 88026 47354
rect 88026 47302 88056 47354
rect 88080 47302 88090 47354
rect 88090 47302 88136 47354
rect 87840 47300 87896 47302
rect 87920 47300 87976 47302
rect 88000 47300 88056 47302
rect 88080 47300 88136 47302
rect 84326 42984 84382 43040
rect 84326 41896 84382 41952
rect 84326 39720 84382 39776
rect 84326 37544 84382 37600
rect 84326 36456 84382 36512
rect 84326 34280 84382 34336
rect 84326 32104 84382 32160
rect 84326 31016 84382 31072
rect 84326 28840 84382 28896
rect 84326 26664 84382 26720
rect 84326 25576 84382 25632
rect 84326 23400 84382 23456
rect 84326 22312 84382 22368
rect 84326 21224 84382 21280
rect 84326 20136 84382 20192
rect 84326 16872 84382 16928
rect 84326 15784 84382 15840
rect 84326 14696 84382 14752
rect 9806 10616 9862 10672
rect 11122 10616 11178 10672
rect 12226 10480 12282 10536
rect 13330 10344 13386 10400
rect 46698 10344 46754 10400
rect 14434 10208 14490 10264
rect 12226 10072 12282 10128
rect 13330 10072 13386 10128
rect 12658 9936 12714 9992
rect 14682 9936 14738 9992
rect 15418 9936 15474 9992
rect 8426 8440 8482 8496
rect 6696 8186 6752 8188
rect 6776 8186 6832 8188
rect 6856 8186 6912 8188
rect 6936 8186 6992 8188
rect 6696 8134 6742 8186
rect 6742 8134 6752 8186
rect 6776 8134 6806 8186
rect 6806 8134 6818 8186
rect 6818 8134 6832 8186
rect 6856 8134 6870 8186
rect 6870 8134 6882 8186
rect 6882 8134 6912 8186
rect 6936 8134 6946 8186
rect 6946 8134 6992 8186
rect 6696 8132 6752 8134
rect 6776 8132 6832 8134
rect 6856 8132 6912 8134
rect 6936 8132 6992 8134
rect 5960 7642 6016 7644
rect 6040 7642 6096 7644
rect 6120 7642 6176 7644
rect 6200 7642 6256 7644
rect 5960 7590 6006 7642
rect 6006 7590 6016 7642
rect 6040 7590 6070 7642
rect 6070 7590 6082 7642
rect 6082 7590 6096 7642
rect 6120 7590 6134 7642
rect 6134 7590 6146 7642
rect 6146 7590 6176 7642
rect 6200 7590 6210 7642
rect 6210 7590 6256 7642
rect 5960 7588 6016 7590
rect 6040 7588 6096 7590
rect 6120 7588 6176 7590
rect 6200 7588 6256 7590
rect 6696 7098 6752 7100
rect 6776 7098 6832 7100
rect 6856 7098 6912 7100
rect 6936 7098 6992 7100
rect 6696 7046 6742 7098
rect 6742 7046 6752 7098
rect 6776 7046 6806 7098
rect 6806 7046 6818 7098
rect 6818 7046 6832 7098
rect 6856 7046 6870 7098
rect 6870 7046 6882 7098
rect 6882 7046 6912 7098
rect 6936 7046 6946 7098
rect 6946 7046 6992 7098
rect 6696 7044 6752 7046
rect 6776 7044 6832 7046
rect 6856 7044 6912 7046
rect 6936 7044 6992 7046
rect 18728 7642 18784 7644
rect 18808 7642 18864 7644
rect 18888 7642 18944 7644
rect 18968 7642 19024 7644
rect 18728 7590 18774 7642
rect 18774 7590 18784 7642
rect 18808 7590 18838 7642
rect 18838 7590 18850 7642
rect 18850 7590 18864 7642
rect 18888 7590 18902 7642
rect 18902 7590 18914 7642
rect 18914 7590 18944 7642
rect 18968 7590 18978 7642
rect 18978 7590 19024 7642
rect 18728 7588 18784 7590
rect 18808 7588 18864 7590
rect 18888 7588 18944 7590
rect 18968 7588 19024 7590
rect 18728 6554 18784 6556
rect 18808 6554 18864 6556
rect 18888 6554 18944 6556
rect 18968 6554 19024 6556
rect 18728 6502 18774 6554
rect 18774 6502 18784 6554
rect 18808 6502 18838 6554
rect 18838 6502 18850 6554
rect 18850 6502 18864 6554
rect 18888 6502 18902 6554
rect 18902 6502 18914 6554
rect 18914 6502 18944 6554
rect 18968 6502 18978 6554
rect 18978 6502 19024 6554
rect 18728 6500 18784 6502
rect 18808 6500 18864 6502
rect 18888 6500 18944 6502
rect 18968 6500 19024 6502
rect 18728 5466 18784 5468
rect 18808 5466 18864 5468
rect 18888 5466 18944 5468
rect 18968 5466 19024 5468
rect 18728 5414 18774 5466
rect 18774 5414 18784 5466
rect 18808 5414 18838 5466
rect 18838 5414 18850 5466
rect 18850 5414 18864 5466
rect 18888 5414 18902 5466
rect 18902 5414 18914 5466
rect 18914 5414 18944 5466
rect 18968 5414 18978 5466
rect 18978 5414 19024 5466
rect 18728 5412 18784 5414
rect 18808 5412 18864 5414
rect 18888 5412 18944 5414
rect 18968 5412 19024 5414
rect 19388 7098 19444 7100
rect 19468 7098 19524 7100
rect 19548 7098 19604 7100
rect 19628 7098 19684 7100
rect 19388 7046 19434 7098
rect 19434 7046 19444 7098
rect 19468 7046 19498 7098
rect 19498 7046 19510 7098
rect 19510 7046 19524 7098
rect 19548 7046 19562 7098
rect 19562 7046 19574 7098
rect 19574 7046 19604 7098
rect 19628 7046 19638 7098
rect 19638 7046 19684 7098
rect 19388 7044 19444 7046
rect 19468 7044 19524 7046
rect 19548 7044 19604 7046
rect 19628 7044 19684 7046
rect 19388 6010 19444 6012
rect 19468 6010 19524 6012
rect 19548 6010 19604 6012
rect 19628 6010 19684 6012
rect 19388 5958 19434 6010
rect 19434 5958 19444 6010
rect 19468 5958 19498 6010
rect 19498 5958 19510 6010
rect 19510 5958 19524 6010
rect 19548 5958 19562 6010
rect 19562 5958 19574 6010
rect 19574 5958 19604 6010
rect 19628 5958 19638 6010
rect 19638 5958 19684 6010
rect 19388 5956 19444 5958
rect 19468 5956 19524 5958
rect 19548 5956 19604 5958
rect 19628 5956 19684 5958
rect 87104 46810 87160 46812
rect 87184 46810 87240 46812
rect 87264 46810 87320 46812
rect 87344 46810 87400 46812
rect 87104 46758 87150 46810
rect 87150 46758 87160 46810
rect 87184 46758 87214 46810
rect 87214 46758 87226 46810
rect 87226 46758 87240 46810
rect 87264 46758 87278 46810
rect 87278 46758 87290 46810
rect 87290 46758 87320 46810
rect 87344 46758 87354 46810
rect 87354 46758 87400 46810
rect 87104 46756 87160 46758
rect 87184 46756 87240 46758
rect 87264 46756 87320 46758
rect 87344 46756 87400 46758
rect 88558 46520 88614 46576
rect 87840 46266 87896 46268
rect 87920 46266 87976 46268
rect 88000 46266 88056 46268
rect 88080 46266 88136 46268
rect 87840 46214 87886 46266
rect 87886 46214 87896 46266
rect 87920 46214 87950 46266
rect 87950 46214 87962 46266
rect 87962 46214 87976 46266
rect 88000 46214 88014 46266
rect 88014 46214 88026 46266
rect 88026 46214 88056 46266
rect 88080 46214 88090 46266
rect 88090 46214 88136 46266
rect 87840 46212 87896 46214
rect 87920 46212 87976 46214
rect 88000 46212 88056 46214
rect 88080 46212 88136 46214
rect 87104 45722 87160 45724
rect 87184 45722 87240 45724
rect 87264 45722 87320 45724
rect 87344 45722 87400 45724
rect 87104 45670 87150 45722
rect 87150 45670 87160 45722
rect 87184 45670 87214 45722
rect 87214 45670 87226 45722
rect 87226 45670 87240 45722
rect 87264 45670 87278 45722
rect 87278 45670 87290 45722
rect 87290 45670 87320 45722
rect 87344 45670 87354 45722
rect 87354 45670 87400 45722
rect 87104 45668 87160 45670
rect 87184 45668 87240 45670
rect 87264 45668 87320 45670
rect 87344 45668 87400 45670
rect 87840 45178 87896 45180
rect 87920 45178 87976 45180
rect 88000 45178 88056 45180
rect 88080 45178 88136 45180
rect 87840 45126 87886 45178
rect 87886 45126 87896 45178
rect 87920 45126 87950 45178
rect 87950 45126 87962 45178
rect 87962 45126 87976 45178
rect 88000 45126 88014 45178
rect 88014 45126 88026 45178
rect 88026 45126 88056 45178
rect 88080 45126 88090 45178
rect 88090 45126 88136 45178
rect 87840 45124 87896 45126
rect 87920 45124 87976 45126
rect 88000 45124 88056 45126
rect 88080 45124 88136 45126
rect 87104 44634 87160 44636
rect 87184 44634 87240 44636
rect 87264 44634 87320 44636
rect 87344 44634 87400 44636
rect 87104 44582 87150 44634
rect 87150 44582 87160 44634
rect 87184 44582 87214 44634
rect 87214 44582 87226 44634
rect 87226 44582 87240 44634
rect 87264 44582 87278 44634
rect 87278 44582 87290 44634
rect 87290 44582 87320 44634
rect 87344 44582 87354 44634
rect 87354 44582 87400 44634
rect 87104 44580 87160 44582
rect 87184 44580 87240 44582
rect 87264 44580 87320 44582
rect 87344 44580 87400 44582
rect 87840 44090 87896 44092
rect 87920 44090 87976 44092
rect 88000 44090 88056 44092
rect 88080 44090 88136 44092
rect 87840 44038 87886 44090
rect 87886 44038 87896 44090
rect 87920 44038 87950 44090
rect 87950 44038 87962 44090
rect 87962 44038 87976 44090
rect 88000 44038 88014 44090
rect 88014 44038 88026 44090
rect 88026 44038 88056 44090
rect 88080 44038 88090 44090
rect 88090 44038 88136 44090
rect 87840 44036 87896 44038
rect 87920 44036 87976 44038
rect 88000 44036 88056 44038
rect 88080 44036 88136 44038
rect 87104 43546 87160 43548
rect 87184 43546 87240 43548
rect 87264 43546 87320 43548
rect 87344 43546 87400 43548
rect 87104 43494 87150 43546
rect 87150 43494 87160 43546
rect 87184 43494 87214 43546
rect 87214 43494 87226 43546
rect 87226 43494 87240 43546
rect 87264 43494 87278 43546
rect 87278 43494 87290 43546
rect 87290 43494 87320 43546
rect 87344 43494 87354 43546
rect 87354 43494 87400 43546
rect 87104 43492 87160 43494
rect 87184 43492 87240 43494
rect 87264 43492 87320 43494
rect 87344 43492 87400 43494
rect 89938 43120 89994 43176
rect 87840 43002 87896 43004
rect 87920 43002 87976 43004
rect 88000 43002 88056 43004
rect 88080 43002 88136 43004
rect 87840 42950 87886 43002
rect 87886 42950 87896 43002
rect 87920 42950 87950 43002
rect 87950 42950 87962 43002
rect 87962 42950 87976 43002
rect 88000 42950 88014 43002
rect 88014 42950 88026 43002
rect 88026 42950 88056 43002
rect 88080 42950 88090 43002
rect 88090 42950 88136 43002
rect 87840 42948 87896 42950
rect 87920 42948 87976 42950
rect 88000 42948 88056 42950
rect 88080 42948 88136 42950
rect 87104 42458 87160 42460
rect 87184 42458 87240 42460
rect 87264 42458 87320 42460
rect 87344 42458 87400 42460
rect 87104 42406 87150 42458
rect 87150 42406 87160 42458
rect 87184 42406 87214 42458
rect 87214 42406 87226 42458
rect 87226 42406 87240 42458
rect 87264 42406 87278 42458
rect 87278 42406 87290 42458
rect 87290 42406 87320 42458
rect 87344 42406 87354 42458
rect 87354 42406 87400 42458
rect 87104 42404 87160 42406
rect 87184 42404 87240 42406
rect 87264 42404 87320 42406
rect 87344 42404 87400 42406
rect 87840 41914 87896 41916
rect 87920 41914 87976 41916
rect 88000 41914 88056 41916
rect 88080 41914 88136 41916
rect 87840 41862 87886 41914
rect 87886 41862 87896 41914
rect 87920 41862 87950 41914
rect 87950 41862 87962 41914
rect 87962 41862 87976 41914
rect 88000 41862 88014 41914
rect 88014 41862 88026 41914
rect 88026 41862 88056 41914
rect 88080 41862 88090 41914
rect 88090 41862 88136 41914
rect 87840 41860 87896 41862
rect 87920 41860 87976 41862
rect 88000 41860 88056 41862
rect 88080 41860 88136 41862
rect 88558 41760 88614 41816
rect 87104 41370 87160 41372
rect 87184 41370 87240 41372
rect 87264 41370 87320 41372
rect 87344 41370 87400 41372
rect 87104 41318 87150 41370
rect 87150 41318 87160 41370
rect 87184 41318 87214 41370
rect 87214 41318 87226 41370
rect 87226 41318 87240 41370
rect 87264 41318 87278 41370
rect 87278 41318 87290 41370
rect 87290 41318 87320 41370
rect 87344 41318 87354 41370
rect 87354 41318 87400 41370
rect 87104 41316 87160 41318
rect 87184 41316 87240 41318
rect 87264 41316 87320 41318
rect 87344 41316 87400 41318
rect 89938 41080 89994 41136
rect 87454 40808 87510 40864
rect 87840 40826 87896 40828
rect 87920 40826 87976 40828
rect 88000 40826 88056 40828
rect 88080 40826 88136 40828
rect 87840 40774 87886 40826
rect 87886 40774 87896 40826
rect 87920 40774 87950 40826
rect 87950 40774 87962 40826
rect 87962 40774 87976 40826
rect 88000 40774 88014 40826
rect 88014 40774 88026 40826
rect 88026 40774 88056 40826
rect 88080 40774 88090 40826
rect 88090 40774 88136 40826
rect 87840 40772 87896 40774
rect 87920 40772 87976 40774
rect 88000 40772 88056 40774
rect 88080 40772 88136 40774
rect 87104 40282 87160 40284
rect 87184 40282 87240 40284
rect 87264 40282 87320 40284
rect 87344 40282 87400 40284
rect 87104 40230 87150 40282
rect 87150 40230 87160 40282
rect 87184 40230 87214 40282
rect 87214 40230 87226 40282
rect 87226 40230 87240 40282
rect 87264 40230 87278 40282
rect 87278 40230 87290 40282
rect 87290 40230 87320 40282
rect 87344 40230 87354 40282
rect 87354 40230 87400 40282
rect 87104 40228 87160 40230
rect 87184 40228 87240 40230
rect 87264 40228 87320 40230
rect 87344 40228 87400 40230
rect 87840 39738 87896 39740
rect 87920 39738 87976 39740
rect 88000 39738 88056 39740
rect 88080 39738 88136 39740
rect 87840 39686 87886 39738
rect 87886 39686 87896 39738
rect 87920 39686 87950 39738
rect 87950 39686 87962 39738
rect 87962 39686 87976 39738
rect 88000 39686 88014 39738
rect 88014 39686 88026 39738
rect 88026 39686 88056 39738
rect 88080 39686 88090 39738
rect 88090 39686 88136 39738
rect 89938 39720 89994 39776
rect 87840 39684 87896 39686
rect 87920 39684 87976 39686
rect 88000 39684 88056 39686
rect 88080 39684 88136 39686
rect 87104 39194 87160 39196
rect 87184 39194 87240 39196
rect 87264 39194 87320 39196
rect 87344 39194 87400 39196
rect 87104 39142 87150 39194
rect 87150 39142 87160 39194
rect 87184 39142 87214 39194
rect 87214 39142 87226 39194
rect 87226 39142 87240 39194
rect 87264 39142 87278 39194
rect 87278 39142 87290 39194
rect 87290 39142 87320 39194
rect 87344 39142 87354 39194
rect 87354 39142 87400 39194
rect 87104 39140 87160 39142
rect 87184 39140 87240 39142
rect 87264 39140 87320 39142
rect 87344 39140 87400 39142
rect 87178 38632 87234 38688
rect 87840 38650 87896 38652
rect 87920 38650 87976 38652
rect 88000 38650 88056 38652
rect 88080 38650 88136 38652
rect 87840 38598 87886 38650
rect 87886 38598 87896 38650
rect 87920 38598 87950 38650
rect 87950 38598 87962 38650
rect 87962 38598 87976 38650
rect 88000 38598 88014 38650
rect 88014 38598 88026 38650
rect 88026 38598 88056 38650
rect 88080 38598 88090 38650
rect 88090 38598 88136 38650
rect 87840 38596 87896 38598
rect 87920 38596 87976 38598
rect 88000 38596 88056 38598
rect 88080 38596 88136 38598
rect 89294 38360 89350 38416
rect 87104 38106 87160 38108
rect 87184 38106 87240 38108
rect 87264 38106 87320 38108
rect 87344 38106 87400 38108
rect 87104 38054 87150 38106
rect 87150 38054 87160 38106
rect 87184 38054 87214 38106
rect 87214 38054 87226 38106
rect 87226 38054 87240 38106
rect 87264 38054 87278 38106
rect 87278 38054 87290 38106
rect 87290 38054 87320 38106
rect 87344 38054 87354 38106
rect 87354 38054 87400 38106
rect 87104 38052 87160 38054
rect 87184 38052 87240 38054
rect 87264 38052 87320 38054
rect 87344 38052 87400 38054
rect 89938 37716 89940 37736
rect 89940 37716 89992 37736
rect 89992 37716 89994 37736
rect 89938 37680 89994 37716
rect 87840 37562 87896 37564
rect 87920 37562 87976 37564
rect 88000 37562 88056 37564
rect 88080 37562 88136 37564
rect 87840 37510 87886 37562
rect 87886 37510 87896 37562
rect 87920 37510 87950 37562
rect 87950 37510 87962 37562
rect 87962 37510 87976 37562
rect 88000 37510 88014 37562
rect 88014 37510 88026 37562
rect 88026 37510 88056 37562
rect 88080 37510 88090 37562
rect 88090 37510 88136 37562
rect 87840 37508 87896 37510
rect 87920 37508 87976 37510
rect 88000 37508 88056 37510
rect 88080 37508 88136 37510
rect 87104 37018 87160 37020
rect 87184 37018 87240 37020
rect 87264 37018 87320 37020
rect 87344 37018 87400 37020
rect 87104 36966 87150 37018
rect 87150 36966 87160 37018
rect 87184 36966 87214 37018
rect 87214 36966 87226 37018
rect 87226 36966 87240 37018
rect 87264 36966 87278 37018
rect 87278 36966 87290 37018
rect 87290 36966 87320 37018
rect 87344 36966 87354 37018
rect 87354 36966 87400 37018
rect 87104 36964 87160 36966
rect 87184 36964 87240 36966
rect 87264 36964 87320 36966
rect 87344 36964 87400 36966
rect 87840 36474 87896 36476
rect 87920 36474 87976 36476
rect 88000 36474 88056 36476
rect 88080 36474 88136 36476
rect 87840 36422 87886 36474
rect 87886 36422 87896 36474
rect 87920 36422 87950 36474
rect 87950 36422 87962 36474
rect 87962 36422 87976 36474
rect 88000 36422 88014 36474
rect 88014 36422 88026 36474
rect 88026 36422 88056 36474
rect 88080 36422 88090 36474
rect 88090 36422 88136 36474
rect 87840 36420 87896 36422
rect 87920 36420 87976 36422
rect 88000 36420 88056 36422
rect 88080 36420 88136 36422
rect 89938 36320 89994 36376
rect 87104 35930 87160 35932
rect 87184 35930 87240 35932
rect 87264 35930 87320 35932
rect 87344 35930 87400 35932
rect 87104 35878 87150 35930
rect 87150 35878 87160 35930
rect 87184 35878 87214 35930
rect 87214 35878 87226 35930
rect 87226 35878 87240 35930
rect 87264 35878 87278 35930
rect 87278 35878 87290 35930
rect 87290 35878 87320 35930
rect 87344 35878 87354 35930
rect 87354 35878 87400 35930
rect 87104 35876 87160 35878
rect 87184 35876 87240 35878
rect 87264 35876 87320 35878
rect 87344 35876 87400 35878
rect 90122 35640 90178 35696
rect 87454 35368 87510 35424
rect 87840 35386 87896 35388
rect 87920 35386 87976 35388
rect 88000 35386 88056 35388
rect 88080 35386 88136 35388
rect 87840 35334 87886 35386
rect 87886 35334 87896 35386
rect 87920 35334 87950 35386
rect 87950 35334 87962 35386
rect 87962 35334 87976 35386
rect 88000 35334 88014 35386
rect 88014 35334 88026 35386
rect 88026 35334 88056 35386
rect 88080 35334 88090 35386
rect 88090 35334 88136 35386
rect 87840 35332 87896 35334
rect 87920 35332 87976 35334
rect 88000 35332 88056 35334
rect 88080 35332 88136 35334
rect 87104 34842 87160 34844
rect 87184 34842 87240 34844
rect 87264 34842 87320 34844
rect 87344 34842 87400 34844
rect 87104 34790 87150 34842
rect 87150 34790 87160 34842
rect 87184 34790 87214 34842
rect 87214 34790 87226 34842
rect 87226 34790 87240 34842
rect 87264 34790 87278 34842
rect 87278 34790 87290 34842
rect 87290 34790 87320 34842
rect 87344 34790 87354 34842
rect 87354 34790 87400 34842
rect 87104 34788 87160 34790
rect 87184 34788 87240 34790
rect 87264 34788 87320 34790
rect 87344 34788 87400 34790
rect 87840 34298 87896 34300
rect 87920 34298 87976 34300
rect 88000 34298 88056 34300
rect 88080 34298 88136 34300
rect 87840 34246 87886 34298
rect 87886 34246 87896 34298
rect 87920 34246 87950 34298
rect 87950 34246 87962 34298
rect 87962 34246 87976 34298
rect 88000 34246 88014 34298
rect 88014 34246 88026 34298
rect 88026 34246 88056 34298
rect 88080 34246 88090 34298
rect 88090 34246 88136 34298
rect 88558 34280 88614 34336
rect 87840 34244 87896 34246
rect 87920 34244 87976 34246
rect 88000 34244 88056 34246
rect 88080 34244 88136 34246
rect 87104 33754 87160 33756
rect 87184 33754 87240 33756
rect 87264 33754 87320 33756
rect 87344 33754 87400 33756
rect 87104 33702 87150 33754
rect 87150 33702 87160 33754
rect 87184 33702 87214 33754
rect 87214 33702 87226 33754
rect 87226 33702 87240 33754
rect 87264 33702 87278 33754
rect 87278 33702 87290 33754
rect 87290 33702 87320 33754
rect 87344 33702 87354 33754
rect 87354 33702 87400 33754
rect 87104 33700 87160 33702
rect 87184 33700 87240 33702
rect 87264 33700 87320 33702
rect 87344 33700 87400 33702
rect 87178 33192 87234 33248
rect 87840 33210 87896 33212
rect 87920 33210 87976 33212
rect 88000 33210 88056 33212
rect 88080 33210 88136 33212
rect 87840 33158 87886 33210
rect 87886 33158 87896 33210
rect 87920 33158 87950 33210
rect 87950 33158 87962 33210
rect 87962 33158 87976 33210
rect 88000 33158 88014 33210
rect 88014 33158 88026 33210
rect 88026 33158 88056 33210
rect 88080 33158 88090 33210
rect 88090 33158 88136 33210
rect 87840 33156 87896 33158
rect 87920 33156 87976 33158
rect 88000 33156 88056 33158
rect 88080 33156 88136 33158
rect 89938 32920 89994 32976
rect 87104 32666 87160 32668
rect 87184 32666 87240 32668
rect 87264 32666 87320 32668
rect 87344 32666 87400 32668
rect 87104 32614 87150 32666
rect 87150 32614 87160 32666
rect 87184 32614 87214 32666
rect 87214 32614 87226 32666
rect 87226 32614 87240 32666
rect 87264 32614 87278 32666
rect 87278 32614 87290 32666
rect 87290 32614 87320 32666
rect 87344 32614 87354 32666
rect 87354 32614 87400 32666
rect 87104 32612 87160 32614
rect 87184 32612 87240 32614
rect 87264 32612 87320 32614
rect 87344 32612 87400 32614
rect 89938 32276 89940 32296
rect 89940 32276 89992 32296
rect 89992 32276 89994 32296
rect 89938 32240 89994 32276
rect 87840 32122 87896 32124
rect 87920 32122 87976 32124
rect 88000 32122 88056 32124
rect 88080 32122 88136 32124
rect 87840 32070 87886 32122
rect 87886 32070 87896 32122
rect 87920 32070 87950 32122
rect 87950 32070 87962 32122
rect 87962 32070 87976 32122
rect 88000 32070 88014 32122
rect 88014 32070 88026 32122
rect 88026 32070 88056 32122
rect 88080 32070 88090 32122
rect 88090 32070 88136 32122
rect 87840 32068 87896 32070
rect 87920 32068 87976 32070
rect 88000 32068 88056 32070
rect 88080 32068 88136 32070
rect 87104 31578 87160 31580
rect 87184 31578 87240 31580
rect 87264 31578 87320 31580
rect 87344 31578 87400 31580
rect 87104 31526 87150 31578
rect 87150 31526 87160 31578
rect 87184 31526 87214 31578
rect 87214 31526 87226 31578
rect 87226 31526 87240 31578
rect 87264 31526 87278 31578
rect 87278 31526 87290 31578
rect 87290 31526 87320 31578
rect 87344 31526 87354 31578
rect 87354 31526 87400 31578
rect 87104 31524 87160 31526
rect 87184 31524 87240 31526
rect 87264 31524 87320 31526
rect 87344 31524 87400 31526
rect 87840 31034 87896 31036
rect 87920 31034 87976 31036
rect 88000 31034 88056 31036
rect 88080 31034 88136 31036
rect 87840 30982 87886 31034
rect 87886 30982 87896 31034
rect 87920 30982 87950 31034
rect 87950 30982 87962 31034
rect 87962 30982 87976 31034
rect 88000 30982 88014 31034
rect 88014 30982 88026 31034
rect 88026 30982 88056 31034
rect 88080 30982 88090 31034
rect 88090 30982 88136 31034
rect 87840 30980 87896 30982
rect 87920 30980 87976 30982
rect 88000 30980 88056 30982
rect 88080 30980 88136 30982
rect 88558 30880 88614 30936
rect 87104 30490 87160 30492
rect 87184 30490 87240 30492
rect 87264 30490 87320 30492
rect 87344 30490 87400 30492
rect 87104 30438 87150 30490
rect 87150 30438 87160 30490
rect 87184 30438 87214 30490
rect 87214 30438 87226 30490
rect 87226 30438 87240 30490
rect 87264 30438 87278 30490
rect 87278 30438 87290 30490
rect 87290 30438 87320 30490
rect 87344 30438 87354 30490
rect 87354 30438 87400 30490
rect 87104 30436 87160 30438
rect 87184 30436 87240 30438
rect 87264 30436 87320 30438
rect 87344 30436 87400 30438
rect 87454 30200 87510 30256
rect 89938 30200 89994 30256
rect 87840 29946 87896 29948
rect 87920 29946 87976 29948
rect 88000 29946 88056 29948
rect 88080 29946 88136 29948
rect 87840 29894 87886 29946
rect 87886 29894 87896 29946
rect 87920 29894 87950 29946
rect 87950 29894 87962 29946
rect 87962 29894 87976 29946
rect 88000 29894 88014 29946
rect 88014 29894 88026 29946
rect 88026 29894 88056 29946
rect 88080 29894 88090 29946
rect 88090 29894 88136 29946
rect 87840 29892 87896 29894
rect 87920 29892 87976 29894
rect 88000 29892 88056 29894
rect 88080 29892 88136 29894
rect 87104 29402 87160 29404
rect 87184 29402 87240 29404
rect 87264 29402 87320 29404
rect 87344 29402 87400 29404
rect 87104 29350 87150 29402
rect 87150 29350 87160 29402
rect 87184 29350 87214 29402
rect 87214 29350 87226 29402
rect 87226 29350 87240 29402
rect 87264 29350 87278 29402
rect 87278 29350 87290 29402
rect 87290 29350 87320 29402
rect 87344 29350 87354 29402
rect 87354 29350 87400 29402
rect 87104 29348 87160 29350
rect 87184 29348 87240 29350
rect 87264 29348 87320 29350
rect 87344 29348 87400 29350
rect 87840 28858 87896 28860
rect 87920 28858 87976 28860
rect 88000 28858 88056 28860
rect 88080 28858 88136 28860
rect 87840 28806 87886 28858
rect 87886 28806 87896 28858
rect 87920 28806 87950 28858
rect 87950 28806 87962 28858
rect 87962 28806 87976 28858
rect 88000 28806 88014 28858
rect 88014 28806 88026 28858
rect 88026 28806 88056 28858
rect 88080 28806 88090 28858
rect 88090 28806 88136 28858
rect 88558 28840 88614 28896
rect 87840 28804 87896 28806
rect 87920 28804 87976 28806
rect 88000 28804 88056 28806
rect 88080 28804 88136 28806
rect 87104 28314 87160 28316
rect 87184 28314 87240 28316
rect 87264 28314 87320 28316
rect 87344 28314 87400 28316
rect 87104 28262 87150 28314
rect 87150 28262 87160 28314
rect 87184 28262 87214 28314
rect 87214 28262 87226 28314
rect 87226 28262 87240 28314
rect 87264 28262 87278 28314
rect 87278 28262 87290 28314
rect 87290 28262 87320 28314
rect 87344 28262 87354 28314
rect 87354 28262 87400 28314
rect 87104 28260 87160 28262
rect 87184 28260 87240 28262
rect 87264 28260 87320 28262
rect 87344 28260 87400 28262
rect 87546 27752 87602 27808
rect 87840 27770 87896 27772
rect 87920 27770 87976 27772
rect 88000 27770 88056 27772
rect 88080 27770 88136 27772
rect 87840 27718 87886 27770
rect 87886 27718 87896 27770
rect 87920 27718 87950 27770
rect 87950 27718 87962 27770
rect 87962 27718 87976 27770
rect 88000 27718 88014 27770
rect 88014 27718 88026 27770
rect 88026 27718 88056 27770
rect 88080 27718 88090 27770
rect 88090 27718 88136 27770
rect 87840 27716 87896 27718
rect 87920 27716 87976 27718
rect 88000 27716 88056 27718
rect 88080 27716 88136 27718
rect 89938 27480 89994 27536
rect 87104 27226 87160 27228
rect 87184 27226 87240 27228
rect 87264 27226 87320 27228
rect 87344 27226 87400 27228
rect 87104 27174 87150 27226
rect 87150 27174 87160 27226
rect 87184 27174 87214 27226
rect 87214 27174 87226 27226
rect 87226 27174 87240 27226
rect 87264 27174 87278 27226
rect 87278 27174 87290 27226
rect 87290 27174 87320 27226
rect 87344 27174 87354 27226
rect 87354 27174 87400 27226
rect 87104 27172 87160 27174
rect 87184 27172 87240 27174
rect 87264 27172 87320 27174
rect 87344 27172 87400 27174
rect 89938 26820 89994 26856
rect 89938 26800 89940 26820
rect 89940 26800 89992 26820
rect 89992 26800 89994 26820
rect 87840 26682 87896 26684
rect 87920 26682 87976 26684
rect 88000 26682 88056 26684
rect 88080 26682 88136 26684
rect 87840 26630 87886 26682
rect 87886 26630 87896 26682
rect 87920 26630 87950 26682
rect 87950 26630 87962 26682
rect 87962 26630 87976 26682
rect 88000 26630 88014 26682
rect 88014 26630 88026 26682
rect 88026 26630 88056 26682
rect 88080 26630 88090 26682
rect 88090 26630 88136 26682
rect 87840 26628 87896 26630
rect 87920 26628 87976 26630
rect 88000 26628 88056 26630
rect 88080 26628 88136 26630
rect 87104 26138 87160 26140
rect 87184 26138 87240 26140
rect 87264 26138 87320 26140
rect 87344 26138 87400 26140
rect 87104 26086 87150 26138
rect 87150 26086 87160 26138
rect 87184 26086 87214 26138
rect 87214 26086 87226 26138
rect 87226 26086 87240 26138
rect 87264 26086 87278 26138
rect 87278 26086 87290 26138
rect 87290 26086 87320 26138
rect 87344 26086 87354 26138
rect 87354 26086 87400 26138
rect 87104 26084 87160 26086
rect 87184 26084 87240 26086
rect 87264 26084 87320 26086
rect 87344 26084 87400 26086
rect 87840 25594 87896 25596
rect 87920 25594 87976 25596
rect 88000 25594 88056 25596
rect 88080 25594 88136 25596
rect 87840 25542 87886 25594
rect 87886 25542 87896 25594
rect 87920 25542 87950 25594
rect 87950 25542 87962 25594
rect 87962 25542 87976 25594
rect 88000 25542 88014 25594
rect 88014 25542 88026 25594
rect 88026 25542 88056 25594
rect 88080 25542 88090 25594
rect 88090 25542 88136 25594
rect 87840 25540 87896 25542
rect 87920 25540 87976 25542
rect 88000 25540 88056 25542
rect 88080 25540 88136 25542
rect 89938 25440 89994 25496
rect 87104 25050 87160 25052
rect 87184 25050 87240 25052
rect 87264 25050 87320 25052
rect 87344 25050 87400 25052
rect 87104 24998 87150 25050
rect 87150 24998 87160 25050
rect 87184 24998 87214 25050
rect 87214 24998 87226 25050
rect 87226 24998 87240 25050
rect 87264 24998 87278 25050
rect 87278 24998 87290 25050
rect 87290 24998 87320 25050
rect 87344 24998 87354 25050
rect 87354 24998 87400 25050
rect 87104 24996 87160 24998
rect 87184 24996 87240 24998
rect 87264 24996 87320 24998
rect 87344 24996 87400 24998
rect 88374 24760 88430 24816
rect 89938 24760 89994 24816
rect 87840 24506 87896 24508
rect 87920 24506 87976 24508
rect 88000 24506 88056 24508
rect 88080 24506 88136 24508
rect 87840 24454 87886 24506
rect 87886 24454 87896 24506
rect 87920 24454 87950 24506
rect 87950 24454 87962 24506
rect 87962 24454 87976 24506
rect 88000 24454 88014 24506
rect 88014 24454 88026 24506
rect 88026 24454 88056 24506
rect 88080 24454 88090 24506
rect 88090 24454 88136 24506
rect 87840 24452 87896 24454
rect 87920 24452 87976 24454
rect 88000 24452 88056 24454
rect 88080 24452 88136 24454
rect 87104 23962 87160 23964
rect 87184 23962 87240 23964
rect 87264 23962 87320 23964
rect 87344 23962 87400 23964
rect 87104 23910 87150 23962
rect 87150 23910 87160 23962
rect 87184 23910 87214 23962
rect 87214 23910 87226 23962
rect 87226 23910 87240 23962
rect 87264 23910 87278 23962
rect 87278 23910 87290 23962
rect 87290 23910 87320 23962
rect 87344 23910 87354 23962
rect 87354 23910 87400 23962
rect 87104 23908 87160 23910
rect 87184 23908 87240 23910
rect 87264 23908 87320 23910
rect 87344 23908 87400 23910
rect 87840 23418 87896 23420
rect 87920 23418 87976 23420
rect 88000 23418 88056 23420
rect 88080 23418 88136 23420
rect 87840 23366 87886 23418
rect 87886 23366 87896 23418
rect 87920 23366 87950 23418
rect 87950 23366 87962 23418
rect 87962 23366 87976 23418
rect 88000 23366 88014 23418
rect 88014 23366 88026 23418
rect 88026 23366 88056 23418
rect 88080 23366 88090 23418
rect 88090 23366 88136 23418
rect 89938 23400 89994 23456
rect 87840 23364 87896 23366
rect 87920 23364 87976 23366
rect 88000 23364 88056 23366
rect 88080 23364 88136 23366
rect 87104 22874 87160 22876
rect 87184 22874 87240 22876
rect 87264 22874 87320 22876
rect 87344 22874 87400 22876
rect 87104 22822 87150 22874
rect 87150 22822 87160 22874
rect 87184 22822 87214 22874
rect 87214 22822 87226 22874
rect 87226 22822 87240 22874
rect 87264 22822 87278 22874
rect 87278 22822 87290 22874
rect 87290 22822 87320 22874
rect 87344 22822 87354 22874
rect 87354 22822 87400 22874
rect 87104 22820 87160 22822
rect 87184 22820 87240 22822
rect 87264 22820 87320 22822
rect 87344 22820 87400 22822
rect 87840 22330 87896 22332
rect 87920 22330 87976 22332
rect 88000 22330 88056 22332
rect 88080 22330 88136 22332
rect 87840 22278 87886 22330
rect 87886 22278 87896 22330
rect 87920 22278 87950 22330
rect 87950 22278 87962 22330
rect 87962 22278 87976 22330
rect 88000 22278 88014 22330
rect 88014 22278 88026 22330
rect 88026 22278 88056 22330
rect 88080 22278 88090 22330
rect 88090 22278 88136 22330
rect 87840 22276 87896 22278
rect 87920 22276 87976 22278
rect 88000 22276 88056 22278
rect 88080 22276 88136 22278
rect 89938 22040 89994 22096
rect 87104 21786 87160 21788
rect 87184 21786 87240 21788
rect 87264 21786 87320 21788
rect 87344 21786 87400 21788
rect 87104 21734 87150 21786
rect 87150 21734 87160 21786
rect 87184 21734 87214 21786
rect 87214 21734 87226 21786
rect 87226 21734 87240 21786
rect 87264 21734 87278 21786
rect 87278 21734 87290 21786
rect 87290 21734 87320 21786
rect 87344 21734 87354 21786
rect 87354 21734 87400 21786
rect 87104 21732 87160 21734
rect 87184 21732 87240 21734
rect 87264 21732 87320 21734
rect 87344 21732 87400 21734
rect 89938 21380 89994 21416
rect 89938 21360 89940 21380
rect 89940 21360 89992 21380
rect 89992 21360 89994 21380
rect 87840 21242 87896 21244
rect 87920 21242 87976 21244
rect 88000 21242 88056 21244
rect 88080 21242 88136 21244
rect 87840 21190 87886 21242
rect 87886 21190 87896 21242
rect 87920 21190 87950 21242
rect 87950 21190 87962 21242
rect 87962 21190 87976 21242
rect 88000 21190 88014 21242
rect 88014 21190 88026 21242
rect 88026 21190 88056 21242
rect 88080 21190 88090 21242
rect 88090 21190 88136 21242
rect 87840 21188 87896 21190
rect 87920 21188 87976 21190
rect 88000 21188 88056 21190
rect 88080 21188 88136 21190
rect 87104 20698 87160 20700
rect 87184 20698 87240 20700
rect 87264 20698 87320 20700
rect 87344 20698 87400 20700
rect 87104 20646 87150 20698
rect 87150 20646 87160 20698
rect 87184 20646 87214 20698
rect 87214 20646 87226 20698
rect 87226 20646 87240 20698
rect 87264 20646 87278 20698
rect 87278 20646 87290 20698
rect 87290 20646 87320 20698
rect 87344 20646 87354 20698
rect 87354 20646 87400 20698
rect 87104 20644 87160 20646
rect 87184 20644 87240 20646
rect 87264 20644 87320 20646
rect 87344 20644 87400 20646
rect 87840 20154 87896 20156
rect 87920 20154 87976 20156
rect 88000 20154 88056 20156
rect 88080 20154 88136 20156
rect 87840 20102 87886 20154
rect 87886 20102 87896 20154
rect 87920 20102 87950 20154
rect 87950 20102 87962 20154
rect 87962 20102 87976 20154
rect 88000 20102 88014 20154
rect 88014 20102 88026 20154
rect 88026 20102 88056 20154
rect 88080 20102 88090 20154
rect 88090 20102 88136 20154
rect 87840 20100 87896 20102
rect 87920 20100 87976 20102
rect 88000 20100 88056 20102
rect 88080 20100 88136 20102
rect 89938 20000 89994 20056
rect 87104 19610 87160 19612
rect 87184 19610 87240 19612
rect 87264 19610 87320 19612
rect 87344 19610 87400 19612
rect 87104 19558 87150 19610
rect 87150 19558 87160 19610
rect 87184 19558 87214 19610
rect 87214 19558 87226 19610
rect 87226 19558 87240 19610
rect 87264 19558 87278 19610
rect 87278 19558 87290 19610
rect 87290 19558 87320 19610
rect 87344 19558 87354 19610
rect 87354 19558 87400 19610
rect 87104 19556 87160 19558
rect 87184 19556 87240 19558
rect 87264 19556 87320 19558
rect 87344 19556 87400 19558
rect 88374 19320 88430 19376
rect 90030 19320 90086 19376
rect 87840 19066 87896 19068
rect 87920 19066 87976 19068
rect 88000 19066 88056 19068
rect 88080 19066 88136 19068
rect 87840 19014 87886 19066
rect 87886 19014 87896 19066
rect 87920 19014 87950 19066
rect 87950 19014 87962 19066
rect 87962 19014 87976 19066
rect 88000 19014 88014 19066
rect 88014 19014 88026 19066
rect 88026 19014 88056 19066
rect 88080 19014 88090 19066
rect 88090 19014 88136 19066
rect 87840 19012 87896 19014
rect 87920 19012 87976 19014
rect 88000 19012 88056 19014
rect 88080 19012 88136 19014
rect 87104 18522 87160 18524
rect 87184 18522 87240 18524
rect 87264 18522 87320 18524
rect 87344 18522 87400 18524
rect 87104 18470 87150 18522
rect 87150 18470 87160 18522
rect 87184 18470 87214 18522
rect 87214 18470 87226 18522
rect 87226 18470 87240 18522
rect 87264 18470 87278 18522
rect 87278 18470 87290 18522
rect 87290 18470 87320 18522
rect 87344 18470 87354 18522
rect 87354 18470 87400 18522
rect 87104 18468 87160 18470
rect 87184 18468 87240 18470
rect 87264 18468 87320 18470
rect 87344 18468 87400 18470
rect 88190 18096 88246 18152
rect 87840 17978 87896 17980
rect 87920 17978 87976 17980
rect 88000 17978 88056 17980
rect 88080 17978 88136 17980
rect 87840 17926 87886 17978
rect 87886 17926 87896 17978
rect 87920 17926 87950 17978
rect 87950 17926 87962 17978
rect 87962 17926 87976 17978
rect 88000 17926 88014 17978
rect 88014 17926 88026 17978
rect 88026 17926 88056 17978
rect 88080 17926 88090 17978
rect 88090 17926 88136 17978
rect 89938 17960 89994 18016
rect 87840 17924 87896 17926
rect 87920 17924 87976 17926
rect 88000 17924 88056 17926
rect 88080 17924 88136 17926
rect 87104 17434 87160 17436
rect 87184 17434 87240 17436
rect 87264 17434 87320 17436
rect 87344 17434 87400 17436
rect 87104 17382 87150 17434
rect 87150 17382 87160 17434
rect 87184 17382 87214 17434
rect 87214 17382 87226 17434
rect 87226 17382 87240 17434
rect 87264 17382 87278 17434
rect 87278 17382 87290 17434
rect 87290 17382 87320 17434
rect 87344 17382 87354 17434
rect 87354 17382 87400 17434
rect 87104 17380 87160 17382
rect 87184 17380 87240 17382
rect 87264 17380 87320 17382
rect 87344 17380 87400 17382
rect 87840 16890 87896 16892
rect 87920 16890 87976 16892
rect 88000 16890 88056 16892
rect 88080 16890 88136 16892
rect 87840 16838 87886 16890
rect 87886 16838 87896 16890
rect 87920 16838 87950 16890
rect 87950 16838 87962 16890
rect 87962 16838 87976 16890
rect 88000 16838 88014 16890
rect 88014 16838 88026 16890
rect 88026 16838 88056 16890
rect 88080 16838 88090 16890
rect 88090 16838 88136 16890
rect 87840 16836 87896 16838
rect 87920 16836 87976 16838
rect 88000 16836 88056 16838
rect 88080 16836 88136 16838
rect 89938 16600 89994 16656
rect 87104 16346 87160 16348
rect 87184 16346 87240 16348
rect 87264 16346 87320 16348
rect 87344 16346 87400 16348
rect 87104 16294 87150 16346
rect 87150 16294 87160 16346
rect 87184 16294 87214 16346
rect 87214 16294 87226 16346
rect 87226 16294 87240 16346
rect 87264 16294 87278 16346
rect 87278 16294 87290 16346
rect 87290 16294 87320 16346
rect 87344 16294 87354 16346
rect 87354 16294 87400 16346
rect 87104 16292 87160 16294
rect 87184 16292 87240 16294
rect 87264 16292 87320 16294
rect 87344 16292 87400 16294
rect 89938 15940 89994 15976
rect 89938 15920 89940 15940
rect 89940 15920 89992 15940
rect 89992 15920 89994 15940
rect 87840 15802 87896 15804
rect 87920 15802 87976 15804
rect 88000 15802 88056 15804
rect 88080 15802 88136 15804
rect 87840 15750 87886 15802
rect 87886 15750 87896 15802
rect 87920 15750 87950 15802
rect 87950 15750 87962 15802
rect 87962 15750 87976 15802
rect 88000 15750 88014 15802
rect 88014 15750 88026 15802
rect 88026 15750 88056 15802
rect 88080 15750 88090 15802
rect 88090 15750 88136 15802
rect 87840 15748 87896 15750
rect 87920 15748 87976 15750
rect 88000 15748 88056 15750
rect 88080 15748 88136 15750
rect 87104 15258 87160 15260
rect 87184 15258 87240 15260
rect 87264 15258 87320 15260
rect 87344 15258 87400 15260
rect 87104 15206 87150 15258
rect 87150 15206 87160 15258
rect 87184 15206 87214 15258
rect 87214 15206 87226 15258
rect 87226 15206 87240 15258
rect 87264 15206 87278 15258
rect 87278 15206 87290 15258
rect 87290 15206 87320 15258
rect 87344 15206 87354 15258
rect 87354 15206 87400 15258
rect 87104 15204 87160 15206
rect 87184 15204 87240 15206
rect 87264 15204 87320 15206
rect 87344 15204 87400 15206
rect 87840 14714 87896 14716
rect 87920 14714 87976 14716
rect 88000 14714 88056 14716
rect 88080 14714 88136 14716
rect 87840 14662 87886 14714
rect 87886 14662 87896 14714
rect 87920 14662 87950 14714
rect 87950 14662 87962 14714
rect 87962 14662 87976 14714
rect 88000 14662 88014 14714
rect 88014 14662 88026 14714
rect 88026 14662 88056 14714
rect 88080 14662 88090 14714
rect 88090 14662 88136 14714
rect 87840 14660 87896 14662
rect 87920 14660 87976 14662
rect 88000 14660 88056 14662
rect 88080 14660 88136 14662
rect 89938 14560 89994 14616
rect 87104 14170 87160 14172
rect 87184 14170 87240 14172
rect 87264 14170 87320 14172
rect 87344 14170 87400 14172
rect 87104 14118 87150 14170
rect 87150 14118 87160 14170
rect 87184 14118 87214 14170
rect 87214 14118 87226 14170
rect 87226 14118 87240 14170
rect 87264 14118 87278 14170
rect 87278 14118 87290 14170
rect 87290 14118 87320 14170
rect 87344 14118 87354 14170
rect 87354 14118 87400 14170
rect 87104 14116 87160 14118
rect 87184 14116 87240 14118
rect 87264 14116 87320 14118
rect 87344 14116 87400 14118
rect 88374 13880 88430 13936
rect 89938 13880 89994 13936
rect 87840 13626 87896 13628
rect 87920 13626 87976 13628
rect 88000 13626 88056 13628
rect 88080 13626 88136 13628
rect 87840 13574 87886 13626
rect 87886 13574 87896 13626
rect 87920 13574 87950 13626
rect 87950 13574 87962 13626
rect 87962 13574 87976 13626
rect 88000 13574 88014 13626
rect 88014 13574 88026 13626
rect 88026 13574 88056 13626
rect 88080 13574 88090 13626
rect 88090 13574 88136 13626
rect 87840 13572 87896 13574
rect 87920 13572 87976 13574
rect 88000 13572 88056 13574
rect 88080 13572 88136 13574
rect 87104 13082 87160 13084
rect 87184 13082 87240 13084
rect 87264 13082 87320 13084
rect 87344 13082 87400 13084
rect 87104 13030 87150 13082
rect 87150 13030 87160 13082
rect 87184 13030 87214 13082
rect 87214 13030 87226 13082
rect 87226 13030 87240 13082
rect 87264 13030 87278 13082
rect 87278 13030 87290 13082
rect 87290 13030 87320 13082
rect 87344 13030 87354 13082
rect 87354 13030 87400 13082
rect 87104 13028 87160 13030
rect 87184 13028 87240 13030
rect 87264 13028 87320 13030
rect 87344 13028 87400 13030
rect 87840 12538 87896 12540
rect 87920 12538 87976 12540
rect 88000 12538 88056 12540
rect 88080 12538 88136 12540
rect 87840 12486 87886 12538
rect 87886 12486 87896 12538
rect 87920 12486 87950 12538
rect 87950 12486 87962 12538
rect 87962 12486 87976 12538
rect 88000 12486 88014 12538
rect 88014 12486 88026 12538
rect 88026 12486 88056 12538
rect 88080 12486 88090 12538
rect 88090 12486 88136 12538
rect 87840 12484 87896 12486
rect 87920 12484 87976 12486
rect 88000 12484 88056 12486
rect 88080 12484 88136 12486
rect 87104 11994 87160 11996
rect 87184 11994 87240 11996
rect 87264 11994 87320 11996
rect 87344 11994 87400 11996
rect 87104 11942 87150 11994
rect 87150 11942 87160 11994
rect 87184 11942 87214 11994
rect 87214 11942 87226 11994
rect 87226 11942 87240 11994
rect 87264 11942 87278 11994
rect 87278 11942 87290 11994
rect 87290 11942 87320 11994
rect 87344 11942 87354 11994
rect 87354 11942 87400 11994
rect 87104 11940 87160 11942
rect 87184 11940 87240 11942
rect 87264 11940 87320 11942
rect 87344 11940 87400 11942
rect 87840 11450 87896 11452
rect 87920 11450 87976 11452
rect 88000 11450 88056 11452
rect 88080 11450 88136 11452
rect 87840 11398 87886 11450
rect 87886 11398 87896 11450
rect 87920 11398 87950 11450
rect 87950 11398 87962 11450
rect 87962 11398 87976 11450
rect 88000 11398 88014 11450
rect 88014 11398 88026 11450
rect 88026 11398 88056 11450
rect 88080 11398 88090 11450
rect 88090 11398 88136 11450
rect 87840 11396 87896 11398
rect 87920 11396 87976 11398
rect 88000 11396 88056 11398
rect 88080 11396 88136 11398
rect 87104 10906 87160 10908
rect 87184 10906 87240 10908
rect 87264 10906 87320 10908
rect 87344 10906 87400 10908
rect 87104 10854 87150 10906
rect 87150 10854 87160 10906
rect 87184 10854 87214 10906
rect 87214 10854 87226 10906
rect 87226 10854 87240 10906
rect 87264 10854 87278 10906
rect 87278 10854 87290 10906
rect 87290 10854 87320 10906
rect 87344 10854 87354 10906
rect 87354 10854 87400 10906
rect 87104 10852 87160 10854
rect 87184 10852 87240 10854
rect 87264 10852 87320 10854
rect 87344 10852 87400 10854
rect 87840 10362 87896 10364
rect 87920 10362 87976 10364
rect 88000 10362 88056 10364
rect 88080 10362 88136 10364
rect 87840 10310 87886 10362
rect 87886 10310 87896 10362
rect 87920 10310 87950 10362
rect 87950 10310 87962 10362
rect 87962 10310 87976 10362
rect 88000 10310 88014 10362
rect 88014 10310 88026 10362
rect 88026 10310 88056 10362
rect 88080 10310 88090 10362
rect 88090 10310 88136 10362
rect 87840 10308 87896 10310
rect 87920 10308 87976 10310
rect 88000 10308 88056 10310
rect 88080 10308 88136 10310
rect 84418 10208 84474 10264
rect 46698 9936 46754 9992
rect 49090 9936 49146 9992
rect 37728 7642 37784 7644
rect 37808 7642 37864 7644
rect 37888 7642 37944 7644
rect 37968 7642 38024 7644
rect 37728 7590 37774 7642
rect 37774 7590 37784 7642
rect 37808 7590 37838 7642
rect 37838 7590 37850 7642
rect 37850 7590 37864 7642
rect 37888 7590 37902 7642
rect 37902 7590 37914 7642
rect 37914 7590 37944 7642
rect 37968 7590 37978 7642
rect 37978 7590 38024 7642
rect 37728 7588 37784 7590
rect 37808 7588 37864 7590
rect 37888 7588 37944 7590
rect 37968 7588 38024 7590
rect 38388 7098 38444 7100
rect 38468 7098 38524 7100
rect 38548 7098 38604 7100
rect 38628 7098 38684 7100
rect 38388 7046 38434 7098
rect 38434 7046 38444 7098
rect 38468 7046 38498 7098
rect 38498 7046 38510 7098
rect 38510 7046 38524 7098
rect 38548 7046 38562 7098
rect 38562 7046 38574 7098
rect 38574 7046 38604 7098
rect 38628 7046 38638 7098
rect 38638 7046 38684 7098
rect 38388 7044 38444 7046
rect 38468 7044 38524 7046
rect 38548 7044 38604 7046
rect 38628 7044 38684 7046
rect 37728 6554 37784 6556
rect 37808 6554 37864 6556
rect 37888 6554 37944 6556
rect 37968 6554 38024 6556
rect 37728 6502 37774 6554
rect 37774 6502 37784 6554
rect 37808 6502 37838 6554
rect 37838 6502 37850 6554
rect 37850 6502 37864 6554
rect 37888 6502 37902 6554
rect 37902 6502 37914 6554
rect 37914 6502 37944 6554
rect 37968 6502 37978 6554
rect 37978 6502 38024 6554
rect 37728 6500 37784 6502
rect 37808 6500 37864 6502
rect 37888 6500 37944 6502
rect 37968 6500 38024 6502
rect 38388 6010 38444 6012
rect 38468 6010 38524 6012
rect 38548 6010 38604 6012
rect 38628 6010 38684 6012
rect 38388 5958 38434 6010
rect 38434 5958 38444 6010
rect 38468 5958 38498 6010
rect 38498 5958 38510 6010
rect 38510 5958 38524 6010
rect 38548 5958 38562 6010
rect 38562 5958 38574 6010
rect 38574 5958 38604 6010
rect 38628 5958 38638 6010
rect 38638 5958 38684 6010
rect 38388 5956 38444 5958
rect 38468 5956 38524 5958
rect 38548 5956 38604 5958
rect 38628 5956 38684 5958
rect 37728 5466 37784 5468
rect 37808 5466 37864 5468
rect 37888 5466 37944 5468
rect 37968 5466 38024 5468
rect 37728 5414 37774 5466
rect 37774 5414 37784 5466
rect 37808 5414 37838 5466
rect 37838 5414 37850 5466
rect 37850 5414 37864 5466
rect 37888 5414 37902 5466
rect 37902 5414 37914 5466
rect 37914 5414 37944 5466
rect 37968 5414 37978 5466
rect 37978 5414 38024 5466
rect 37728 5412 37784 5414
rect 37808 5412 37864 5414
rect 37888 5412 37944 5414
rect 37968 5412 38024 5414
rect 50194 9936 50250 9992
rect 51574 9936 51630 9992
rect 48078 8440 48134 8496
rect 19388 4922 19444 4924
rect 19468 4922 19524 4924
rect 19548 4922 19604 4924
rect 19628 4922 19684 4924
rect 19388 4870 19434 4922
rect 19434 4870 19444 4922
rect 19468 4870 19498 4922
rect 19498 4870 19510 4922
rect 19510 4870 19524 4922
rect 19548 4870 19562 4922
rect 19562 4870 19574 4922
rect 19574 4870 19604 4922
rect 19628 4870 19638 4922
rect 19638 4870 19684 4922
rect 19388 4868 19444 4870
rect 19468 4868 19524 4870
rect 19548 4868 19604 4870
rect 19628 4868 19684 4870
rect 56728 7642 56784 7644
rect 56808 7642 56864 7644
rect 56888 7642 56944 7644
rect 56968 7642 57024 7644
rect 56728 7590 56774 7642
rect 56774 7590 56784 7642
rect 56808 7590 56838 7642
rect 56838 7590 56850 7642
rect 56850 7590 56864 7642
rect 56888 7590 56902 7642
rect 56902 7590 56914 7642
rect 56914 7590 56944 7642
rect 56968 7590 56978 7642
rect 56978 7590 57024 7642
rect 56728 7588 56784 7590
rect 56808 7588 56864 7590
rect 56888 7588 56944 7590
rect 56968 7588 57024 7590
rect 56728 6554 56784 6556
rect 56808 6554 56864 6556
rect 56888 6554 56944 6556
rect 56968 6554 57024 6556
rect 56728 6502 56774 6554
rect 56774 6502 56784 6554
rect 56808 6502 56838 6554
rect 56838 6502 56850 6554
rect 56850 6502 56864 6554
rect 56888 6502 56902 6554
rect 56902 6502 56914 6554
rect 56914 6502 56944 6554
rect 56968 6502 56978 6554
rect 56978 6502 57024 6554
rect 56728 6500 56784 6502
rect 56808 6500 56864 6502
rect 56888 6500 56944 6502
rect 56968 6500 57024 6502
rect 56728 5466 56784 5468
rect 56808 5466 56864 5468
rect 56888 5466 56944 5468
rect 56968 5466 57024 5468
rect 56728 5414 56774 5466
rect 56774 5414 56784 5466
rect 56808 5414 56838 5466
rect 56838 5414 56850 5466
rect 56850 5414 56864 5466
rect 56888 5414 56902 5466
rect 56902 5414 56914 5466
rect 56914 5414 56944 5466
rect 56968 5414 56978 5466
rect 56978 5414 57024 5466
rect 56728 5412 56784 5414
rect 56808 5412 56864 5414
rect 56888 5412 56944 5414
rect 56968 5412 57024 5414
rect 57388 7098 57444 7100
rect 57468 7098 57524 7100
rect 57548 7098 57604 7100
rect 57628 7098 57684 7100
rect 57388 7046 57434 7098
rect 57434 7046 57444 7098
rect 57468 7046 57498 7098
rect 57498 7046 57510 7098
rect 57510 7046 57524 7098
rect 57548 7046 57562 7098
rect 57562 7046 57574 7098
rect 57574 7046 57604 7098
rect 57628 7046 57638 7098
rect 57638 7046 57684 7098
rect 57388 7044 57444 7046
rect 57468 7044 57524 7046
rect 57548 7044 57604 7046
rect 57628 7044 57684 7046
rect 57388 6010 57444 6012
rect 57468 6010 57524 6012
rect 57548 6010 57604 6012
rect 57628 6010 57684 6012
rect 57388 5958 57434 6010
rect 57434 5958 57444 6010
rect 57468 5958 57498 6010
rect 57498 5958 57510 6010
rect 57510 5958 57524 6010
rect 57548 5958 57562 6010
rect 57562 5958 57574 6010
rect 57574 5958 57604 6010
rect 57628 5958 57638 6010
rect 57638 5958 57684 6010
rect 57388 5956 57444 5958
rect 57468 5956 57524 5958
rect 57548 5956 57604 5958
rect 57628 5956 57684 5958
rect 75728 7642 75784 7644
rect 75808 7642 75864 7644
rect 75888 7642 75944 7644
rect 75968 7642 76024 7644
rect 75728 7590 75774 7642
rect 75774 7590 75784 7642
rect 75808 7590 75838 7642
rect 75838 7590 75850 7642
rect 75850 7590 75864 7642
rect 75888 7590 75902 7642
rect 75902 7590 75914 7642
rect 75914 7590 75944 7642
rect 75968 7590 75978 7642
rect 75978 7590 76024 7642
rect 75728 7588 75784 7590
rect 75808 7588 75864 7590
rect 75888 7588 75944 7590
rect 75968 7588 76024 7590
rect 76388 7098 76444 7100
rect 76468 7098 76524 7100
rect 76548 7098 76604 7100
rect 76628 7098 76684 7100
rect 76388 7046 76434 7098
rect 76434 7046 76444 7098
rect 76468 7046 76498 7098
rect 76498 7046 76510 7098
rect 76510 7046 76524 7098
rect 76548 7046 76562 7098
rect 76562 7046 76574 7098
rect 76574 7046 76604 7098
rect 76628 7046 76638 7098
rect 76638 7046 76684 7098
rect 76388 7044 76444 7046
rect 76468 7044 76524 7046
rect 76548 7044 76604 7046
rect 76628 7044 76684 7046
rect 75728 6554 75784 6556
rect 75808 6554 75864 6556
rect 75888 6554 75944 6556
rect 75968 6554 76024 6556
rect 75728 6502 75774 6554
rect 75774 6502 75784 6554
rect 75808 6502 75838 6554
rect 75838 6502 75850 6554
rect 75850 6502 75864 6554
rect 75888 6502 75902 6554
rect 75902 6502 75914 6554
rect 75914 6502 75944 6554
rect 75968 6502 75978 6554
rect 75978 6502 76024 6554
rect 75728 6500 75784 6502
rect 75808 6500 75864 6502
rect 75888 6500 75944 6502
rect 75968 6500 76024 6502
rect 76388 6010 76444 6012
rect 76468 6010 76524 6012
rect 76548 6010 76604 6012
rect 76628 6010 76684 6012
rect 76388 5958 76434 6010
rect 76434 5958 76444 6010
rect 76468 5958 76498 6010
rect 76498 5958 76510 6010
rect 76510 5958 76524 6010
rect 76548 5958 76562 6010
rect 76562 5958 76574 6010
rect 76574 5958 76604 6010
rect 76628 5958 76638 6010
rect 76638 5958 76684 6010
rect 76388 5956 76444 5958
rect 76468 5956 76524 5958
rect 76548 5956 76604 5958
rect 76628 5956 76684 5958
rect 75728 5466 75784 5468
rect 75808 5466 75864 5468
rect 75888 5466 75944 5468
rect 75968 5466 76024 5468
rect 75728 5414 75774 5466
rect 75774 5414 75784 5466
rect 75808 5414 75838 5466
rect 75838 5414 75850 5466
rect 75850 5414 75864 5466
rect 75888 5414 75902 5466
rect 75902 5414 75914 5466
rect 75914 5414 75944 5466
rect 75968 5414 75978 5466
rect 75978 5414 76024 5466
rect 75728 5412 75784 5414
rect 75808 5412 75864 5414
rect 75888 5412 75944 5414
rect 75968 5412 76024 5414
rect 38388 4922 38444 4924
rect 38468 4922 38524 4924
rect 38548 4922 38604 4924
rect 38628 4922 38684 4924
rect 38388 4870 38434 4922
rect 38434 4870 38444 4922
rect 38468 4870 38498 4922
rect 38498 4870 38510 4922
rect 38510 4870 38524 4922
rect 38548 4870 38562 4922
rect 38562 4870 38574 4922
rect 38574 4870 38604 4922
rect 38628 4870 38638 4922
rect 38638 4870 38684 4922
rect 38388 4868 38444 4870
rect 38468 4868 38524 4870
rect 38548 4868 38604 4870
rect 38628 4868 38684 4870
rect 57388 4922 57444 4924
rect 57468 4922 57524 4924
rect 57548 4922 57604 4924
rect 57628 4922 57684 4924
rect 57388 4870 57434 4922
rect 57434 4870 57444 4922
rect 57468 4870 57498 4922
rect 57498 4870 57510 4922
rect 57510 4870 57524 4922
rect 57548 4870 57562 4922
rect 57562 4870 57574 4922
rect 57574 4870 57604 4922
rect 57628 4870 57638 4922
rect 57638 4870 57684 4922
rect 57388 4868 57444 4870
rect 57468 4868 57524 4870
rect 57548 4868 57604 4870
rect 57628 4868 57684 4870
rect 76388 4922 76444 4924
rect 76468 4922 76524 4924
rect 76548 4922 76604 4924
rect 76628 4922 76684 4924
rect 76388 4870 76434 4922
rect 76434 4870 76444 4922
rect 76468 4870 76498 4922
rect 76498 4870 76510 4922
rect 76510 4870 76524 4922
rect 76548 4870 76562 4922
rect 76562 4870 76574 4922
rect 76574 4870 76604 4922
rect 76628 4870 76638 4922
rect 76638 4870 76684 4922
rect 76388 4868 76444 4870
rect 76468 4868 76524 4870
rect 76548 4868 76604 4870
rect 76628 4868 76684 4870
rect 87104 9818 87160 9820
rect 87184 9818 87240 9820
rect 87264 9818 87320 9820
rect 87344 9818 87400 9820
rect 87104 9766 87150 9818
rect 87150 9766 87160 9818
rect 87184 9766 87214 9818
rect 87214 9766 87226 9818
rect 87226 9766 87240 9818
rect 87264 9766 87278 9818
rect 87278 9766 87290 9818
rect 87290 9766 87320 9818
rect 87344 9766 87354 9818
rect 87354 9766 87400 9818
rect 87104 9764 87160 9766
rect 87184 9764 87240 9766
rect 87264 9764 87320 9766
rect 87344 9764 87400 9766
rect 87840 9274 87896 9276
rect 87920 9274 87976 9276
rect 88000 9274 88056 9276
rect 88080 9274 88136 9276
rect 87840 9222 87886 9274
rect 87886 9222 87896 9274
rect 87920 9222 87950 9274
rect 87950 9222 87962 9274
rect 87962 9222 87976 9274
rect 88000 9222 88014 9274
rect 88014 9222 88026 9274
rect 88026 9222 88056 9274
rect 88080 9222 88090 9274
rect 88090 9222 88136 9274
rect 87840 9220 87896 9222
rect 87920 9220 87976 9222
rect 88000 9220 88056 9222
rect 88080 9220 88136 9222
rect 87104 8730 87160 8732
rect 87184 8730 87240 8732
rect 87264 8730 87320 8732
rect 87344 8730 87400 8732
rect 87104 8678 87150 8730
rect 87150 8678 87160 8730
rect 87184 8678 87214 8730
rect 87214 8678 87226 8730
rect 87226 8678 87240 8730
rect 87264 8678 87278 8730
rect 87278 8678 87290 8730
rect 87290 8678 87320 8730
rect 87344 8678 87354 8730
rect 87354 8678 87400 8730
rect 87104 8676 87160 8678
rect 87184 8676 87240 8678
rect 87264 8676 87320 8678
rect 87344 8676 87400 8678
rect 87840 8186 87896 8188
rect 87920 8186 87976 8188
rect 88000 8186 88056 8188
rect 88080 8186 88136 8188
rect 87840 8134 87886 8186
rect 87886 8134 87896 8186
rect 87920 8134 87950 8186
rect 87950 8134 87962 8186
rect 87962 8134 87976 8186
rect 88000 8134 88014 8186
rect 88014 8134 88026 8186
rect 88026 8134 88056 8186
rect 88080 8134 88090 8186
rect 88090 8134 88136 8186
rect 87840 8132 87896 8134
rect 87920 8132 87976 8134
rect 88000 8132 88056 8134
rect 88080 8132 88136 8134
rect 87104 7642 87160 7644
rect 87184 7642 87240 7644
rect 87264 7642 87320 7644
rect 87344 7642 87400 7644
rect 87104 7590 87150 7642
rect 87150 7590 87160 7642
rect 87184 7590 87214 7642
rect 87214 7590 87226 7642
rect 87226 7590 87240 7642
rect 87264 7590 87278 7642
rect 87278 7590 87290 7642
rect 87290 7590 87320 7642
rect 87344 7590 87354 7642
rect 87354 7590 87400 7642
rect 87104 7588 87160 7590
rect 87184 7588 87240 7590
rect 87264 7588 87320 7590
rect 87344 7588 87400 7590
rect 87840 7098 87896 7100
rect 87920 7098 87976 7100
rect 88000 7098 88056 7100
rect 88080 7098 88136 7100
rect 87840 7046 87886 7098
rect 87886 7046 87896 7098
rect 87920 7046 87950 7098
rect 87950 7046 87962 7098
rect 87962 7046 87976 7098
rect 88000 7046 88014 7098
rect 88014 7046 88026 7098
rect 88026 7046 88056 7098
rect 88080 7046 88090 7098
rect 88090 7046 88136 7098
rect 87840 7044 87896 7046
rect 87920 7044 87976 7046
rect 88000 7044 88056 7046
rect 88080 7044 88136 7046
<< metal3 >>
rect 18718 89248 19034 89249
rect 18718 89184 18724 89248
rect 18788 89184 18804 89248
rect 18868 89184 18884 89248
rect 18948 89184 18964 89248
rect 19028 89184 19034 89248
rect 18718 89183 19034 89184
rect 37718 89248 38034 89249
rect 37718 89184 37724 89248
rect 37788 89184 37804 89248
rect 37868 89184 37884 89248
rect 37948 89184 37964 89248
rect 38028 89184 38034 89248
rect 37718 89183 38034 89184
rect 56718 89248 57034 89249
rect 56718 89184 56724 89248
rect 56788 89184 56804 89248
rect 56868 89184 56884 89248
rect 56948 89184 56964 89248
rect 57028 89184 57034 89248
rect 56718 89183 57034 89184
rect 75718 89248 76034 89249
rect 75718 89184 75724 89248
rect 75788 89184 75804 89248
rect 75868 89184 75884 89248
rect 75948 89184 75964 89248
rect 76028 89184 76034 89248
rect 75718 89183 76034 89184
rect 19378 88704 19694 88705
rect 19378 88640 19384 88704
rect 19448 88640 19464 88704
rect 19528 88640 19544 88704
rect 19608 88640 19624 88704
rect 19688 88640 19694 88704
rect 19378 88639 19694 88640
rect 38378 88704 38694 88705
rect 38378 88640 38384 88704
rect 38448 88640 38464 88704
rect 38528 88640 38544 88704
rect 38608 88640 38624 88704
rect 38688 88640 38694 88704
rect 38378 88639 38694 88640
rect 57378 88704 57694 88705
rect 57378 88640 57384 88704
rect 57448 88640 57464 88704
rect 57528 88640 57544 88704
rect 57608 88640 57624 88704
rect 57688 88640 57694 88704
rect 57378 88639 57694 88640
rect 76378 88704 76694 88705
rect 76378 88640 76384 88704
rect 76448 88640 76464 88704
rect 76528 88640 76544 88704
rect 76608 88640 76624 88704
rect 76688 88640 76694 88704
rect 76378 88639 76694 88640
rect 18718 88160 19034 88161
rect 18718 88096 18724 88160
rect 18788 88096 18804 88160
rect 18868 88096 18884 88160
rect 18948 88096 18964 88160
rect 19028 88096 19034 88160
rect 18718 88095 19034 88096
rect 37718 88160 38034 88161
rect 37718 88096 37724 88160
rect 37788 88096 37804 88160
rect 37868 88096 37884 88160
rect 37948 88096 37964 88160
rect 38028 88096 38034 88160
rect 37718 88095 38034 88096
rect 56718 88160 57034 88161
rect 56718 88096 56724 88160
rect 56788 88096 56804 88160
rect 56868 88096 56884 88160
rect 56948 88096 56964 88160
rect 57028 88096 57034 88160
rect 56718 88095 57034 88096
rect 75718 88160 76034 88161
rect 75718 88096 75724 88160
rect 75788 88096 75804 88160
rect 75868 88096 75884 88160
rect 75948 88096 75964 88160
rect 76028 88096 76034 88160
rect 75718 88095 76034 88096
rect 19378 87616 19694 87617
rect 19378 87552 19384 87616
rect 19448 87552 19464 87616
rect 19528 87552 19544 87616
rect 19608 87552 19624 87616
rect 19688 87552 19694 87616
rect 19378 87551 19694 87552
rect 38378 87616 38694 87617
rect 38378 87552 38384 87616
rect 38448 87552 38464 87616
rect 38528 87552 38544 87616
rect 38608 87552 38624 87616
rect 38688 87552 38694 87616
rect 38378 87551 38694 87552
rect 57378 87616 57694 87617
rect 57378 87552 57384 87616
rect 57448 87552 57464 87616
rect 57528 87552 57544 87616
rect 57608 87552 57624 87616
rect 57688 87552 57694 87616
rect 57378 87551 57694 87552
rect 76378 87616 76694 87617
rect 76378 87552 76384 87616
rect 76448 87552 76464 87616
rect 76528 87552 76544 87616
rect 76608 87552 76624 87616
rect 76688 87552 76694 87616
rect 76378 87551 76694 87552
rect 5950 87072 6266 87073
rect 5950 87008 5956 87072
rect 6020 87008 6036 87072
rect 6100 87008 6116 87072
rect 6180 87008 6196 87072
rect 6260 87008 6266 87072
rect 5950 87007 6266 87008
rect 18718 87072 19034 87073
rect 18718 87008 18724 87072
rect 18788 87008 18804 87072
rect 18868 87008 18884 87072
rect 18948 87008 18964 87072
rect 19028 87008 19034 87072
rect 18718 87007 19034 87008
rect 37718 87072 38034 87073
rect 37718 87008 37724 87072
rect 37788 87008 37804 87072
rect 37868 87008 37884 87072
rect 37948 87008 37964 87072
rect 38028 87008 38034 87072
rect 37718 87007 38034 87008
rect 56718 87072 57034 87073
rect 56718 87008 56724 87072
rect 56788 87008 56804 87072
rect 56868 87008 56884 87072
rect 56948 87008 56964 87072
rect 57028 87008 57034 87072
rect 56718 87007 57034 87008
rect 75718 87072 76034 87073
rect 75718 87008 75724 87072
rect 75788 87008 75804 87072
rect 75868 87008 75884 87072
rect 75948 87008 75964 87072
rect 76028 87008 76034 87072
rect 75718 87007 76034 87008
rect 87094 87072 87410 87073
rect 87094 87008 87100 87072
rect 87164 87008 87180 87072
rect 87244 87008 87260 87072
rect 87324 87008 87340 87072
rect 87404 87008 87410 87072
rect 87094 87007 87410 87008
rect 6686 86528 7002 86529
rect 6686 86464 6692 86528
rect 6756 86464 6772 86528
rect 6836 86464 6852 86528
rect 6916 86464 6932 86528
rect 6996 86464 7002 86528
rect 6686 86463 7002 86464
rect 19378 86528 19694 86529
rect 19378 86464 19384 86528
rect 19448 86464 19464 86528
rect 19528 86464 19544 86528
rect 19608 86464 19624 86528
rect 19688 86464 19694 86528
rect 19378 86463 19694 86464
rect 38378 86528 38694 86529
rect 38378 86464 38384 86528
rect 38448 86464 38464 86528
rect 38528 86464 38544 86528
rect 38608 86464 38624 86528
rect 38688 86464 38694 86528
rect 38378 86463 38694 86464
rect 57378 86528 57694 86529
rect 57378 86464 57384 86528
rect 57448 86464 57464 86528
rect 57528 86464 57544 86528
rect 57608 86464 57624 86528
rect 57688 86464 57694 86528
rect 57378 86463 57694 86464
rect 76378 86528 76694 86529
rect 76378 86464 76384 86528
rect 76448 86464 76464 86528
rect 76528 86464 76544 86528
rect 76608 86464 76624 86528
rect 76688 86464 76694 86528
rect 76378 86463 76694 86464
rect 87830 86528 88146 86529
rect 87830 86464 87836 86528
rect 87900 86464 87916 86528
rect 87980 86464 87996 86528
rect 88060 86464 88076 86528
rect 88140 86464 88146 86528
rect 87830 86463 88146 86464
rect 5950 85984 6266 85985
rect 5950 85920 5956 85984
rect 6020 85920 6036 85984
rect 6100 85920 6116 85984
rect 6180 85920 6196 85984
rect 6260 85920 6266 85984
rect 5950 85919 6266 85920
rect 87094 85984 87410 85985
rect 87094 85920 87100 85984
rect 87164 85920 87180 85984
rect 87244 85920 87260 85984
rect 87324 85920 87340 85984
rect 87404 85920 87410 85984
rect 87094 85919 87410 85920
rect 6686 85440 7002 85441
rect 6686 85376 6692 85440
rect 6756 85376 6772 85440
rect 6836 85376 6852 85440
rect 6916 85376 6932 85440
rect 6996 85376 7002 85440
rect 6686 85375 7002 85376
rect 87830 85440 88146 85441
rect 87830 85376 87836 85440
rect 87900 85376 87916 85440
rect 87980 85376 87996 85440
rect 88060 85376 88076 85440
rect 88140 85376 88146 85440
rect 87830 85375 88146 85376
rect 5950 84896 6266 84897
rect 5950 84832 5956 84896
rect 6020 84832 6036 84896
rect 6100 84832 6116 84896
rect 6180 84832 6196 84896
rect 6260 84832 6266 84896
rect 5950 84831 6266 84832
rect 87094 84896 87410 84897
rect 87094 84832 87100 84896
rect 87164 84832 87180 84896
rect 87244 84832 87260 84896
rect 87324 84832 87340 84896
rect 87404 84832 87410 84896
rect 87094 84831 87410 84832
rect 8421 84386 8487 84389
rect 14401 84386 14467 84389
rect 8421 84384 14467 84386
rect 6686 84352 7002 84353
rect 6686 84288 6692 84352
rect 6756 84288 6772 84352
rect 6836 84288 6852 84352
rect 6916 84288 6932 84352
rect 6996 84288 7002 84352
rect 8421 84328 8426 84384
rect 8482 84328 14406 84384
rect 14462 84328 14467 84384
rect 8421 84326 14467 84328
rect 8421 84323 8487 84326
rect 14401 84323 14467 84326
rect 87830 84352 88146 84353
rect 6686 84287 7002 84288
rect 87830 84288 87836 84352
rect 87900 84288 87916 84352
rect 87980 84288 87996 84352
rect 88060 84288 88076 84352
rect 88140 84288 88146 84352
rect 87830 84287 88146 84288
rect 9801 84250 9867 84253
rect 51431 84250 51497 84253
rect 9801 84248 51497 84250
rect 9801 84192 9806 84248
rect 9862 84192 51436 84248
rect 51492 84192 51497 84248
rect 9801 84190 51497 84192
rect 9801 84187 9867 84190
rect 51431 84187 51497 84190
rect 5950 83808 6266 83809
rect 5950 83744 5956 83808
rect 6020 83744 6036 83808
rect 6100 83744 6116 83808
rect 6180 83744 6196 83808
rect 6260 83744 6266 83808
rect 5950 83743 6266 83744
rect 87094 83808 87410 83809
rect 87094 83744 87100 83808
rect 87164 83744 87180 83808
rect 87244 83744 87260 83808
rect 87324 83744 87340 83808
rect 87404 83744 87410 83808
rect 87094 83743 87410 83744
rect 6686 83264 7002 83265
rect 6686 83200 6692 83264
rect 6756 83200 6772 83264
rect 6836 83200 6852 83264
rect 6916 83200 6932 83264
rect 6996 83200 7002 83264
rect 6686 83199 7002 83200
rect 87830 83264 88146 83265
rect 87830 83200 87836 83264
rect 87900 83200 87916 83264
rect 87980 83200 87996 83264
rect 88060 83200 88076 83264
rect 88140 83200 88146 83264
rect 87830 83199 88146 83200
rect 5950 82720 6266 82721
rect 5950 82656 5956 82720
rect 6020 82656 6036 82720
rect 6100 82656 6116 82720
rect 6180 82656 6196 82720
rect 6260 82656 6266 82720
rect 5950 82655 6266 82656
rect 87094 82720 87410 82721
rect 87094 82656 87100 82720
rect 87164 82656 87180 82720
rect 87244 82656 87260 82720
rect 87324 82656 87340 82720
rect 87404 82656 87410 82720
rect 87094 82655 87410 82656
rect 6686 82176 7002 82177
rect 6686 82112 6692 82176
rect 6756 82112 6772 82176
rect 6836 82112 6852 82176
rect 6916 82112 6932 82176
rect 6996 82112 7002 82176
rect 6686 82111 7002 82112
rect 87830 82176 88146 82177
rect 87830 82112 87836 82176
rect 87900 82112 87916 82176
rect 87980 82112 87996 82176
rect 88060 82112 88076 82176
rect 88140 82112 88146 82176
rect 87830 82111 88146 82112
rect 5950 81632 6266 81633
rect 5950 81568 5956 81632
rect 6020 81568 6036 81632
rect 6100 81568 6116 81632
rect 6180 81568 6196 81632
rect 6260 81568 6266 81632
rect 5950 81567 6266 81568
rect 87094 81632 87410 81633
rect 87094 81568 87100 81632
rect 87164 81568 87180 81632
rect 87244 81568 87260 81632
rect 87324 81568 87340 81632
rect 87404 81568 87410 81632
rect 87094 81567 87410 81568
rect 6686 81088 7002 81089
rect 6686 81024 6692 81088
rect 6756 81024 6772 81088
rect 6836 81024 6852 81088
rect 6916 81024 6932 81088
rect 6996 81024 7002 81088
rect 6686 81023 7002 81024
rect 87830 81088 88146 81089
rect 87830 81024 87836 81088
rect 87900 81024 87916 81088
rect 87980 81024 87996 81088
rect 88060 81024 88076 81088
rect 88140 81024 88146 81088
rect 87830 81023 88146 81024
rect 1600 80578 2400 80608
rect 2901 80578 2967 80581
rect 1600 80576 2967 80578
rect 1600 80520 2906 80576
rect 2962 80520 2967 80576
rect 88645 80578 88711 80581
rect 91400 80578 92200 80608
rect 88645 80576 92200 80578
rect 1600 80518 2967 80520
rect 1600 80488 2400 80518
rect 2901 80515 2967 80518
rect 5950 80544 6266 80545
rect 5950 80480 5956 80544
rect 6020 80480 6036 80544
rect 6100 80480 6116 80544
rect 6180 80480 6196 80544
rect 6260 80480 6266 80544
rect 5950 80479 6266 80480
rect 87094 80544 87410 80545
rect 87094 80480 87100 80544
rect 87164 80480 87180 80544
rect 87244 80480 87260 80544
rect 87324 80480 87340 80544
rect 87404 80480 87410 80544
rect 88645 80520 88650 80576
rect 88706 80520 92200 80576
rect 88645 80518 92200 80520
rect 88645 80515 88711 80518
rect 91400 80488 92200 80518
rect 87094 80479 87410 80480
rect 7133 80442 7199 80445
rect 84321 80442 84387 80445
rect 7133 80440 9634 80442
rect 7133 80384 7138 80440
rect 7194 80410 9634 80440
rect 83940 80440 84387 80442
rect 7194 80384 10156 80410
rect 7133 80382 10156 80384
rect 83940 80384 84326 80440
rect 84382 80384 84387 80440
rect 83940 80382 84387 80384
rect 7133 80379 7199 80382
rect 9574 80350 10156 80382
rect 84321 80379 84387 80382
rect 6686 80000 7002 80001
rect 6686 79936 6692 80000
rect 6756 79936 6772 80000
rect 6836 79936 6852 80000
rect 6916 79936 6932 80000
rect 6996 79936 7002 80000
rect 6686 79935 7002 79936
rect 87830 80000 88146 80001
rect 87830 79936 87836 80000
rect 87900 79936 87916 80000
rect 87980 79936 87996 80000
rect 88060 79936 88076 80000
rect 88140 79936 88146 80000
rect 87830 79935 88146 79936
rect 5950 79456 6266 79457
rect 5950 79392 5956 79456
rect 6020 79392 6036 79456
rect 6100 79392 6116 79456
rect 6180 79392 6196 79456
rect 6260 79392 6266 79456
rect 5950 79391 6266 79392
rect 87094 79456 87410 79457
rect 87094 79392 87100 79456
rect 87164 79392 87180 79456
rect 87244 79392 87260 79456
rect 87324 79392 87340 79456
rect 87404 79392 87410 79456
rect 87094 79391 87410 79392
rect 7133 79354 7199 79357
rect 84321 79354 84387 79357
rect 7133 79352 9634 79354
rect 7133 79296 7138 79352
rect 7194 79322 9634 79352
rect 83940 79352 84387 79354
rect 7194 79296 10156 79322
rect 7133 79294 10156 79296
rect 83940 79296 84326 79352
rect 84382 79296 84387 79352
rect 83940 79294 84387 79296
rect 7133 79291 7199 79294
rect 9574 79262 10156 79294
rect 84321 79291 84387 79294
rect 1600 79218 2400 79248
rect 2717 79218 2783 79221
rect 1600 79216 2783 79218
rect 1600 79160 2722 79216
rect 2778 79160 2783 79216
rect 1600 79158 2783 79160
rect 1600 79128 2400 79158
rect 2717 79155 2783 79158
rect 88645 79218 88711 79221
rect 91400 79218 92200 79248
rect 88645 79216 92200 79218
rect 88645 79160 88650 79216
rect 88706 79160 92200 79216
rect 88645 79158 92200 79160
rect 88645 79155 88711 79158
rect 91400 79128 92200 79158
rect 6686 78912 7002 78913
rect 6686 78848 6692 78912
rect 6756 78848 6772 78912
rect 6836 78848 6852 78912
rect 6916 78848 6932 78912
rect 6996 78848 7002 78912
rect 6686 78847 7002 78848
rect 87830 78912 88146 78913
rect 87830 78848 87836 78912
rect 87900 78848 87916 78912
rect 87980 78848 87996 78912
rect 88060 78848 88076 78912
rect 88140 78848 88146 78912
rect 87830 78847 88146 78848
rect 1600 78538 2400 78568
rect 2901 78538 2967 78541
rect 1600 78536 2967 78538
rect 1600 78480 2906 78536
rect 2962 78480 2967 78536
rect 1600 78478 2967 78480
rect 1600 78448 2400 78478
rect 2901 78475 2967 78478
rect 88645 78538 88711 78541
rect 91400 78538 92200 78568
rect 88645 78536 92200 78538
rect 88645 78480 88650 78536
rect 88706 78480 92200 78536
rect 88645 78478 92200 78480
rect 88645 78475 88711 78478
rect 91400 78448 92200 78478
rect 5950 78368 6266 78369
rect 5950 78304 5956 78368
rect 6020 78304 6036 78368
rect 6100 78304 6116 78368
rect 6180 78304 6196 78368
rect 6260 78304 6266 78368
rect 5950 78303 6266 78304
rect 87094 78368 87410 78369
rect 87094 78304 87100 78368
rect 87164 78304 87180 78368
rect 87244 78304 87260 78368
rect 87324 78304 87340 78368
rect 87404 78304 87410 78368
rect 87094 78303 87410 78304
rect 7133 78266 7199 78269
rect 84321 78266 84387 78269
rect 7133 78264 9634 78266
rect 7133 78208 7138 78264
rect 7194 78234 9634 78264
rect 83940 78264 84387 78266
rect 7194 78208 10156 78234
rect 7133 78206 10156 78208
rect 83940 78208 84326 78264
rect 84382 78208 84387 78264
rect 83940 78206 84387 78208
rect 7133 78203 7199 78206
rect 9574 78174 10156 78206
rect 84321 78203 84387 78206
rect 6686 77824 7002 77825
rect 6686 77760 6692 77824
rect 6756 77760 6772 77824
rect 6836 77760 6852 77824
rect 6916 77760 6932 77824
rect 6996 77760 7002 77824
rect 6686 77759 7002 77760
rect 87830 77824 88146 77825
rect 87830 77760 87836 77824
rect 87900 77760 87916 77824
rect 87980 77760 87996 77824
rect 88060 77760 88076 77824
rect 88140 77760 88146 77824
rect 87830 77759 88146 77760
rect 5950 77280 6266 77281
rect 5950 77216 5956 77280
rect 6020 77216 6036 77280
rect 6100 77216 6116 77280
rect 6180 77216 6196 77280
rect 6260 77216 6266 77280
rect 5950 77215 6266 77216
rect 87094 77280 87410 77281
rect 87094 77216 87100 77280
rect 87164 77216 87180 77280
rect 87244 77216 87260 77280
rect 87324 77216 87340 77280
rect 87404 77216 87410 77280
rect 87094 77215 87410 77216
rect 1600 77178 2400 77208
rect 4373 77178 4439 77181
rect 84321 77178 84387 77181
rect 1600 77176 4439 77178
rect 1600 77120 4378 77176
rect 4434 77120 4439 77176
rect 83940 77176 84387 77178
rect 1600 77118 4439 77120
rect 1600 77088 2400 77118
rect 4373 77115 4439 77118
rect 9574 77086 10156 77146
rect 83940 77120 84326 77176
rect 84382 77120 84387 77176
rect 83940 77118 84387 77120
rect 84321 77115 84387 77118
rect 90025 77178 90091 77181
rect 91400 77178 92200 77208
rect 90025 77176 92200 77178
rect 90025 77120 90030 77176
rect 90086 77120 92200 77176
rect 90025 77118 92200 77120
rect 90025 77115 90091 77118
rect 91400 77088 92200 77118
rect 5661 77042 5727 77045
rect 9574 77042 9634 77086
rect 5661 77040 9634 77042
rect 5661 76984 5666 77040
rect 5722 76984 9634 77040
rect 5661 76982 9634 76984
rect 5661 76979 5727 76982
rect 6686 76736 7002 76737
rect 6686 76672 6692 76736
rect 6756 76672 6772 76736
rect 6836 76672 6852 76736
rect 6916 76672 6932 76736
rect 6996 76672 7002 76736
rect 6686 76671 7002 76672
rect 87830 76736 88146 76737
rect 87830 76672 87836 76736
rect 87900 76672 87916 76736
rect 87980 76672 87996 76736
rect 88060 76672 88076 76736
rect 88140 76672 88146 76736
rect 87830 76671 88146 76672
rect 5950 76192 6266 76193
rect 5950 76128 5956 76192
rect 6020 76128 6036 76192
rect 6100 76128 6116 76192
rect 6180 76128 6196 76192
rect 6260 76128 6266 76192
rect 5950 76127 6266 76128
rect 87094 76192 87410 76193
rect 87094 76128 87100 76192
rect 87164 76128 87180 76192
rect 87244 76128 87260 76192
rect 87324 76128 87340 76192
rect 87404 76128 87410 76192
rect 87094 76127 87410 76128
rect 7133 76090 7199 76093
rect 7133 76088 9634 76090
rect 7133 76032 7138 76088
rect 7194 76058 9634 76088
rect 7194 76032 10156 76058
rect 7133 76030 10156 76032
rect 7133 76027 7199 76030
rect 9574 75998 10156 76030
rect 84321 76022 84387 76025
rect 83940 76020 84387 76022
rect 83940 75964 84326 76020
rect 84382 75964 84387 76020
rect 83940 75962 84387 75964
rect 84321 75959 84387 75962
rect 1600 75818 2400 75848
rect 2901 75818 2967 75821
rect 1600 75816 2967 75818
rect 1600 75760 2906 75816
rect 2962 75760 2967 75816
rect 1600 75758 2967 75760
rect 1600 75728 2400 75758
rect 2901 75755 2967 75758
rect 88737 75818 88803 75821
rect 91400 75818 92200 75848
rect 88737 75816 92200 75818
rect 88737 75760 88742 75816
rect 88798 75760 92200 75816
rect 88737 75758 92200 75760
rect 88737 75755 88803 75758
rect 91400 75728 92200 75758
rect 6686 75648 7002 75649
rect 6686 75584 6692 75648
rect 6756 75584 6772 75648
rect 6836 75584 6852 75648
rect 6916 75584 6932 75648
rect 6996 75584 7002 75648
rect 6686 75583 7002 75584
rect 87830 75648 88146 75649
rect 87830 75584 87836 75648
rect 87900 75584 87916 75648
rect 87980 75584 87996 75648
rect 88060 75584 88076 75648
rect 88140 75584 88146 75648
rect 87830 75583 88146 75584
rect 1600 75138 2400 75168
rect 2901 75138 2967 75141
rect 1600 75136 2967 75138
rect 1600 75080 2906 75136
rect 2962 75080 2967 75136
rect 88553 75138 88619 75141
rect 91400 75138 92200 75168
rect 88553 75136 92200 75138
rect 1600 75078 2967 75080
rect 1600 75048 2400 75078
rect 2901 75075 2967 75078
rect 5950 75104 6266 75105
rect 5950 75040 5956 75104
rect 6020 75040 6036 75104
rect 6100 75040 6116 75104
rect 6180 75040 6196 75104
rect 6260 75040 6266 75104
rect 5950 75039 6266 75040
rect 87094 75104 87410 75105
rect 87094 75040 87100 75104
rect 87164 75040 87180 75104
rect 87244 75040 87260 75104
rect 87324 75040 87340 75104
rect 87404 75040 87410 75104
rect 88553 75080 88558 75136
rect 88614 75080 92200 75136
rect 88553 75078 92200 75080
rect 88553 75075 88619 75078
rect 91400 75048 92200 75078
rect 87094 75039 87410 75040
rect 7133 75002 7199 75005
rect 84321 75002 84387 75005
rect 7133 75000 9634 75002
rect 7133 74944 7138 75000
rect 7194 74970 9634 75000
rect 83940 75000 84387 75002
rect 7194 74944 10156 74970
rect 7133 74942 10156 74944
rect 83940 74944 84326 75000
rect 84382 74944 84387 75000
rect 83940 74942 84387 74944
rect 7133 74939 7199 74942
rect 9574 74910 10156 74942
rect 84321 74939 84387 74942
rect 6686 74560 7002 74561
rect 6686 74496 6692 74560
rect 6756 74496 6772 74560
rect 6836 74496 6852 74560
rect 6916 74496 6932 74560
rect 6996 74496 7002 74560
rect 6686 74495 7002 74496
rect 87830 74560 88146 74561
rect 87830 74496 87836 74560
rect 87900 74496 87916 74560
rect 87980 74496 87996 74560
rect 88060 74496 88076 74560
rect 88140 74496 88146 74560
rect 87830 74495 88146 74496
rect 5950 74016 6266 74017
rect 5950 73952 5956 74016
rect 6020 73952 6036 74016
rect 6100 73952 6116 74016
rect 6180 73952 6196 74016
rect 6260 73952 6266 74016
rect 5950 73951 6266 73952
rect 87094 74016 87410 74017
rect 87094 73952 87100 74016
rect 87164 73952 87180 74016
rect 87244 73952 87260 74016
rect 87324 73952 87340 74016
rect 87404 73952 87410 74016
rect 87094 73951 87410 73952
rect 7133 73914 7199 73917
rect 84321 73914 84387 73917
rect 7133 73912 9634 73914
rect 7133 73856 7138 73912
rect 7194 73882 9634 73912
rect 83940 73912 84387 73914
rect 7194 73856 10156 73882
rect 7133 73854 10156 73856
rect 83940 73856 84326 73912
rect 84382 73856 84387 73912
rect 83940 73854 84387 73856
rect 7133 73851 7199 73854
rect 9574 73822 10156 73854
rect 84321 73851 84387 73854
rect 1600 73778 2400 73808
rect 2901 73778 2967 73781
rect 1600 73776 2967 73778
rect 1600 73720 2906 73776
rect 2962 73720 2967 73776
rect 1600 73718 2967 73720
rect 1600 73688 2400 73718
rect 2901 73715 2967 73718
rect 88553 73778 88619 73781
rect 91400 73778 92200 73808
rect 88553 73776 92200 73778
rect 88553 73720 88558 73776
rect 88614 73720 92200 73776
rect 88553 73718 92200 73720
rect 88553 73715 88619 73718
rect 91400 73688 92200 73718
rect 6686 73472 7002 73473
rect 6686 73408 6692 73472
rect 6756 73408 6772 73472
rect 6836 73408 6852 73472
rect 6916 73408 6932 73472
rect 6996 73408 7002 73472
rect 6686 73407 7002 73408
rect 87830 73472 88146 73473
rect 87830 73408 87836 73472
rect 87900 73408 87916 73472
rect 87980 73408 87996 73472
rect 88060 73408 88076 73472
rect 88140 73408 88146 73472
rect 87830 73407 88146 73408
rect 1600 73098 2400 73128
rect 2901 73098 2967 73101
rect 1600 73096 2967 73098
rect 1600 73040 2906 73096
rect 2962 73040 2967 73096
rect 1600 73038 2967 73040
rect 1600 73008 2400 73038
rect 2901 73035 2967 73038
rect 88645 73098 88711 73101
rect 91400 73098 92200 73128
rect 88645 73096 92200 73098
rect 88645 73040 88650 73096
rect 88706 73040 92200 73096
rect 88645 73038 92200 73040
rect 88645 73035 88711 73038
rect 91400 73008 92200 73038
rect 5950 72928 6266 72929
rect 5950 72864 5956 72928
rect 6020 72864 6036 72928
rect 6100 72864 6116 72928
rect 6180 72864 6196 72928
rect 6260 72864 6266 72928
rect 5950 72863 6266 72864
rect 87094 72928 87410 72929
rect 87094 72864 87100 72928
rect 87164 72864 87180 72928
rect 87244 72864 87260 72928
rect 87324 72864 87340 72928
rect 87404 72864 87410 72928
rect 87094 72863 87410 72864
rect 7133 72826 7199 72829
rect 84321 72826 84387 72829
rect 7133 72824 9634 72826
rect 7133 72768 7138 72824
rect 7194 72794 9634 72824
rect 83940 72824 84387 72826
rect 7194 72768 10156 72794
rect 7133 72766 10156 72768
rect 83940 72768 84326 72824
rect 84382 72768 84387 72824
rect 83940 72766 84387 72768
rect 7133 72763 7199 72766
rect 9574 72734 10156 72766
rect 84321 72763 84387 72766
rect 6686 72384 7002 72385
rect 6686 72320 6692 72384
rect 6756 72320 6772 72384
rect 6836 72320 6852 72384
rect 6916 72320 6932 72384
rect 6996 72320 7002 72384
rect 6686 72319 7002 72320
rect 87830 72384 88146 72385
rect 87830 72320 87836 72384
rect 87900 72320 87916 72384
rect 87980 72320 87996 72384
rect 88060 72320 88076 72384
rect 88140 72320 88146 72384
rect 87830 72319 88146 72320
rect 87173 72010 87239 72013
rect 83910 72008 87239 72010
rect 83910 71952 87178 72008
rect 87234 71952 87239 72008
rect 83910 71950 87239 71952
rect 5950 71840 6266 71841
rect 5950 71776 5956 71840
rect 6020 71776 6036 71840
rect 6100 71776 6116 71840
rect 6180 71776 6196 71840
rect 6260 71776 6266 71840
rect 5950 71775 6266 71776
rect 1600 71738 2400 71768
rect 4373 71738 4439 71741
rect 1600 71736 4439 71738
rect 1600 71680 4378 71736
rect 4434 71680 4439 71736
rect 83910 71708 83970 71950
rect 87173 71947 87239 71950
rect 87094 71840 87410 71841
rect 87094 71776 87100 71840
rect 87164 71776 87180 71840
rect 87244 71776 87260 71840
rect 87324 71776 87340 71840
rect 87404 71776 87410 71840
rect 87094 71775 87410 71776
rect 90117 71738 90183 71741
rect 91400 71738 92200 71768
rect 90117 71736 92200 71738
rect 1600 71678 4439 71680
rect 1600 71648 2400 71678
rect 4373 71675 4439 71678
rect 9574 71646 10156 71706
rect 90117 71680 90122 71736
rect 90178 71680 92200 71736
rect 90117 71678 92200 71680
rect 90117 71675 90183 71678
rect 91400 71648 92200 71678
rect 5661 71602 5727 71605
rect 9574 71602 9634 71646
rect 5661 71600 9634 71602
rect 5661 71544 5666 71600
rect 5722 71544 9634 71600
rect 5661 71542 9634 71544
rect 5661 71539 5727 71542
rect 6686 71296 7002 71297
rect 6686 71232 6692 71296
rect 6756 71232 6772 71296
rect 6836 71232 6852 71296
rect 6916 71232 6932 71296
rect 6996 71232 7002 71296
rect 6686 71231 7002 71232
rect 87830 71296 88146 71297
rect 87830 71232 87836 71296
rect 87900 71232 87916 71296
rect 87980 71232 87996 71296
rect 88060 71232 88076 71296
rect 88140 71232 88146 71296
rect 87830 71231 88146 71232
rect 5661 70922 5727 70925
rect 5661 70920 9818 70922
rect 5661 70864 5666 70920
rect 5722 70864 9818 70920
rect 5661 70862 9818 70864
rect 5661 70859 5727 70862
rect 5950 70752 6266 70753
rect 5950 70688 5956 70752
rect 6020 70688 6036 70752
rect 6100 70688 6116 70752
rect 6180 70688 6196 70752
rect 6260 70688 6266 70752
rect 5950 70687 6266 70688
rect 9758 70618 9818 70862
rect 87094 70752 87410 70753
rect 87094 70688 87100 70752
rect 87164 70688 87180 70752
rect 87244 70688 87260 70752
rect 87324 70688 87340 70752
rect 87404 70688 87410 70752
rect 87094 70687 87410 70688
rect 84321 70650 84387 70653
rect 83940 70648 84387 70650
rect 9758 70558 10156 70618
rect 83940 70592 84326 70648
rect 84382 70592 84387 70648
rect 83940 70590 84387 70592
rect 84321 70587 84387 70590
rect 1600 70378 2400 70408
rect 2901 70378 2967 70381
rect 1600 70376 2967 70378
rect 1600 70320 2906 70376
rect 2962 70320 2967 70376
rect 1600 70318 2967 70320
rect 1600 70288 2400 70318
rect 2901 70315 2967 70318
rect 89933 70378 89999 70381
rect 91400 70378 92200 70408
rect 89933 70376 92200 70378
rect 89933 70320 89938 70376
rect 89994 70320 92200 70376
rect 89933 70318 92200 70320
rect 89933 70315 89999 70318
rect 91400 70288 92200 70318
rect 6686 70208 7002 70209
rect 6686 70144 6692 70208
rect 6756 70144 6772 70208
rect 6836 70144 6852 70208
rect 6916 70144 6932 70208
rect 6996 70144 7002 70208
rect 6686 70143 7002 70144
rect 87830 70208 88146 70209
rect 87830 70144 87836 70208
rect 87900 70144 87916 70208
rect 87980 70144 87996 70208
rect 88060 70144 88076 70208
rect 88140 70144 88146 70208
rect 87830 70143 88146 70144
rect 1600 69698 2400 69728
rect 2901 69698 2967 69701
rect 1600 69696 2967 69698
rect 1600 69640 2906 69696
rect 2962 69640 2967 69696
rect 88553 69698 88619 69701
rect 91400 69698 92200 69728
rect 88553 69696 92200 69698
rect 1600 69638 2967 69640
rect 1600 69608 2400 69638
rect 2901 69635 2967 69638
rect 5950 69664 6266 69665
rect 5950 69600 5956 69664
rect 6020 69600 6036 69664
rect 6100 69600 6116 69664
rect 6180 69600 6196 69664
rect 6260 69600 6266 69664
rect 5950 69599 6266 69600
rect 87094 69664 87410 69665
rect 87094 69600 87100 69664
rect 87164 69600 87180 69664
rect 87244 69600 87260 69664
rect 87324 69600 87340 69664
rect 87404 69600 87410 69664
rect 88553 69640 88558 69696
rect 88614 69640 92200 69696
rect 88553 69638 92200 69640
rect 88553 69635 88619 69638
rect 91400 69608 92200 69638
rect 87094 69599 87410 69600
rect 7133 69562 7199 69565
rect 84321 69562 84387 69565
rect 7133 69560 9634 69562
rect 7133 69504 7138 69560
rect 7194 69530 9634 69560
rect 83940 69560 84387 69562
rect 7194 69504 10156 69530
rect 7133 69502 10156 69504
rect 83940 69504 84326 69560
rect 84382 69504 84387 69560
rect 83940 69502 84387 69504
rect 7133 69499 7199 69502
rect 9574 69470 10156 69502
rect 84321 69499 84387 69502
rect 6686 69120 7002 69121
rect 6686 69056 6692 69120
rect 6756 69056 6772 69120
rect 6836 69056 6852 69120
rect 6916 69056 6932 69120
rect 6996 69056 7002 69120
rect 6686 69055 7002 69056
rect 87830 69120 88146 69121
rect 87830 69056 87836 69120
rect 87900 69056 87916 69120
rect 87980 69056 87996 69120
rect 88060 69056 88076 69120
rect 88140 69056 88146 69120
rect 87830 69055 88146 69056
rect 89933 69018 89999 69021
rect 91400 69018 92200 69048
rect 89933 69016 92200 69018
rect 89933 68960 89938 69016
rect 89994 68960 92200 69016
rect 89933 68958 92200 68960
rect 89933 68955 89999 68958
rect 91400 68928 92200 68958
rect 5950 68576 6266 68577
rect 5950 68512 5956 68576
rect 6020 68512 6036 68576
rect 6100 68512 6116 68576
rect 6180 68512 6196 68576
rect 6260 68512 6266 68576
rect 5950 68511 6266 68512
rect 87094 68576 87410 68577
rect 87094 68512 87100 68576
rect 87164 68512 87180 68576
rect 87244 68512 87260 68576
rect 87324 68512 87340 68576
rect 87404 68512 87410 68576
rect 87094 68511 87410 68512
rect 7133 68474 7199 68477
rect 84321 68474 84387 68477
rect 7133 68472 9634 68474
rect 7133 68416 7138 68472
rect 7194 68442 9634 68472
rect 83940 68472 84387 68474
rect 7194 68416 10156 68442
rect 7133 68414 10156 68416
rect 83940 68416 84326 68472
rect 84382 68416 84387 68472
rect 83940 68414 84387 68416
rect 7133 68411 7199 68414
rect 9574 68382 10156 68414
rect 84321 68411 84387 68414
rect 1600 68338 2400 68368
rect 2901 68338 2967 68341
rect 1600 68336 2967 68338
rect 1600 68280 2906 68336
rect 2962 68280 2967 68336
rect 1600 68278 2967 68280
rect 1600 68248 2400 68278
rect 2901 68275 2967 68278
rect 88645 68338 88711 68341
rect 91400 68338 92200 68368
rect 88645 68336 92200 68338
rect 88645 68280 88650 68336
rect 88706 68280 92200 68336
rect 88645 68278 92200 68280
rect 88645 68275 88711 68278
rect 91400 68248 92200 68278
rect 6686 68032 7002 68033
rect 6686 67968 6692 68032
rect 6756 67968 6772 68032
rect 6836 67968 6852 68032
rect 6916 67968 6932 68032
rect 6996 67968 7002 68032
rect 6686 67967 7002 67968
rect 87830 68032 88146 68033
rect 87830 67968 87836 68032
rect 87900 67968 87916 68032
rect 87980 67968 87996 68032
rect 88060 67968 88076 68032
rect 88140 67968 88146 68032
rect 87830 67967 88146 67968
rect 1600 67658 2400 67688
rect 2901 67658 2967 67661
rect 1600 67656 2967 67658
rect 1600 67600 2906 67656
rect 2962 67600 2967 67656
rect 1600 67598 2967 67600
rect 1600 67568 2400 67598
rect 2901 67595 2967 67598
rect 88645 67658 88711 67661
rect 91400 67658 92200 67688
rect 88645 67656 92200 67658
rect 88645 67600 88650 67656
rect 88706 67600 92200 67656
rect 88645 67598 92200 67600
rect 88645 67595 88711 67598
rect 91400 67568 92200 67598
rect 5950 67488 6266 67489
rect 5950 67424 5956 67488
rect 6020 67424 6036 67488
rect 6100 67424 6116 67488
rect 6180 67424 6196 67488
rect 6260 67424 6266 67488
rect 5950 67423 6266 67424
rect 87094 67488 87410 67489
rect 87094 67424 87100 67488
rect 87164 67424 87180 67488
rect 87244 67424 87260 67488
rect 87324 67424 87340 67488
rect 87404 67424 87410 67488
rect 87094 67423 87410 67424
rect 7133 67386 7199 67389
rect 84321 67386 84387 67389
rect 7133 67384 9634 67386
rect 7133 67328 7138 67384
rect 7194 67354 9634 67384
rect 83940 67384 84387 67386
rect 7194 67328 10156 67354
rect 7133 67326 10156 67328
rect 83940 67328 84326 67384
rect 84382 67328 84387 67384
rect 83940 67326 84387 67328
rect 7133 67323 7199 67326
rect 9574 67294 10156 67326
rect 84321 67323 84387 67326
rect 6686 66944 7002 66945
rect 6686 66880 6692 66944
rect 6756 66880 6772 66944
rect 6836 66880 6852 66944
rect 6916 66880 6932 66944
rect 6996 66880 7002 66944
rect 6686 66879 7002 66880
rect 87830 66944 88146 66945
rect 87830 66880 87836 66944
rect 87900 66880 87916 66944
rect 87980 66880 87996 66944
rect 88060 66880 88076 66944
rect 88140 66880 88146 66944
rect 87830 66879 88146 66880
rect 5950 66400 6266 66401
rect 5950 66336 5956 66400
rect 6020 66336 6036 66400
rect 6100 66336 6116 66400
rect 6180 66336 6196 66400
rect 6260 66336 6266 66400
rect 5950 66335 6266 66336
rect 87094 66400 87410 66401
rect 87094 66336 87100 66400
rect 87164 66336 87180 66400
rect 87244 66336 87260 66400
rect 87324 66336 87340 66400
rect 87404 66336 87410 66400
rect 87094 66335 87410 66336
rect 1600 66298 2400 66328
rect 4373 66298 4439 66301
rect 90117 66298 90183 66301
rect 91400 66298 92200 66328
rect 1600 66296 4439 66298
rect 1600 66240 4378 66296
rect 4434 66240 4439 66296
rect 1600 66238 4439 66240
rect 1600 66208 2400 66238
rect 4373 66235 4439 66238
rect 9574 66206 10156 66266
rect 83940 66238 85810 66298
rect 5477 66162 5543 66165
rect 9574 66162 9634 66206
rect 5477 66160 9634 66162
rect 5477 66104 5482 66160
rect 5538 66104 9634 66160
rect 5477 66102 9634 66104
rect 85750 66162 85810 66238
rect 90117 66296 92200 66298
rect 90117 66240 90122 66296
rect 90178 66240 92200 66296
rect 90117 66238 92200 66240
rect 90117 66235 90183 66238
rect 91400 66208 92200 66238
rect 87449 66162 87515 66165
rect 85750 66160 87515 66162
rect 85750 66104 87454 66160
rect 87510 66104 87515 66160
rect 85750 66102 87515 66104
rect 5477 66099 5543 66102
rect 87449 66099 87515 66102
rect 6686 65856 7002 65857
rect 6686 65792 6692 65856
rect 6756 65792 6772 65856
rect 6836 65792 6852 65856
rect 6916 65792 6932 65856
rect 6996 65792 7002 65856
rect 6686 65791 7002 65792
rect 87830 65856 88146 65857
rect 87830 65792 87836 65856
rect 87900 65792 87916 65856
rect 87980 65792 87996 65856
rect 88060 65792 88076 65856
rect 88140 65792 88146 65856
rect 87830 65791 88146 65792
rect 5385 65482 5451 65485
rect 5385 65480 9634 65482
rect 5385 65424 5390 65480
rect 5446 65424 9634 65480
rect 5385 65422 9634 65424
rect 5385 65419 5451 65422
rect 5950 65312 6266 65313
rect 5950 65248 5956 65312
rect 6020 65248 6036 65312
rect 6100 65248 6116 65312
rect 6180 65248 6196 65312
rect 6260 65248 6266 65312
rect 5950 65247 6266 65248
rect 9574 65178 9634 65422
rect 87094 65312 87410 65313
rect 87094 65248 87100 65312
rect 87164 65248 87180 65312
rect 87244 65248 87260 65312
rect 87324 65248 87340 65312
rect 87404 65248 87410 65312
rect 87094 65247 87410 65248
rect 9574 65118 10156 65178
rect 84321 65142 84387 65145
rect 83940 65140 84387 65142
rect 83940 65084 84326 65140
rect 84382 65084 84387 65140
rect 83940 65082 84387 65084
rect 84321 65079 84387 65082
rect 1600 64938 2400 64968
rect 2901 64938 2967 64941
rect 1600 64936 2967 64938
rect 1600 64880 2906 64936
rect 2962 64880 2967 64936
rect 1600 64878 2967 64880
rect 1600 64848 2400 64878
rect 2901 64875 2967 64878
rect 89933 64938 89999 64941
rect 91400 64938 92200 64968
rect 89933 64936 92200 64938
rect 89933 64880 89938 64936
rect 89994 64880 92200 64936
rect 89933 64878 92200 64880
rect 89933 64875 89999 64878
rect 91400 64848 92200 64878
rect 6686 64768 7002 64769
rect 6686 64704 6692 64768
rect 6756 64704 6772 64768
rect 6836 64704 6852 64768
rect 6916 64704 6932 64768
rect 6996 64704 7002 64768
rect 6686 64703 7002 64704
rect 87830 64768 88146 64769
rect 87830 64704 87836 64768
rect 87900 64704 87916 64768
rect 87980 64704 87996 64768
rect 88060 64704 88076 64768
rect 88140 64704 88146 64768
rect 87830 64703 88146 64704
rect 1600 64258 2400 64288
rect 2901 64258 2967 64261
rect 1600 64256 2967 64258
rect 1600 64200 2906 64256
rect 2962 64200 2967 64256
rect 88553 64258 88619 64261
rect 91400 64258 92200 64288
rect 88553 64256 92200 64258
rect 1600 64198 2967 64200
rect 1600 64168 2400 64198
rect 2901 64195 2967 64198
rect 5950 64224 6266 64225
rect 5950 64160 5956 64224
rect 6020 64160 6036 64224
rect 6100 64160 6116 64224
rect 6180 64160 6196 64224
rect 6260 64160 6266 64224
rect 5950 64159 6266 64160
rect 87094 64224 87410 64225
rect 87094 64160 87100 64224
rect 87164 64160 87180 64224
rect 87244 64160 87260 64224
rect 87324 64160 87340 64224
rect 87404 64160 87410 64224
rect 88553 64200 88558 64256
rect 88614 64200 92200 64256
rect 88553 64198 92200 64200
rect 88553 64195 88619 64198
rect 91400 64168 92200 64198
rect 87094 64159 87410 64160
rect 7225 64122 7291 64125
rect 84321 64122 84387 64125
rect 7225 64120 9634 64122
rect 7225 64064 7230 64120
rect 7286 64090 9634 64120
rect 83940 64120 84387 64122
rect 7286 64064 10156 64090
rect 7225 64062 10156 64064
rect 83940 64064 84326 64120
rect 84382 64064 84387 64120
rect 83940 64062 84387 64064
rect 7225 64059 7291 64062
rect 9574 64030 10156 64062
rect 84321 64059 84387 64062
rect 6686 63680 7002 63681
rect 6686 63616 6692 63680
rect 6756 63616 6772 63680
rect 6836 63616 6852 63680
rect 6916 63616 6932 63680
rect 6996 63616 7002 63680
rect 6686 63615 7002 63616
rect 87830 63680 88146 63681
rect 87830 63616 87836 63680
rect 87900 63616 87916 63680
rect 87980 63616 87996 63680
rect 88060 63616 88076 63680
rect 88140 63616 88146 63680
rect 87830 63615 88146 63616
rect 5950 63136 6266 63137
rect 5950 63072 5956 63136
rect 6020 63072 6036 63136
rect 6100 63072 6116 63136
rect 6180 63072 6196 63136
rect 6260 63072 6266 63136
rect 5950 63071 6266 63072
rect 87094 63136 87410 63137
rect 87094 63072 87100 63136
rect 87164 63072 87180 63136
rect 87244 63072 87260 63136
rect 87324 63072 87340 63136
rect 87404 63072 87410 63136
rect 87094 63071 87410 63072
rect 7225 63034 7291 63037
rect 84321 63034 84387 63037
rect 7225 63032 9634 63034
rect 7225 62976 7230 63032
rect 7286 63002 9634 63032
rect 83940 63032 84387 63034
rect 7286 62976 10156 63002
rect 7225 62974 10156 62976
rect 83940 62976 84326 63032
rect 84382 62976 84387 63032
rect 83940 62974 84387 62976
rect 7225 62971 7291 62974
rect 9574 62942 10156 62974
rect 84321 62971 84387 62974
rect 1600 62898 2400 62928
rect 2901 62898 2967 62901
rect 1600 62896 2967 62898
rect 1600 62840 2906 62896
rect 2962 62840 2967 62896
rect 1600 62838 2967 62840
rect 1600 62808 2400 62838
rect 2901 62835 2967 62838
rect 88553 62898 88619 62901
rect 91400 62898 92200 62928
rect 88553 62896 92200 62898
rect 88553 62840 88558 62896
rect 88614 62840 92200 62896
rect 88553 62838 92200 62840
rect 88553 62835 88619 62838
rect 91400 62808 92200 62838
rect 6686 62592 7002 62593
rect 6686 62528 6692 62592
rect 6756 62528 6772 62592
rect 6836 62528 6852 62592
rect 6916 62528 6932 62592
rect 6996 62528 7002 62592
rect 6686 62527 7002 62528
rect 87830 62592 88146 62593
rect 87830 62528 87836 62592
rect 87900 62528 87916 62592
rect 87980 62528 87996 62592
rect 88060 62528 88076 62592
rect 88140 62528 88146 62592
rect 87830 62527 88146 62528
rect 1600 62218 2400 62248
rect 5201 62218 5267 62221
rect 88369 62218 88435 62221
rect 1600 62216 5267 62218
rect 1600 62160 5206 62216
rect 5262 62160 5267 62216
rect 1600 62158 5267 62160
rect 1600 62128 2400 62158
rect 5201 62155 5267 62158
rect 83910 62216 88435 62218
rect 83910 62160 88374 62216
rect 88430 62160 88435 62216
rect 83910 62158 88435 62160
rect 5950 62048 6266 62049
rect 5950 61984 5956 62048
rect 6020 61984 6036 62048
rect 6100 61984 6116 62048
rect 6180 61984 6196 62048
rect 6260 61984 6266 62048
rect 5950 61983 6266 61984
rect 9617 61914 9683 61917
rect 83910 61916 83970 62158
rect 88369 62155 88435 62158
rect 89933 62218 89999 62221
rect 91400 62218 92200 62248
rect 89933 62216 92200 62218
rect 89933 62160 89938 62216
rect 89994 62160 92200 62216
rect 89933 62158 92200 62160
rect 89933 62155 89999 62158
rect 91400 62128 92200 62158
rect 87094 62048 87410 62049
rect 87094 61984 87100 62048
rect 87164 61984 87180 62048
rect 87244 61984 87260 62048
rect 87324 61984 87340 62048
rect 87404 61984 87410 62048
rect 87094 61983 87410 61984
rect 9617 61912 10156 61914
rect 9617 61856 9622 61912
rect 9678 61856 10156 61912
rect 9617 61854 10156 61856
rect 9617 61851 9683 61854
rect 6686 61504 7002 61505
rect 6686 61440 6692 61504
rect 6756 61440 6772 61504
rect 6836 61440 6852 61504
rect 6916 61440 6932 61504
rect 6996 61440 7002 61504
rect 6686 61439 7002 61440
rect 87830 61504 88146 61505
rect 87830 61440 87836 61504
rect 87900 61440 87916 61504
rect 87980 61440 87996 61504
rect 88060 61440 88076 61504
rect 88140 61440 88146 61504
rect 87830 61439 88146 61440
rect 5950 60960 6266 60961
rect 5950 60896 5956 60960
rect 6020 60896 6036 60960
rect 6100 60896 6116 60960
rect 6180 60896 6196 60960
rect 6260 60896 6266 60960
rect 5950 60895 6266 60896
rect 87094 60960 87410 60961
rect 87094 60896 87100 60960
rect 87164 60896 87180 60960
rect 87244 60896 87260 60960
rect 87324 60896 87340 60960
rect 87404 60896 87410 60960
rect 87094 60895 87410 60896
rect 1600 60858 2400 60888
rect 5201 60858 5267 60861
rect 89933 60858 89999 60861
rect 91400 60858 92200 60888
rect 1600 60856 5267 60858
rect 1600 60800 5206 60856
rect 5262 60800 5267 60856
rect 1600 60798 5267 60800
rect 1600 60768 2400 60798
rect 5201 60795 5267 60798
rect 9617 60826 9683 60829
rect 9617 60824 10156 60826
rect 9617 60768 9622 60824
rect 9678 60768 10156 60824
rect 83940 60798 85810 60858
rect 9617 60766 10156 60768
rect 9617 60763 9683 60766
rect 85750 60722 85810 60798
rect 89933 60856 92200 60858
rect 89933 60800 89938 60856
rect 89994 60800 92200 60856
rect 89933 60798 92200 60800
rect 89933 60795 89999 60798
rect 91400 60768 92200 60798
rect 88369 60722 88435 60725
rect 85750 60720 88435 60722
rect 85750 60664 88374 60720
rect 88430 60664 88435 60720
rect 85750 60662 88435 60664
rect 88369 60659 88435 60662
rect 6686 60416 7002 60417
rect 6686 60352 6692 60416
rect 6756 60352 6772 60416
rect 6836 60352 6852 60416
rect 6916 60352 6932 60416
rect 6996 60352 7002 60416
rect 6686 60351 7002 60352
rect 87830 60416 88146 60417
rect 87830 60352 87836 60416
rect 87900 60352 87916 60416
rect 87980 60352 87996 60416
rect 88060 60352 88076 60416
rect 88140 60352 88146 60416
rect 87830 60351 88146 60352
rect 5950 59872 6266 59873
rect 5950 59808 5956 59872
rect 6020 59808 6036 59872
rect 6100 59808 6116 59872
rect 6180 59808 6196 59872
rect 6260 59808 6266 59872
rect 5950 59807 6266 59808
rect 87094 59872 87410 59873
rect 87094 59808 87100 59872
rect 87164 59808 87180 59872
rect 87244 59808 87260 59872
rect 87324 59808 87340 59872
rect 87404 59808 87410 59872
rect 87094 59807 87410 59808
rect 9574 59678 10156 59738
rect 84321 59702 84387 59705
rect 83940 59700 84387 59702
rect 5661 59634 5727 59637
rect 9574 59634 9634 59678
rect 83940 59644 84326 59700
rect 84382 59644 84387 59700
rect 83940 59642 84387 59644
rect 84321 59639 84387 59642
rect 5661 59632 9634 59634
rect 5661 59576 5666 59632
rect 5722 59576 9634 59632
rect 5661 59574 9634 59576
rect 5661 59571 5727 59574
rect 1600 59498 2400 59528
rect 2901 59498 2967 59501
rect 1600 59496 2967 59498
rect 1600 59440 2906 59496
rect 2962 59440 2967 59496
rect 1600 59438 2967 59440
rect 1600 59408 2400 59438
rect 2901 59435 2967 59438
rect 89933 59498 89999 59501
rect 91400 59498 92200 59528
rect 89933 59496 92200 59498
rect 89933 59440 89938 59496
rect 89994 59440 92200 59496
rect 89933 59438 92200 59440
rect 89933 59435 89999 59438
rect 91400 59408 92200 59438
rect 6686 59328 7002 59329
rect 6686 59264 6692 59328
rect 6756 59264 6772 59328
rect 6836 59264 6852 59328
rect 6916 59264 6932 59328
rect 6996 59264 7002 59328
rect 6686 59263 7002 59264
rect 87830 59328 88146 59329
rect 87830 59264 87836 59328
rect 87900 59264 87916 59328
rect 87980 59264 87996 59328
rect 88060 59264 88076 59328
rect 88140 59264 88146 59328
rect 87830 59263 88146 59264
rect 1600 58818 2400 58848
rect 2901 58818 2967 58821
rect 1600 58816 2967 58818
rect 1600 58760 2906 58816
rect 2962 58760 2967 58816
rect 88553 58818 88619 58821
rect 91400 58818 92200 58848
rect 88553 58816 92200 58818
rect 1600 58758 2967 58760
rect 1600 58728 2400 58758
rect 2901 58755 2967 58758
rect 5950 58784 6266 58785
rect 5950 58720 5956 58784
rect 6020 58720 6036 58784
rect 6100 58720 6116 58784
rect 6180 58720 6196 58784
rect 6260 58720 6266 58784
rect 5950 58719 6266 58720
rect 87094 58784 87410 58785
rect 87094 58720 87100 58784
rect 87164 58720 87180 58784
rect 87244 58720 87260 58784
rect 87324 58720 87340 58784
rect 87404 58720 87410 58784
rect 88553 58760 88558 58816
rect 88614 58760 92200 58816
rect 88553 58758 92200 58760
rect 88553 58755 88619 58758
rect 91400 58728 92200 58758
rect 87094 58719 87410 58720
rect 7225 58682 7291 58685
rect 84321 58682 84387 58685
rect 7225 58680 9634 58682
rect 7225 58624 7230 58680
rect 7286 58650 9634 58680
rect 83940 58680 84387 58682
rect 7286 58624 10156 58650
rect 7225 58622 10156 58624
rect 83940 58624 84326 58680
rect 84382 58624 84387 58680
rect 83940 58622 84387 58624
rect 7225 58619 7291 58622
rect 9574 58590 10156 58622
rect 84321 58619 84387 58622
rect 6686 58240 7002 58241
rect 6686 58176 6692 58240
rect 6756 58176 6772 58240
rect 6836 58176 6852 58240
rect 6916 58176 6932 58240
rect 6996 58176 7002 58240
rect 6686 58175 7002 58176
rect 87830 58240 88146 58241
rect 87830 58176 87836 58240
rect 87900 58176 87916 58240
rect 87980 58176 87996 58240
rect 88060 58176 88076 58240
rect 88140 58176 88146 58240
rect 87830 58175 88146 58176
rect 5950 57696 6266 57697
rect 5950 57632 5956 57696
rect 6020 57632 6036 57696
rect 6100 57632 6116 57696
rect 6180 57632 6196 57696
rect 6260 57632 6266 57696
rect 5950 57631 6266 57632
rect 87094 57696 87410 57697
rect 87094 57632 87100 57696
rect 87164 57632 87180 57696
rect 87244 57632 87260 57696
rect 87324 57632 87340 57696
rect 87404 57632 87410 57696
rect 87094 57631 87410 57632
rect 7225 57594 7291 57597
rect 84321 57594 84387 57597
rect 7225 57592 9634 57594
rect 7225 57536 7230 57592
rect 7286 57562 9634 57592
rect 83940 57592 84387 57594
rect 7286 57536 10156 57562
rect 7225 57534 10156 57536
rect 83940 57536 84326 57592
rect 84382 57536 84387 57592
rect 83940 57534 84387 57536
rect 7225 57531 7291 57534
rect 9574 57502 10156 57534
rect 84321 57531 84387 57534
rect 1600 57458 2400 57488
rect 2901 57458 2967 57461
rect 1600 57456 2967 57458
rect 1600 57400 2906 57456
rect 2962 57400 2967 57456
rect 1600 57398 2967 57400
rect 1600 57368 2400 57398
rect 2901 57395 2967 57398
rect 88553 57458 88619 57461
rect 91400 57458 92200 57488
rect 88553 57456 92200 57458
rect 88553 57400 88558 57456
rect 88614 57400 92200 57456
rect 88553 57398 92200 57400
rect 88553 57395 88619 57398
rect 91400 57368 92200 57398
rect 6686 57152 7002 57153
rect 6686 57088 6692 57152
rect 6756 57088 6772 57152
rect 6836 57088 6852 57152
rect 6916 57088 6932 57152
rect 6996 57088 7002 57152
rect 6686 57087 7002 57088
rect 87830 57152 88146 57153
rect 87830 57088 87836 57152
rect 87900 57088 87916 57152
rect 87980 57088 87996 57152
rect 88060 57088 88076 57152
rect 88140 57088 88146 57152
rect 87830 57087 88146 57088
rect 1600 56778 2400 56808
rect 4925 56778 4991 56781
rect 88277 56778 88343 56781
rect 1600 56776 4991 56778
rect 1600 56720 4930 56776
rect 4986 56720 4991 56776
rect 1600 56718 4991 56720
rect 1600 56688 2400 56718
rect 4925 56715 4991 56718
rect 83910 56776 88343 56778
rect 83910 56720 88282 56776
rect 88338 56720 88343 56776
rect 83910 56718 88343 56720
rect 5950 56608 6266 56609
rect 5950 56544 5956 56608
rect 6020 56544 6036 56608
rect 6100 56544 6116 56608
rect 6180 56544 6196 56608
rect 6260 56544 6266 56608
rect 5950 56543 6266 56544
rect 83910 56476 83970 56718
rect 88277 56715 88343 56718
rect 89933 56778 89999 56781
rect 91400 56778 92200 56808
rect 89933 56776 92200 56778
rect 89933 56720 89938 56776
rect 89994 56720 92200 56776
rect 89933 56718 92200 56720
rect 89933 56715 89999 56718
rect 91400 56688 92200 56718
rect 87094 56608 87410 56609
rect 87094 56544 87100 56608
rect 87164 56544 87180 56608
rect 87244 56544 87260 56608
rect 87324 56544 87340 56608
rect 87404 56544 87410 56608
rect 87094 56543 87410 56544
rect 9574 56414 10156 56474
rect 5385 56370 5451 56373
rect 9574 56370 9634 56414
rect 5385 56368 9634 56370
rect 5385 56312 5390 56368
rect 5446 56312 9634 56368
rect 5385 56310 9634 56312
rect 5385 56307 5451 56310
rect 6686 56064 7002 56065
rect 6686 56000 6692 56064
rect 6756 56000 6772 56064
rect 6836 56000 6852 56064
rect 6916 56000 6932 56064
rect 6996 56000 7002 56064
rect 6686 55999 7002 56000
rect 87830 56064 88146 56065
rect 87830 56000 87836 56064
rect 87900 56000 87916 56064
rect 87980 56000 87996 56064
rect 88060 56000 88076 56064
rect 88140 56000 88146 56064
rect 87830 55999 88146 56000
rect 5950 55520 6266 55521
rect 5950 55456 5956 55520
rect 6020 55456 6036 55520
rect 6100 55456 6116 55520
rect 6180 55456 6196 55520
rect 6260 55456 6266 55520
rect 5950 55455 6266 55456
rect 87094 55520 87410 55521
rect 87094 55456 87100 55520
rect 87164 55456 87180 55520
rect 87244 55456 87260 55520
rect 87324 55456 87340 55520
rect 87404 55456 87410 55520
rect 87094 55455 87410 55456
rect 1600 55418 2400 55448
rect 5017 55418 5083 55421
rect 89933 55418 89999 55421
rect 91400 55418 92200 55448
rect 1600 55416 5083 55418
rect 1600 55360 5022 55416
rect 5078 55360 5083 55416
rect 1600 55358 5083 55360
rect 1600 55328 2400 55358
rect 5017 55355 5083 55358
rect 9574 55326 10156 55386
rect 83940 55358 85810 55418
rect 5661 55282 5727 55285
rect 9574 55282 9634 55326
rect 5661 55280 9634 55282
rect 5661 55224 5666 55280
rect 5722 55224 9634 55280
rect 5661 55222 9634 55224
rect 85750 55282 85810 55358
rect 89933 55416 92200 55418
rect 89933 55360 89938 55416
rect 89994 55360 92200 55416
rect 89933 55358 92200 55360
rect 89933 55355 89999 55358
rect 91400 55328 92200 55358
rect 88369 55282 88435 55285
rect 85750 55280 88435 55282
rect 85750 55224 88374 55280
rect 88430 55224 88435 55280
rect 85750 55222 88435 55224
rect 5661 55219 5727 55222
rect 88369 55219 88435 55222
rect 6686 54976 7002 54977
rect 6686 54912 6692 54976
rect 6756 54912 6772 54976
rect 6836 54912 6852 54976
rect 6916 54912 6932 54976
rect 6996 54912 7002 54976
rect 6686 54911 7002 54912
rect 87830 54976 88146 54977
rect 87830 54912 87836 54976
rect 87900 54912 87916 54976
rect 87980 54912 87996 54976
rect 88060 54912 88076 54976
rect 88140 54912 88146 54976
rect 87830 54911 88146 54912
rect 1600 54738 2400 54768
rect 2533 54738 2599 54741
rect 1600 54736 2599 54738
rect 1600 54680 2538 54736
rect 2594 54680 2599 54736
rect 1600 54678 2599 54680
rect 1600 54648 2400 54678
rect 2533 54675 2599 54678
rect 5950 54432 6266 54433
rect 5950 54368 5956 54432
rect 6020 54368 6036 54432
rect 6100 54368 6116 54432
rect 6180 54368 6196 54432
rect 6260 54368 6266 54432
rect 5950 54367 6266 54368
rect 87094 54432 87410 54433
rect 87094 54368 87100 54432
rect 87164 54368 87180 54432
rect 87244 54368 87260 54432
rect 87324 54368 87340 54432
rect 87404 54368 87410 54432
rect 87094 54367 87410 54368
rect 9574 54238 10156 54298
rect 84321 54262 84387 54265
rect 83940 54260 84387 54262
rect 5661 54194 5727 54197
rect 9574 54194 9634 54238
rect 83940 54204 84326 54260
rect 84382 54204 84387 54260
rect 83940 54202 84387 54204
rect 84321 54199 84387 54202
rect 5661 54192 9634 54194
rect 5661 54136 5666 54192
rect 5722 54136 9634 54192
rect 5661 54134 9634 54136
rect 5661 54131 5727 54134
rect 1600 54058 2400 54088
rect 5201 54058 5267 54061
rect 1600 54056 5267 54058
rect 1600 54000 5206 54056
rect 5262 54000 5267 54056
rect 1600 53998 5267 54000
rect 1600 53968 2400 53998
rect 5201 53995 5267 53998
rect 89933 54058 89999 54061
rect 91400 54058 92200 54088
rect 89933 54056 92200 54058
rect 89933 54000 89938 54056
rect 89994 54000 92200 54056
rect 89933 53998 92200 54000
rect 89933 53995 89999 53998
rect 91400 53968 92200 53998
rect 6686 53888 7002 53889
rect 6686 53824 6692 53888
rect 6756 53824 6772 53888
rect 6836 53824 6852 53888
rect 6916 53824 6932 53888
rect 6996 53824 7002 53888
rect 6686 53823 7002 53824
rect 87830 53888 88146 53889
rect 87830 53824 87836 53888
rect 87900 53824 87916 53888
rect 87980 53824 87996 53888
rect 88060 53824 88076 53888
rect 88140 53824 88146 53888
rect 87830 53823 88146 53824
rect 1600 53378 2400 53408
rect 2901 53378 2967 53381
rect 1600 53376 2967 53378
rect 1600 53320 2906 53376
rect 2962 53320 2967 53376
rect 88553 53378 88619 53381
rect 91400 53378 92200 53408
rect 88553 53376 92200 53378
rect 1600 53318 2967 53320
rect 1600 53288 2400 53318
rect 2901 53315 2967 53318
rect 5950 53344 6266 53345
rect 5950 53280 5956 53344
rect 6020 53280 6036 53344
rect 6100 53280 6116 53344
rect 6180 53280 6196 53344
rect 6260 53280 6266 53344
rect 5950 53279 6266 53280
rect 87094 53344 87410 53345
rect 87094 53280 87100 53344
rect 87164 53280 87180 53344
rect 87244 53280 87260 53344
rect 87324 53280 87340 53344
rect 87404 53280 87410 53344
rect 88553 53320 88558 53376
rect 88614 53320 92200 53376
rect 88553 53318 92200 53320
rect 88553 53315 88619 53318
rect 91400 53288 92200 53318
rect 87094 53279 87410 53280
rect 7133 53242 7199 53245
rect 84321 53242 84387 53245
rect 7133 53240 9634 53242
rect 7133 53184 7138 53240
rect 7194 53210 9634 53240
rect 83940 53240 84387 53242
rect 7194 53184 10156 53210
rect 7133 53182 10156 53184
rect 83940 53184 84326 53240
rect 84382 53184 84387 53240
rect 83940 53182 84387 53184
rect 7133 53179 7199 53182
rect 9574 53150 10156 53182
rect 84321 53179 84387 53182
rect 6686 52800 7002 52801
rect 6686 52736 6692 52800
rect 6756 52736 6772 52800
rect 6836 52736 6852 52800
rect 6916 52736 6932 52800
rect 6996 52736 7002 52800
rect 6686 52735 7002 52736
rect 87830 52800 88146 52801
rect 87830 52736 87836 52800
rect 87900 52736 87916 52800
rect 87980 52736 87996 52800
rect 88060 52736 88076 52800
rect 88140 52736 88146 52800
rect 87830 52735 88146 52736
rect 1600 52698 2400 52728
rect 2901 52698 2967 52701
rect 1600 52696 2967 52698
rect 1600 52640 2906 52696
rect 2962 52640 2967 52696
rect 1600 52638 2967 52640
rect 1600 52608 2400 52638
rect 2901 52635 2967 52638
rect 89933 52698 89999 52701
rect 91400 52698 92200 52728
rect 89933 52696 92200 52698
rect 89933 52640 89938 52696
rect 89994 52640 92200 52696
rect 89933 52638 92200 52640
rect 89933 52635 89999 52638
rect 91400 52608 92200 52638
rect 5950 52256 6266 52257
rect 5950 52192 5956 52256
rect 6020 52192 6036 52256
rect 6100 52192 6116 52256
rect 6180 52192 6196 52256
rect 6260 52192 6266 52256
rect 5950 52191 6266 52192
rect 87094 52256 87410 52257
rect 87094 52192 87100 52256
rect 87164 52192 87180 52256
rect 87244 52192 87260 52256
rect 87324 52192 87340 52256
rect 87404 52192 87410 52256
rect 87094 52191 87410 52192
rect 7133 52154 7199 52157
rect 84321 52154 84387 52157
rect 7133 52152 9634 52154
rect 7133 52096 7138 52152
rect 7194 52122 9634 52152
rect 83940 52152 84387 52154
rect 7194 52096 10156 52122
rect 7133 52094 10156 52096
rect 83940 52096 84326 52152
rect 84382 52096 84387 52152
rect 83940 52094 84387 52096
rect 7133 52091 7199 52094
rect 9574 52062 10156 52094
rect 84321 52091 84387 52094
rect 1600 52018 2400 52048
rect 2901 52018 2967 52021
rect 1600 52016 2967 52018
rect 1600 51960 2906 52016
rect 2962 51960 2967 52016
rect 1600 51958 2967 51960
rect 1600 51928 2400 51958
rect 2901 51955 2967 51958
rect 88553 52018 88619 52021
rect 91400 52018 92200 52048
rect 88553 52016 92200 52018
rect 88553 51960 88558 52016
rect 88614 51960 92200 52016
rect 88553 51958 92200 51960
rect 88553 51955 88619 51958
rect 91400 51928 92200 51958
rect 6686 51712 7002 51713
rect 6686 51648 6692 51712
rect 6756 51648 6772 51712
rect 6836 51648 6852 51712
rect 6916 51648 6932 51712
rect 6996 51648 7002 51712
rect 6686 51647 7002 51648
rect 87830 51712 88146 51713
rect 87830 51648 87836 51712
rect 87900 51648 87916 51712
rect 87980 51648 87996 51712
rect 88060 51648 88076 51712
rect 88140 51648 88146 51712
rect 87830 51647 88146 51648
rect 1600 51338 2400 51368
rect 2901 51338 2967 51341
rect 1600 51336 2967 51338
rect 1600 51280 2906 51336
rect 2962 51280 2967 51336
rect 1600 51278 2967 51280
rect 1600 51248 2400 51278
rect 2901 51275 2967 51278
rect 88553 51338 88619 51341
rect 91400 51338 92200 51368
rect 88553 51336 92200 51338
rect 88553 51280 88558 51336
rect 88614 51280 92200 51336
rect 88553 51278 92200 51280
rect 88553 51275 88619 51278
rect 91400 51248 92200 51278
rect 5950 51168 6266 51169
rect 5950 51104 5956 51168
rect 6020 51104 6036 51168
rect 6100 51104 6116 51168
rect 6180 51104 6196 51168
rect 6260 51104 6266 51168
rect 5950 51103 6266 51104
rect 87094 51168 87410 51169
rect 87094 51104 87100 51168
rect 87164 51104 87180 51168
rect 87244 51104 87260 51168
rect 87324 51104 87340 51168
rect 87404 51104 87410 51168
rect 87094 51103 87410 51104
rect 9574 50974 10156 51034
rect 83940 51006 85810 51066
rect 5661 50930 5727 50933
rect 9574 50930 9634 50974
rect 5661 50928 9634 50930
rect 5661 50872 5666 50928
rect 5722 50872 9634 50928
rect 5661 50870 9634 50872
rect 85750 50930 85810 51006
rect 88369 50930 88435 50933
rect 85750 50928 88435 50930
rect 85750 50872 88374 50928
rect 88430 50872 88435 50928
rect 85750 50870 88435 50872
rect 5661 50867 5727 50870
rect 88369 50867 88435 50870
rect 6686 50624 7002 50625
rect 6686 50560 6692 50624
rect 6756 50560 6772 50624
rect 6836 50560 6852 50624
rect 6916 50560 6932 50624
rect 6996 50560 7002 50624
rect 6686 50559 7002 50560
rect 87830 50624 88146 50625
rect 87830 50560 87836 50624
rect 87900 50560 87916 50624
rect 87980 50560 87996 50624
rect 88060 50560 88076 50624
rect 88140 50560 88146 50624
rect 87830 50559 88146 50560
rect 5950 50080 6266 50081
rect 5950 50016 5956 50080
rect 6020 50016 6036 50080
rect 6100 50016 6116 50080
rect 6180 50016 6196 50080
rect 6260 50016 6266 50080
rect 5950 50015 6266 50016
rect 87094 50080 87410 50081
rect 87094 50016 87100 50080
rect 87164 50016 87180 50080
rect 87244 50016 87260 50080
rect 87324 50016 87340 50080
rect 87404 50016 87410 50080
rect 87094 50015 87410 50016
rect 6686 49536 7002 49537
rect 6686 49472 6692 49536
rect 6756 49472 6772 49536
rect 6836 49472 6852 49536
rect 6916 49472 6932 49536
rect 6996 49472 7002 49536
rect 6686 49471 7002 49472
rect 87830 49536 88146 49537
rect 87830 49472 87836 49536
rect 87900 49472 87916 49536
rect 87980 49472 87996 49536
rect 88060 49472 88076 49536
rect 88140 49472 88146 49536
rect 87830 49471 88146 49472
rect 1600 49298 2400 49328
rect 2901 49298 2967 49301
rect 1600 49296 2967 49298
rect 1600 49240 2906 49296
rect 2962 49240 2967 49296
rect 1600 49238 2967 49240
rect 1600 49208 2400 49238
rect 2901 49235 2967 49238
rect 89933 49298 89999 49301
rect 91400 49298 92200 49328
rect 89933 49296 92200 49298
rect 89933 49240 89938 49296
rect 89994 49240 92200 49296
rect 89933 49238 92200 49240
rect 89933 49235 89999 49238
rect 91400 49208 92200 49238
rect 5950 48992 6266 48993
rect 5950 48928 5956 48992
rect 6020 48928 6036 48992
rect 6100 48928 6116 48992
rect 6180 48928 6196 48992
rect 6260 48928 6266 48992
rect 5950 48927 6266 48928
rect 87094 48992 87410 48993
rect 87094 48928 87100 48992
rect 87164 48928 87180 48992
rect 87244 48928 87260 48992
rect 87324 48928 87340 48992
rect 87404 48928 87410 48992
rect 87094 48927 87410 48928
rect 89933 48618 89999 48621
rect 91400 48618 92200 48648
rect 89933 48616 92200 48618
rect 89933 48560 89938 48616
rect 89994 48560 92200 48616
rect 89933 48558 92200 48560
rect 89933 48555 89999 48558
rect 91400 48528 92200 48558
rect 6686 48448 7002 48449
rect 6686 48384 6692 48448
rect 6756 48384 6772 48448
rect 6836 48384 6852 48448
rect 6916 48384 6932 48448
rect 6996 48384 7002 48448
rect 6686 48383 7002 48384
rect 87830 48448 88146 48449
rect 87830 48384 87836 48448
rect 87900 48384 87916 48448
rect 87980 48384 87996 48448
rect 88060 48384 88076 48448
rect 88140 48384 88146 48448
rect 87830 48383 88146 48384
rect 9801 48074 9867 48077
rect 11117 48074 11183 48077
rect 9801 48072 11183 48074
rect 9801 48016 9806 48072
rect 9862 48016 11122 48072
rect 11178 48016 11183 48072
rect 9801 48014 11183 48016
rect 9801 48011 9867 48014
rect 11117 48011 11183 48014
rect 88553 47938 88619 47941
rect 91400 47938 92200 47968
rect 88553 47936 92200 47938
rect 5950 47904 6266 47905
rect 5950 47840 5956 47904
rect 6020 47840 6036 47904
rect 6100 47840 6116 47904
rect 6180 47840 6196 47904
rect 6260 47840 6266 47904
rect 5950 47839 6266 47840
rect 87094 47904 87410 47905
rect 87094 47840 87100 47904
rect 87164 47840 87180 47904
rect 87244 47840 87260 47904
rect 87324 47840 87340 47904
rect 87404 47840 87410 47904
rect 88553 47880 88558 47936
rect 88614 47880 92200 47936
rect 88553 47878 92200 47880
rect 88553 47875 88619 47878
rect 91400 47848 92200 47878
rect 87094 47839 87410 47840
rect 6686 47360 7002 47361
rect 6686 47296 6692 47360
rect 6756 47296 6772 47360
rect 6836 47296 6852 47360
rect 6916 47296 6932 47360
rect 6996 47296 7002 47360
rect 6686 47295 7002 47296
rect 87830 47360 88146 47361
rect 87830 47296 87836 47360
rect 87900 47296 87916 47360
rect 87980 47296 87996 47360
rect 88060 47296 88076 47360
rect 88140 47296 88146 47360
rect 87830 47295 88146 47296
rect 8329 47258 8395 47261
rect 13325 47258 13391 47261
rect 50327 47258 50393 47261
rect 8329 47256 50393 47258
rect 8329 47200 8334 47256
rect 8390 47200 13330 47256
rect 13386 47200 50332 47256
rect 50388 47200 50393 47256
rect 8329 47198 50393 47200
rect 8329 47195 8395 47198
rect 13325 47195 13391 47198
rect 50327 47195 50393 47198
rect 9801 46850 9867 46853
rect 51431 46850 51497 46853
rect 9801 46848 51497 46850
rect 5950 46816 6266 46817
rect 5950 46752 5956 46816
rect 6020 46752 6036 46816
rect 6100 46752 6116 46816
rect 6180 46752 6196 46816
rect 6260 46752 6266 46816
rect 9801 46792 9806 46848
rect 9862 46792 51436 46848
rect 51492 46792 51497 46848
rect 9801 46790 51497 46792
rect 9801 46787 9867 46790
rect 51431 46787 51497 46790
rect 87094 46816 87410 46817
rect 5950 46751 6266 46752
rect 87094 46752 87100 46816
rect 87164 46752 87180 46816
rect 87244 46752 87260 46816
rect 87324 46752 87340 46816
rect 87404 46752 87410 46816
rect 87094 46751 87410 46752
rect 1600 46578 2400 46608
rect 2901 46578 2967 46581
rect 1600 46576 2967 46578
rect 1600 46520 2906 46576
rect 2962 46520 2967 46576
rect 1600 46518 2967 46520
rect 1600 46488 2400 46518
rect 2901 46515 2967 46518
rect 88553 46578 88619 46581
rect 91400 46578 92200 46608
rect 88553 46576 92200 46578
rect 88553 46520 88558 46576
rect 88614 46520 92200 46576
rect 88553 46518 92200 46520
rect 88553 46515 88619 46518
rect 91400 46488 92200 46518
rect 6686 46272 7002 46273
rect 6686 46208 6692 46272
rect 6756 46208 6772 46272
rect 6836 46208 6852 46272
rect 6916 46208 6932 46272
rect 6996 46208 7002 46272
rect 6686 46207 7002 46208
rect 87830 46272 88146 46273
rect 87830 46208 87836 46272
rect 87900 46208 87916 46272
rect 87980 46208 87996 46272
rect 88060 46208 88076 46272
rect 88140 46208 88146 46272
rect 87830 46207 88146 46208
rect 1600 45898 2400 45928
rect 2901 45898 2967 45901
rect 1600 45896 2967 45898
rect 1600 45840 2906 45896
rect 2962 45840 2967 45896
rect 1600 45838 2967 45840
rect 1600 45808 2400 45838
rect 2901 45835 2967 45838
rect 5950 45728 6266 45729
rect 5950 45664 5956 45728
rect 6020 45664 6036 45728
rect 6100 45664 6116 45728
rect 6180 45664 6196 45728
rect 6260 45664 6266 45728
rect 5950 45663 6266 45664
rect 87094 45728 87410 45729
rect 87094 45664 87100 45728
rect 87164 45664 87180 45728
rect 87244 45664 87260 45728
rect 87324 45664 87340 45728
rect 87404 45664 87410 45728
rect 87094 45663 87410 45664
rect 6686 45184 7002 45185
rect 6686 45120 6692 45184
rect 6756 45120 6772 45184
rect 6836 45120 6852 45184
rect 6916 45120 6932 45184
rect 6996 45120 7002 45184
rect 6686 45119 7002 45120
rect 87830 45184 88146 45185
rect 87830 45120 87836 45184
rect 87900 45120 87916 45184
rect 87980 45120 87996 45184
rect 88060 45120 88076 45184
rect 88140 45120 88146 45184
rect 87830 45119 88146 45120
rect 5950 44640 6266 44641
rect 5950 44576 5956 44640
rect 6020 44576 6036 44640
rect 6100 44576 6116 44640
rect 6180 44576 6196 44640
rect 6260 44576 6266 44640
rect 5950 44575 6266 44576
rect 87094 44640 87410 44641
rect 87094 44576 87100 44640
rect 87164 44576 87180 44640
rect 87244 44576 87260 44640
rect 87324 44576 87340 44640
rect 87404 44576 87410 44640
rect 87094 44575 87410 44576
rect 1600 44538 2400 44568
rect 2533 44538 2599 44541
rect 1600 44536 2599 44538
rect 1600 44480 2538 44536
rect 2594 44480 2599 44536
rect 1600 44478 2599 44480
rect 1600 44448 2400 44478
rect 2533 44475 2599 44478
rect 6686 44096 7002 44097
rect 6686 44032 6692 44096
rect 6756 44032 6772 44096
rect 6836 44032 6852 44096
rect 6916 44032 6932 44096
rect 6996 44032 7002 44096
rect 6686 44031 7002 44032
rect 87830 44096 88146 44097
rect 87830 44032 87836 44096
rect 87900 44032 87916 44096
rect 87980 44032 87996 44096
rect 88060 44032 88076 44096
rect 88140 44032 88146 44096
rect 87830 44031 88146 44032
rect 1600 43858 2400 43888
rect 5201 43858 5267 43861
rect 1600 43856 5267 43858
rect 1600 43800 5206 43856
rect 5262 43800 5267 43856
rect 1600 43798 5267 43800
rect 1600 43768 2400 43798
rect 5201 43795 5267 43798
rect 5950 43552 6266 43553
rect 5950 43488 5956 43552
rect 6020 43488 6036 43552
rect 6100 43488 6116 43552
rect 6180 43488 6196 43552
rect 6260 43488 6266 43552
rect 5950 43487 6266 43488
rect 87094 43552 87410 43553
rect 87094 43488 87100 43552
rect 87164 43488 87180 43552
rect 87244 43488 87260 43552
rect 87324 43488 87340 43552
rect 87404 43488 87410 43552
rect 87094 43487 87410 43488
rect 1600 43178 2400 43208
rect 2901 43178 2967 43181
rect 1600 43176 2967 43178
rect 1600 43120 2906 43176
rect 2962 43120 2967 43176
rect 1600 43118 2967 43120
rect 1600 43088 2400 43118
rect 2901 43115 2967 43118
rect 89933 43178 89999 43181
rect 91400 43178 92200 43208
rect 89933 43176 92200 43178
rect 89933 43120 89938 43176
rect 89994 43120 92200 43176
rect 89933 43118 92200 43120
rect 89933 43115 89999 43118
rect 91400 43088 92200 43118
rect 7133 43042 7199 43045
rect 84321 43042 84387 43045
rect 7133 43040 9818 43042
rect 6686 43008 7002 43009
rect 6686 42944 6692 43008
rect 6756 42944 6772 43008
rect 6836 42944 6852 43008
rect 6916 42944 6932 43008
rect 6996 42944 7002 43008
rect 7133 42984 7138 43040
rect 7194 43010 9818 43040
rect 83940 43040 84387 43042
rect 7194 42984 10156 43010
rect 7133 42982 10156 42984
rect 83940 42984 84326 43040
rect 84382 42984 84387 43040
rect 83940 42982 84387 42984
rect 7133 42979 7199 42982
rect 9758 42950 10156 42982
rect 84321 42979 84387 42982
rect 87830 43008 88146 43009
rect 6686 42943 7002 42944
rect 87830 42944 87836 43008
rect 87900 42944 87916 43008
rect 87980 42944 87996 43008
rect 88060 42944 88076 43008
rect 88140 42944 88146 43008
rect 87830 42943 88146 42944
rect 1600 42498 2400 42528
rect 2901 42498 2967 42501
rect 1600 42496 2967 42498
rect 1600 42440 2906 42496
rect 2962 42440 2967 42496
rect 1600 42438 2967 42440
rect 1600 42408 2400 42438
rect 2901 42435 2967 42438
rect 5950 42464 6266 42465
rect 5950 42400 5956 42464
rect 6020 42400 6036 42464
rect 6100 42400 6116 42464
rect 6180 42400 6196 42464
rect 6260 42400 6266 42464
rect 5950 42399 6266 42400
rect 87094 42464 87410 42465
rect 87094 42400 87100 42464
rect 87164 42400 87180 42464
rect 87244 42400 87260 42464
rect 87324 42400 87340 42464
rect 87404 42400 87410 42464
rect 87094 42399 87410 42400
rect 7133 41954 7199 41957
rect 84321 41954 84387 41957
rect 7133 41952 9634 41954
rect 6686 41920 7002 41921
rect 6686 41856 6692 41920
rect 6756 41856 6772 41920
rect 6836 41856 6852 41920
rect 6916 41856 6932 41920
rect 6996 41856 7002 41920
rect 7133 41896 7138 41952
rect 7194 41922 9634 41952
rect 83940 41952 84387 41954
rect 7194 41896 10156 41922
rect 7133 41894 10156 41896
rect 83940 41896 84326 41952
rect 84382 41896 84387 41952
rect 83940 41894 84387 41896
rect 7133 41891 7199 41894
rect 9574 41862 10156 41894
rect 84321 41891 84387 41894
rect 87830 41920 88146 41921
rect 6686 41855 7002 41856
rect 87830 41856 87836 41920
rect 87900 41856 87916 41920
rect 87980 41856 87996 41920
rect 88060 41856 88076 41920
rect 88140 41856 88146 41920
rect 87830 41855 88146 41856
rect 1600 41818 2400 41848
rect 2901 41818 2967 41821
rect 1600 41816 2967 41818
rect 1600 41760 2906 41816
rect 2962 41760 2967 41816
rect 1600 41758 2967 41760
rect 1600 41728 2400 41758
rect 2901 41755 2967 41758
rect 88553 41818 88619 41821
rect 91400 41818 92200 41848
rect 88553 41816 92200 41818
rect 88553 41760 88558 41816
rect 88614 41760 92200 41816
rect 88553 41758 92200 41760
rect 88553 41755 88619 41758
rect 91400 41728 92200 41758
rect 5950 41376 6266 41377
rect 5950 41312 5956 41376
rect 6020 41312 6036 41376
rect 6100 41312 6116 41376
rect 6180 41312 6196 41376
rect 6260 41312 6266 41376
rect 5950 41311 6266 41312
rect 87094 41376 87410 41377
rect 87094 41312 87100 41376
rect 87164 41312 87180 41376
rect 87244 41312 87260 41376
rect 87324 41312 87340 41376
rect 87404 41312 87410 41376
rect 87094 41311 87410 41312
rect 1600 41138 2400 41168
rect 4373 41138 4439 41141
rect 1600 41136 4439 41138
rect 1600 41080 4378 41136
rect 4434 41080 4439 41136
rect 1600 41078 4439 41080
rect 1600 41048 2400 41078
rect 4373 41075 4439 41078
rect 89933 41138 89999 41141
rect 91400 41138 92200 41168
rect 89933 41136 92200 41138
rect 89933 41080 89938 41136
rect 89994 41080 92200 41136
rect 89933 41078 92200 41080
rect 89933 41075 89999 41078
rect 91400 41048 92200 41078
rect 5661 41002 5727 41005
rect 5661 41000 9634 41002
rect 5661 40944 5666 41000
rect 5722 40944 9634 41000
rect 5661 40942 9634 40944
rect 5661 40939 5727 40942
rect 9574 40834 9634 40942
rect 87449 40866 87515 40869
rect 83940 40864 87515 40866
rect 6686 40832 7002 40833
rect 6686 40768 6692 40832
rect 6756 40768 6772 40832
rect 6836 40768 6852 40832
rect 6916 40768 6932 40832
rect 6996 40768 7002 40832
rect 9574 40774 10156 40834
rect 83940 40808 87454 40864
rect 87510 40808 87515 40864
rect 83940 40806 87515 40808
rect 87449 40803 87515 40806
rect 87830 40832 88146 40833
rect 6686 40767 7002 40768
rect 87830 40768 87836 40832
rect 87900 40768 87916 40832
rect 87980 40768 87996 40832
rect 88060 40768 88076 40832
rect 88140 40768 88146 40832
rect 87830 40767 88146 40768
rect 5950 40288 6266 40289
rect 5950 40224 5956 40288
rect 6020 40224 6036 40288
rect 6100 40224 6116 40288
rect 6180 40224 6196 40288
rect 6260 40224 6266 40288
rect 5950 40223 6266 40224
rect 87094 40288 87410 40289
rect 87094 40224 87100 40288
rect 87164 40224 87180 40288
rect 87244 40224 87260 40288
rect 87324 40224 87340 40288
rect 87404 40224 87410 40288
rect 87094 40223 87410 40224
rect 1600 39778 2400 39808
rect 2901 39778 2967 39781
rect 1600 39776 2967 39778
rect 1600 39720 2906 39776
rect 2962 39720 2967 39776
rect 7133 39778 7199 39781
rect 84321 39778 84387 39781
rect 7133 39776 9634 39778
rect 1600 39718 2967 39720
rect 1600 39688 2400 39718
rect 2901 39715 2967 39718
rect 6686 39744 7002 39745
rect 6686 39680 6692 39744
rect 6756 39680 6772 39744
rect 6836 39680 6852 39744
rect 6916 39680 6932 39744
rect 6996 39680 7002 39744
rect 7133 39720 7138 39776
rect 7194 39746 9634 39776
rect 83940 39776 84387 39778
rect 7194 39720 10156 39746
rect 7133 39718 10156 39720
rect 83940 39720 84326 39776
rect 84382 39720 84387 39776
rect 89933 39778 89999 39781
rect 91400 39778 92200 39808
rect 89933 39776 92200 39778
rect 83940 39718 84387 39720
rect 7133 39715 7199 39718
rect 9574 39686 10156 39718
rect 84321 39715 84387 39718
rect 87830 39744 88146 39745
rect 6686 39679 7002 39680
rect 87830 39680 87836 39744
rect 87900 39680 87916 39744
rect 87980 39680 87996 39744
rect 88060 39680 88076 39744
rect 88140 39680 88146 39744
rect 89933 39720 89938 39776
rect 89994 39720 92200 39776
rect 89933 39718 92200 39720
rect 89933 39715 89999 39718
rect 91400 39688 92200 39718
rect 87830 39679 88146 39680
rect 5950 39200 6266 39201
rect 5950 39136 5956 39200
rect 6020 39136 6036 39200
rect 6100 39136 6116 39200
rect 6180 39136 6196 39200
rect 6260 39136 6266 39200
rect 5950 39135 6266 39136
rect 87094 39200 87410 39201
rect 87094 39136 87100 39200
rect 87164 39136 87180 39200
rect 87244 39136 87260 39200
rect 87324 39136 87340 39200
rect 87404 39136 87410 39200
rect 87094 39135 87410 39136
rect 7409 38690 7475 38693
rect 87173 38690 87239 38693
rect 7409 38688 9634 38690
rect 6686 38656 7002 38657
rect 6686 38592 6692 38656
rect 6756 38592 6772 38656
rect 6836 38592 6852 38656
rect 6916 38592 6932 38656
rect 6996 38592 7002 38656
rect 7409 38632 7414 38688
rect 7470 38658 9634 38688
rect 83940 38688 87239 38690
rect 7470 38632 10156 38658
rect 7409 38630 10156 38632
rect 83940 38632 87178 38688
rect 87234 38632 87239 38688
rect 83940 38630 87239 38632
rect 7409 38627 7475 38630
rect 9574 38598 10156 38630
rect 87173 38627 87239 38630
rect 87830 38656 88146 38657
rect 6686 38591 7002 38592
rect 87830 38592 87836 38656
rect 87900 38592 87916 38656
rect 87980 38592 87996 38656
rect 88060 38592 88076 38656
rect 88140 38592 88146 38656
rect 87830 38591 88146 38592
rect 1600 38418 2400 38448
rect 4373 38418 4439 38421
rect 1600 38416 4439 38418
rect 1600 38360 4378 38416
rect 4434 38360 4439 38416
rect 1600 38358 4439 38360
rect 1600 38328 2400 38358
rect 4373 38355 4439 38358
rect 89289 38418 89355 38421
rect 91400 38418 92200 38448
rect 89289 38416 92200 38418
rect 89289 38360 89294 38416
rect 89350 38360 92200 38416
rect 89289 38358 92200 38360
rect 89289 38355 89355 38358
rect 91400 38328 92200 38358
rect 5950 38112 6266 38113
rect 5950 38048 5956 38112
rect 6020 38048 6036 38112
rect 6100 38048 6116 38112
rect 6180 38048 6196 38112
rect 6260 38048 6266 38112
rect 5950 38047 6266 38048
rect 87094 38112 87410 38113
rect 87094 38048 87100 38112
rect 87164 38048 87180 38112
rect 87244 38048 87260 38112
rect 87324 38048 87340 38112
rect 87404 38048 87410 38112
rect 87094 38047 87410 38048
rect 1600 37738 2400 37768
rect 2901 37738 2967 37741
rect 1600 37736 2967 37738
rect 1600 37680 2906 37736
rect 2962 37680 2967 37736
rect 1600 37678 2967 37680
rect 1600 37648 2400 37678
rect 2901 37675 2967 37678
rect 89933 37738 89999 37741
rect 91400 37738 92200 37768
rect 89933 37736 92200 37738
rect 89933 37680 89938 37736
rect 89994 37680 92200 37736
rect 89933 37678 92200 37680
rect 89933 37675 89999 37678
rect 91400 37648 92200 37678
rect 7133 37602 7199 37605
rect 84321 37602 84387 37605
rect 7133 37600 9634 37602
rect 6686 37568 7002 37569
rect 6686 37504 6692 37568
rect 6756 37504 6772 37568
rect 6836 37504 6852 37568
rect 6916 37504 6932 37568
rect 6996 37504 7002 37568
rect 7133 37544 7138 37600
rect 7194 37570 9634 37600
rect 83940 37600 84387 37602
rect 7194 37544 10156 37570
rect 7133 37542 10156 37544
rect 83940 37544 84326 37600
rect 84382 37544 84387 37600
rect 83940 37542 84387 37544
rect 7133 37539 7199 37542
rect 9574 37510 10156 37542
rect 84321 37539 84387 37542
rect 87830 37568 88146 37569
rect 6686 37503 7002 37504
rect 87830 37504 87836 37568
rect 87900 37504 87916 37568
rect 87980 37504 87996 37568
rect 88060 37504 88076 37568
rect 88140 37504 88146 37568
rect 87830 37503 88146 37504
rect 5950 37024 6266 37025
rect 5950 36960 5956 37024
rect 6020 36960 6036 37024
rect 6100 36960 6116 37024
rect 6180 36960 6196 37024
rect 6260 36960 6266 37024
rect 5950 36959 6266 36960
rect 87094 37024 87410 37025
rect 87094 36960 87100 37024
rect 87164 36960 87180 37024
rect 87244 36960 87260 37024
rect 87324 36960 87340 37024
rect 87404 36960 87410 37024
rect 87094 36959 87410 36960
rect 7133 36514 7199 36517
rect 84321 36514 84387 36517
rect 7133 36512 9634 36514
rect 6686 36480 7002 36481
rect 6686 36416 6692 36480
rect 6756 36416 6772 36480
rect 6836 36416 6852 36480
rect 6916 36416 6932 36480
rect 6996 36416 7002 36480
rect 7133 36456 7138 36512
rect 7194 36482 9634 36512
rect 83940 36512 84387 36514
rect 7194 36456 10156 36482
rect 7133 36454 10156 36456
rect 83940 36456 84326 36512
rect 84382 36456 84387 36512
rect 83940 36454 84387 36456
rect 7133 36451 7199 36454
rect 9574 36422 10156 36454
rect 84321 36451 84387 36454
rect 87830 36480 88146 36481
rect 6686 36415 7002 36416
rect 87830 36416 87836 36480
rect 87900 36416 87916 36480
rect 87980 36416 87996 36480
rect 88060 36416 88076 36480
rect 88140 36416 88146 36480
rect 87830 36415 88146 36416
rect 1600 36378 2400 36408
rect 2901 36378 2967 36381
rect 1600 36376 2967 36378
rect 1600 36320 2906 36376
rect 2962 36320 2967 36376
rect 1600 36318 2967 36320
rect 1600 36288 2400 36318
rect 2901 36315 2967 36318
rect 89933 36378 89999 36381
rect 91400 36378 92200 36408
rect 89933 36376 92200 36378
rect 89933 36320 89938 36376
rect 89994 36320 92200 36376
rect 89933 36318 92200 36320
rect 89933 36315 89999 36318
rect 91400 36288 92200 36318
rect 5950 35936 6266 35937
rect 5950 35872 5956 35936
rect 6020 35872 6036 35936
rect 6100 35872 6116 35936
rect 6180 35872 6196 35936
rect 6260 35872 6266 35936
rect 5950 35871 6266 35872
rect 87094 35936 87410 35937
rect 87094 35872 87100 35936
rect 87164 35872 87180 35936
rect 87244 35872 87260 35936
rect 87324 35872 87340 35936
rect 87404 35872 87410 35936
rect 87094 35871 87410 35872
rect 1600 35698 2400 35728
rect 4373 35698 4439 35701
rect 1600 35696 4439 35698
rect 1600 35640 4378 35696
rect 4434 35640 4439 35696
rect 1600 35638 4439 35640
rect 1600 35608 2400 35638
rect 4373 35635 4439 35638
rect 90117 35698 90183 35701
rect 91400 35698 92200 35728
rect 90117 35696 92200 35698
rect 90117 35640 90122 35696
rect 90178 35640 92200 35696
rect 90117 35638 92200 35640
rect 90117 35635 90183 35638
rect 91400 35608 92200 35638
rect 5661 35562 5727 35565
rect 5661 35560 9634 35562
rect 5661 35504 5666 35560
rect 5722 35504 9634 35560
rect 5661 35502 9634 35504
rect 5661 35499 5727 35502
rect 9574 35394 9634 35502
rect 87449 35426 87515 35429
rect 83940 35424 87515 35426
rect 6686 35392 7002 35393
rect 6686 35328 6692 35392
rect 6756 35328 6772 35392
rect 6836 35328 6852 35392
rect 6916 35328 6932 35392
rect 6996 35328 7002 35392
rect 9574 35334 10156 35394
rect 83940 35368 87454 35424
rect 87510 35368 87515 35424
rect 83940 35366 87515 35368
rect 87449 35363 87515 35366
rect 87830 35392 88146 35393
rect 6686 35327 7002 35328
rect 87830 35328 87836 35392
rect 87900 35328 87916 35392
rect 87980 35328 87996 35392
rect 88060 35328 88076 35392
rect 88140 35328 88146 35392
rect 87830 35327 88146 35328
rect 5950 34848 6266 34849
rect 5950 34784 5956 34848
rect 6020 34784 6036 34848
rect 6100 34784 6116 34848
rect 6180 34784 6196 34848
rect 6260 34784 6266 34848
rect 5950 34783 6266 34784
rect 87094 34848 87410 34849
rect 87094 34784 87100 34848
rect 87164 34784 87180 34848
rect 87244 34784 87260 34848
rect 87324 34784 87340 34848
rect 87404 34784 87410 34848
rect 87094 34783 87410 34784
rect 1600 34338 2400 34368
rect 2901 34338 2967 34341
rect 1600 34336 2967 34338
rect 1600 34280 2906 34336
rect 2962 34280 2967 34336
rect 7133 34338 7199 34341
rect 84321 34338 84387 34341
rect 7133 34336 9634 34338
rect 1600 34278 2967 34280
rect 1600 34248 2400 34278
rect 2901 34275 2967 34278
rect 6686 34304 7002 34305
rect 6686 34240 6692 34304
rect 6756 34240 6772 34304
rect 6836 34240 6852 34304
rect 6916 34240 6932 34304
rect 6996 34240 7002 34304
rect 7133 34280 7138 34336
rect 7194 34306 9634 34336
rect 83940 34336 84387 34338
rect 7194 34280 10156 34306
rect 7133 34278 10156 34280
rect 83940 34280 84326 34336
rect 84382 34280 84387 34336
rect 88553 34338 88619 34341
rect 91400 34338 92200 34368
rect 88553 34336 92200 34338
rect 83940 34278 84387 34280
rect 7133 34275 7199 34278
rect 9574 34246 10156 34278
rect 84321 34275 84387 34278
rect 87830 34304 88146 34305
rect 6686 34239 7002 34240
rect 87830 34240 87836 34304
rect 87900 34240 87916 34304
rect 87980 34240 87996 34304
rect 88060 34240 88076 34304
rect 88140 34240 88146 34304
rect 88553 34280 88558 34336
rect 88614 34280 92200 34336
rect 88553 34278 92200 34280
rect 88553 34275 88619 34278
rect 91400 34248 92200 34278
rect 87830 34239 88146 34240
rect 5950 33760 6266 33761
rect 5950 33696 5956 33760
rect 6020 33696 6036 33760
rect 6100 33696 6116 33760
rect 6180 33696 6196 33760
rect 6260 33696 6266 33760
rect 5950 33695 6266 33696
rect 87094 33760 87410 33761
rect 87094 33696 87100 33760
rect 87164 33696 87180 33760
rect 87244 33696 87260 33760
rect 87324 33696 87340 33760
rect 87404 33696 87410 33760
rect 87094 33695 87410 33696
rect 1600 33658 2400 33688
rect 2901 33658 2967 33661
rect 1600 33656 2967 33658
rect 1600 33600 2906 33656
rect 2962 33600 2967 33656
rect 1600 33598 2967 33600
rect 1600 33568 2400 33598
rect 2901 33595 2967 33598
rect 87173 33250 87239 33253
rect 83940 33248 87239 33250
rect 6686 33216 7002 33217
rect 6686 33152 6692 33216
rect 6756 33152 6772 33216
rect 6836 33152 6852 33216
rect 6916 33152 6932 33216
rect 6996 33152 7002 33216
rect 6686 33151 7002 33152
rect 9574 33158 10156 33218
rect 83940 33192 87178 33248
rect 87234 33192 87239 33248
rect 83940 33190 87239 33192
rect 87173 33187 87239 33190
rect 87830 33216 88146 33217
rect 1600 32978 2400 33008
rect 4373 32978 4439 32981
rect 1600 32976 4439 32978
rect 1600 32920 4378 32976
rect 4434 32920 4439 32976
rect 1600 32918 4439 32920
rect 1600 32888 2400 32918
rect 4373 32915 4439 32918
rect 5661 32978 5727 32981
rect 9574 32978 9634 33158
rect 87830 33152 87836 33216
rect 87900 33152 87916 33216
rect 87980 33152 87996 33216
rect 88060 33152 88076 33216
rect 88140 33152 88146 33216
rect 87830 33151 88146 33152
rect 5661 32976 9634 32978
rect 5661 32920 5666 32976
rect 5722 32920 9634 32976
rect 5661 32918 9634 32920
rect 89933 32978 89999 32981
rect 91400 32978 92200 33008
rect 89933 32976 92200 32978
rect 89933 32920 89938 32976
rect 89994 32920 92200 32976
rect 89933 32918 92200 32920
rect 5661 32915 5727 32918
rect 89933 32915 89999 32918
rect 91400 32888 92200 32918
rect 5950 32672 6266 32673
rect 5950 32608 5956 32672
rect 6020 32608 6036 32672
rect 6100 32608 6116 32672
rect 6180 32608 6196 32672
rect 6260 32608 6266 32672
rect 5950 32607 6266 32608
rect 87094 32672 87410 32673
rect 87094 32608 87100 32672
rect 87164 32608 87180 32672
rect 87244 32608 87260 32672
rect 87324 32608 87340 32672
rect 87404 32608 87410 32672
rect 87094 32607 87410 32608
rect 1600 32298 2400 32328
rect 2901 32298 2967 32301
rect 1600 32296 2967 32298
rect 1600 32240 2906 32296
rect 2962 32240 2967 32296
rect 1600 32238 2967 32240
rect 1600 32208 2400 32238
rect 2901 32235 2967 32238
rect 89933 32298 89999 32301
rect 91400 32298 92200 32328
rect 89933 32296 92200 32298
rect 89933 32240 89938 32296
rect 89994 32240 92200 32296
rect 89933 32238 92200 32240
rect 89933 32235 89999 32238
rect 91400 32208 92200 32238
rect 7133 32162 7199 32165
rect 84321 32162 84387 32165
rect 7133 32160 9634 32162
rect 6686 32128 7002 32129
rect 6686 32064 6692 32128
rect 6756 32064 6772 32128
rect 6836 32064 6852 32128
rect 6916 32064 6932 32128
rect 6996 32064 7002 32128
rect 7133 32104 7138 32160
rect 7194 32130 9634 32160
rect 83940 32160 84387 32162
rect 7194 32104 10156 32130
rect 7133 32102 10156 32104
rect 83940 32104 84326 32160
rect 84382 32104 84387 32160
rect 83940 32102 84387 32104
rect 7133 32099 7199 32102
rect 9574 32070 10156 32102
rect 84321 32099 84387 32102
rect 87830 32128 88146 32129
rect 6686 32063 7002 32064
rect 87830 32064 87836 32128
rect 87900 32064 87916 32128
rect 87980 32064 87996 32128
rect 88060 32064 88076 32128
rect 88140 32064 88146 32128
rect 87830 32063 88146 32064
rect 5950 31584 6266 31585
rect 5950 31520 5956 31584
rect 6020 31520 6036 31584
rect 6100 31520 6116 31584
rect 6180 31520 6196 31584
rect 6260 31520 6266 31584
rect 5950 31519 6266 31520
rect 87094 31584 87410 31585
rect 87094 31520 87100 31584
rect 87164 31520 87180 31584
rect 87244 31520 87260 31584
rect 87324 31520 87340 31584
rect 87404 31520 87410 31584
rect 87094 31519 87410 31520
rect 7133 31074 7199 31077
rect 84321 31074 84387 31077
rect 7133 31072 9634 31074
rect 6686 31040 7002 31041
rect 6686 30976 6692 31040
rect 6756 30976 6772 31040
rect 6836 30976 6852 31040
rect 6916 30976 6932 31040
rect 6996 30976 7002 31040
rect 7133 31016 7138 31072
rect 7194 31042 9634 31072
rect 83940 31072 84387 31074
rect 7194 31016 10156 31042
rect 7133 31014 10156 31016
rect 83940 31016 84326 31072
rect 84382 31016 84387 31072
rect 83940 31014 84387 31016
rect 7133 31011 7199 31014
rect 9574 30982 10156 31014
rect 84321 31011 84387 31014
rect 87830 31040 88146 31041
rect 6686 30975 7002 30976
rect 87830 30976 87836 31040
rect 87900 30976 87916 31040
rect 87980 30976 87996 31040
rect 88060 30976 88076 31040
rect 88140 30976 88146 31040
rect 87830 30975 88146 30976
rect 1600 30938 2400 30968
rect 2901 30938 2967 30941
rect 1600 30936 2967 30938
rect 1600 30880 2906 30936
rect 2962 30880 2967 30936
rect 1600 30878 2967 30880
rect 1600 30848 2400 30878
rect 2901 30875 2967 30878
rect 88553 30938 88619 30941
rect 91400 30938 92200 30968
rect 88553 30936 92200 30938
rect 88553 30880 88558 30936
rect 88614 30880 92200 30936
rect 88553 30878 92200 30880
rect 88553 30875 88619 30878
rect 91400 30848 92200 30878
rect 5950 30496 6266 30497
rect 5950 30432 5956 30496
rect 6020 30432 6036 30496
rect 6100 30432 6116 30496
rect 6180 30432 6196 30496
rect 6260 30432 6266 30496
rect 5950 30431 6266 30432
rect 87094 30496 87410 30497
rect 87094 30432 87100 30496
rect 87164 30432 87180 30496
rect 87244 30432 87260 30496
rect 87324 30432 87340 30496
rect 87404 30432 87410 30496
rect 87094 30431 87410 30432
rect 1600 30258 2400 30288
rect 4373 30258 4439 30261
rect 87449 30258 87515 30261
rect 1600 30256 4439 30258
rect 1600 30200 4378 30256
rect 4434 30200 4439 30256
rect 1600 30198 4439 30200
rect 1600 30168 2400 30198
rect 4373 30195 4439 30198
rect 83910 30256 87515 30258
rect 83910 30200 87454 30256
rect 87510 30200 87515 30256
rect 83910 30198 87515 30200
rect 5661 30122 5727 30125
rect 5661 30120 9634 30122
rect 5661 30064 5666 30120
rect 5722 30064 9634 30120
rect 5661 30062 9634 30064
rect 5661 30059 5727 30062
rect 9574 29954 9634 30062
rect 83910 29956 83970 30198
rect 87449 30195 87515 30198
rect 89933 30258 89999 30261
rect 91400 30258 92200 30288
rect 89933 30256 92200 30258
rect 89933 30200 89938 30256
rect 89994 30200 92200 30256
rect 89933 30198 92200 30200
rect 89933 30195 89999 30198
rect 91400 30168 92200 30198
rect 6686 29952 7002 29953
rect 6686 29888 6692 29952
rect 6756 29888 6772 29952
rect 6836 29888 6852 29952
rect 6916 29888 6932 29952
rect 6996 29888 7002 29952
rect 9574 29894 10156 29954
rect 87830 29952 88146 29953
rect 6686 29887 7002 29888
rect 87830 29888 87836 29952
rect 87900 29888 87916 29952
rect 87980 29888 87996 29952
rect 88060 29888 88076 29952
rect 88140 29888 88146 29952
rect 87830 29887 88146 29888
rect 5950 29408 6266 29409
rect 5950 29344 5956 29408
rect 6020 29344 6036 29408
rect 6100 29344 6116 29408
rect 6180 29344 6196 29408
rect 6260 29344 6266 29408
rect 5950 29343 6266 29344
rect 87094 29408 87410 29409
rect 87094 29344 87100 29408
rect 87164 29344 87180 29408
rect 87244 29344 87260 29408
rect 87324 29344 87340 29408
rect 87404 29344 87410 29408
rect 87094 29343 87410 29344
rect 1600 28898 2400 28928
rect 2901 28898 2967 28901
rect 1600 28896 2967 28898
rect 1600 28840 2906 28896
rect 2962 28840 2967 28896
rect 7133 28898 7199 28901
rect 84321 28898 84387 28901
rect 7133 28896 9634 28898
rect 1600 28838 2967 28840
rect 1600 28808 2400 28838
rect 2901 28835 2967 28838
rect 6686 28864 7002 28865
rect 6686 28800 6692 28864
rect 6756 28800 6772 28864
rect 6836 28800 6852 28864
rect 6916 28800 6932 28864
rect 6996 28800 7002 28864
rect 7133 28840 7138 28896
rect 7194 28866 9634 28896
rect 83940 28896 84387 28898
rect 7194 28840 10156 28866
rect 7133 28838 10156 28840
rect 83940 28840 84326 28896
rect 84382 28840 84387 28896
rect 88553 28898 88619 28901
rect 91400 28898 92200 28928
rect 88553 28896 92200 28898
rect 83940 28838 84387 28840
rect 7133 28835 7199 28838
rect 9574 28806 10156 28838
rect 84321 28835 84387 28838
rect 87830 28864 88146 28865
rect 6686 28799 7002 28800
rect 87830 28800 87836 28864
rect 87900 28800 87916 28864
rect 87980 28800 87996 28864
rect 88060 28800 88076 28864
rect 88140 28800 88146 28864
rect 88553 28840 88558 28896
rect 88614 28840 92200 28896
rect 88553 28838 92200 28840
rect 88553 28835 88619 28838
rect 91400 28808 92200 28838
rect 87830 28799 88146 28800
rect 5950 28320 6266 28321
rect 5950 28256 5956 28320
rect 6020 28256 6036 28320
rect 6100 28256 6116 28320
rect 6180 28256 6196 28320
rect 6260 28256 6266 28320
rect 5950 28255 6266 28256
rect 87094 28320 87410 28321
rect 87094 28256 87100 28320
rect 87164 28256 87180 28320
rect 87244 28256 87260 28320
rect 87324 28256 87340 28320
rect 87404 28256 87410 28320
rect 87094 28255 87410 28256
rect 87541 27810 87607 27813
rect 83940 27808 87607 27810
rect 6686 27776 7002 27777
rect 6686 27712 6692 27776
rect 6756 27712 6772 27776
rect 6836 27712 6852 27776
rect 6916 27712 6932 27776
rect 6996 27712 7002 27776
rect 6686 27711 7002 27712
rect 9574 27718 10156 27778
rect 83940 27752 87546 27808
rect 87602 27752 87607 27808
rect 83940 27750 87607 27752
rect 87541 27747 87607 27750
rect 87830 27776 88146 27777
rect 1600 27538 2400 27568
rect 5109 27538 5175 27541
rect 1600 27536 5175 27538
rect 1600 27480 5114 27536
rect 5170 27480 5175 27536
rect 1600 27478 5175 27480
rect 1600 27448 2400 27478
rect 5109 27475 5175 27478
rect 5385 27538 5451 27541
rect 9574 27538 9634 27718
rect 87830 27712 87836 27776
rect 87900 27712 87916 27776
rect 87980 27712 87996 27776
rect 88060 27712 88076 27776
rect 88140 27712 88146 27776
rect 87830 27711 88146 27712
rect 5385 27536 9634 27538
rect 5385 27480 5390 27536
rect 5446 27480 9634 27536
rect 5385 27478 9634 27480
rect 89933 27538 89999 27541
rect 91400 27538 92200 27568
rect 89933 27536 92200 27538
rect 89933 27480 89938 27536
rect 89994 27480 92200 27536
rect 89933 27478 92200 27480
rect 5385 27475 5451 27478
rect 89933 27475 89999 27478
rect 91400 27448 92200 27478
rect 5950 27232 6266 27233
rect 5950 27168 5956 27232
rect 6020 27168 6036 27232
rect 6100 27168 6116 27232
rect 6180 27168 6196 27232
rect 6260 27168 6266 27232
rect 5950 27167 6266 27168
rect 87094 27232 87410 27233
rect 87094 27168 87100 27232
rect 87164 27168 87180 27232
rect 87244 27168 87260 27232
rect 87324 27168 87340 27232
rect 87404 27168 87410 27232
rect 87094 27167 87410 27168
rect 1600 26858 2400 26888
rect 2901 26858 2967 26861
rect 1600 26856 2967 26858
rect 1600 26800 2906 26856
rect 2962 26800 2967 26856
rect 1600 26798 2967 26800
rect 1600 26768 2400 26798
rect 2901 26795 2967 26798
rect 89933 26858 89999 26861
rect 91400 26858 92200 26888
rect 89933 26856 92200 26858
rect 89933 26800 89938 26856
rect 89994 26800 92200 26856
rect 89933 26798 92200 26800
rect 89933 26795 89999 26798
rect 91400 26768 92200 26798
rect 7133 26722 7199 26725
rect 84321 26722 84387 26725
rect 7133 26720 9634 26722
rect 6686 26688 7002 26689
rect 6686 26624 6692 26688
rect 6756 26624 6772 26688
rect 6836 26624 6852 26688
rect 6916 26624 6932 26688
rect 6996 26624 7002 26688
rect 7133 26664 7138 26720
rect 7194 26690 9634 26720
rect 83940 26720 84387 26722
rect 7194 26664 10156 26690
rect 7133 26662 10156 26664
rect 83940 26664 84326 26720
rect 84382 26664 84387 26720
rect 83940 26662 84387 26664
rect 7133 26659 7199 26662
rect 9574 26630 10156 26662
rect 84321 26659 84387 26662
rect 87830 26688 88146 26689
rect 6686 26623 7002 26624
rect 87830 26624 87836 26688
rect 87900 26624 87916 26688
rect 87980 26624 87996 26688
rect 88060 26624 88076 26688
rect 88140 26624 88146 26688
rect 87830 26623 88146 26624
rect 5950 26144 6266 26145
rect 5950 26080 5956 26144
rect 6020 26080 6036 26144
rect 6100 26080 6116 26144
rect 6180 26080 6196 26144
rect 6260 26080 6266 26144
rect 5950 26079 6266 26080
rect 87094 26144 87410 26145
rect 87094 26080 87100 26144
rect 87164 26080 87180 26144
rect 87244 26080 87260 26144
rect 87324 26080 87340 26144
rect 87404 26080 87410 26144
rect 87094 26079 87410 26080
rect 7133 25634 7199 25637
rect 84321 25634 84387 25637
rect 7133 25632 9634 25634
rect 6686 25600 7002 25601
rect 6686 25536 6692 25600
rect 6756 25536 6772 25600
rect 6836 25536 6852 25600
rect 6916 25536 6932 25600
rect 6996 25536 7002 25600
rect 7133 25576 7138 25632
rect 7194 25602 9634 25632
rect 83940 25632 84387 25634
rect 7194 25576 10156 25602
rect 7133 25574 10156 25576
rect 83940 25576 84326 25632
rect 84382 25576 84387 25632
rect 83940 25574 84387 25576
rect 7133 25571 7199 25574
rect 9574 25542 10156 25574
rect 84321 25571 84387 25574
rect 87830 25600 88146 25601
rect 6686 25535 7002 25536
rect 87830 25536 87836 25600
rect 87900 25536 87916 25600
rect 87980 25536 87996 25600
rect 88060 25536 88076 25600
rect 88140 25536 88146 25600
rect 87830 25535 88146 25536
rect 1600 25498 2400 25528
rect 2901 25498 2967 25501
rect 1600 25496 2967 25498
rect 1600 25440 2906 25496
rect 2962 25440 2967 25496
rect 1600 25438 2967 25440
rect 1600 25408 2400 25438
rect 2901 25435 2967 25438
rect 89933 25498 89999 25501
rect 91400 25498 92200 25528
rect 89933 25496 92200 25498
rect 89933 25440 89938 25496
rect 89994 25440 92200 25496
rect 89933 25438 92200 25440
rect 89933 25435 89999 25438
rect 91400 25408 92200 25438
rect 5950 25056 6266 25057
rect 5950 24992 5956 25056
rect 6020 24992 6036 25056
rect 6100 24992 6116 25056
rect 6180 24992 6196 25056
rect 6260 24992 6266 25056
rect 5950 24991 6266 24992
rect 87094 25056 87410 25057
rect 87094 24992 87100 25056
rect 87164 24992 87180 25056
rect 87244 24992 87260 25056
rect 87324 24992 87340 25056
rect 87404 24992 87410 25056
rect 87094 24991 87410 24992
rect 1600 24818 2400 24848
rect 4925 24818 4991 24821
rect 88369 24818 88435 24821
rect 1600 24816 4991 24818
rect 1600 24760 4930 24816
rect 4986 24760 4991 24816
rect 1600 24758 4991 24760
rect 1600 24728 2400 24758
rect 4925 24755 4991 24758
rect 83910 24816 88435 24818
rect 83910 24760 88374 24816
rect 88430 24760 88435 24816
rect 83910 24758 88435 24760
rect 5661 24682 5727 24685
rect 5661 24680 9634 24682
rect 5661 24624 5666 24680
rect 5722 24624 9634 24680
rect 5661 24622 9634 24624
rect 5661 24619 5727 24622
rect 9574 24514 9634 24622
rect 83910 24516 83970 24758
rect 88369 24755 88435 24758
rect 89933 24818 89999 24821
rect 91400 24818 92200 24848
rect 89933 24816 92200 24818
rect 89933 24760 89938 24816
rect 89994 24760 92200 24816
rect 89933 24758 92200 24760
rect 89933 24755 89999 24758
rect 91400 24728 92200 24758
rect 6686 24512 7002 24513
rect 6686 24448 6692 24512
rect 6756 24448 6772 24512
rect 6836 24448 6852 24512
rect 6916 24448 6932 24512
rect 6996 24448 7002 24512
rect 9574 24454 10156 24514
rect 87830 24512 88146 24513
rect 6686 24447 7002 24448
rect 87830 24448 87836 24512
rect 87900 24448 87916 24512
rect 87980 24448 87996 24512
rect 88060 24448 88076 24512
rect 88140 24448 88146 24512
rect 87830 24447 88146 24448
rect 5950 23968 6266 23969
rect 5950 23904 5956 23968
rect 6020 23904 6036 23968
rect 6100 23904 6116 23968
rect 6180 23904 6196 23968
rect 6260 23904 6266 23968
rect 5950 23903 6266 23904
rect 87094 23968 87410 23969
rect 87094 23904 87100 23968
rect 87164 23904 87180 23968
rect 87244 23904 87260 23968
rect 87324 23904 87340 23968
rect 87404 23904 87410 23968
rect 87094 23903 87410 23904
rect 1600 23458 2400 23488
rect 2901 23458 2967 23461
rect 1600 23456 2967 23458
rect 1600 23400 2906 23456
rect 2962 23400 2967 23456
rect 7133 23458 7199 23461
rect 84321 23458 84387 23461
rect 7133 23456 9634 23458
rect 1600 23398 2967 23400
rect 1600 23368 2400 23398
rect 2901 23395 2967 23398
rect 6686 23424 7002 23425
rect 6686 23360 6692 23424
rect 6756 23360 6772 23424
rect 6836 23360 6852 23424
rect 6916 23360 6932 23424
rect 6996 23360 7002 23424
rect 7133 23400 7138 23456
rect 7194 23426 9634 23456
rect 83940 23456 84387 23458
rect 7194 23400 10156 23426
rect 7133 23398 10156 23400
rect 83940 23400 84326 23456
rect 84382 23400 84387 23456
rect 89933 23458 89999 23461
rect 91400 23458 92200 23488
rect 89933 23456 92200 23458
rect 83940 23398 84387 23400
rect 7133 23395 7199 23398
rect 9574 23366 10156 23398
rect 84321 23395 84387 23398
rect 87830 23424 88146 23425
rect 6686 23359 7002 23360
rect 87830 23360 87836 23424
rect 87900 23360 87916 23424
rect 87980 23360 87996 23424
rect 88060 23360 88076 23424
rect 88140 23360 88146 23424
rect 89933 23400 89938 23456
rect 89994 23400 92200 23456
rect 89933 23398 92200 23400
rect 89933 23395 89999 23398
rect 91400 23368 92200 23398
rect 87830 23359 88146 23360
rect 5950 22880 6266 22881
rect 5950 22816 5956 22880
rect 6020 22816 6036 22880
rect 6100 22816 6116 22880
rect 6180 22816 6196 22880
rect 6260 22816 6266 22880
rect 5950 22815 6266 22816
rect 87094 22880 87410 22881
rect 87094 22816 87100 22880
rect 87164 22816 87180 22880
rect 87244 22816 87260 22880
rect 87324 22816 87340 22880
rect 87404 22816 87410 22880
rect 87094 22815 87410 22816
rect 7133 22370 7199 22373
rect 84321 22370 84387 22373
rect 7133 22368 9634 22370
rect 6686 22336 7002 22337
rect 6686 22272 6692 22336
rect 6756 22272 6772 22336
rect 6836 22272 6852 22336
rect 6916 22272 6932 22336
rect 6996 22272 7002 22336
rect 7133 22312 7138 22368
rect 7194 22338 9634 22368
rect 83940 22368 84387 22370
rect 7194 22312 10156 22338
rect 7133 22310 10156 22312
rect 83940 22312 84326 22368
rect 84382 22312 84387 22368
rect 83940 22310 84387 22312
rect 7133 22307 7199 22310
rect 9574 22278 10156 22310
rect 84321 22307 84387 22310
rect 87830 22336 88146 22337
rect 6686 22271 7002 22272
rect 87830 22272 87836 22336
rect 87900 22272 87916 22336
rect 87980 22272 87996 22336
rect 88060 22272 88076 22336
rect 88140 22272 88146 22336
rect 87830 22271 88146 22272
rect 1600 22098 2400 22128
rect 5201 22098 5267 22101
rect 1600 22096 5267 22098
rect 1600 22040 5206 22096
rect 5262 22040 5267 22096
rect 1600 22038 5267 22040
rect 1600 22008 2400 22038
rect 5201 22035 5267 22038
rect 89933 22098 89999 22101
rect 91400 22098 92200 22128
rect 89933 22096 92200 22098
rect 89933 22040 89938 22096
rect 89994 22040 92200 22096
rect 89933 22038 92200 22040
rect 89933 22035 89999 22038
rect 91400 22008 92200 22038
rect 5950 21792 6266 21793
rect 5950 21728 5956 21792
rect 6020 21728 6036 21792
rect 6100 21728 6116 21792
rect 6180 21728 6196 21792
rect 6260 21728 6266 21792
rect 5950 21727 6266 21728
rect 87094 21792 87410 21793
rect 87094 21728 87100 21792
rect 87164 21728 87180 21792
rect 87244 21728 87260 21792
rect 87324 21728 87340 21792
rect 87404 21728 87410 21792
rect 87094 21727 87410 21728
rect 1600 21418 2400 21448
rect 2901 21418 2967 21421
rect 1600 21416 2967 21418
rect 1600 21360 2906 21416
rect 2962 21360 2967 21416
rect 1600 21358 2967 21360
rect 1600 21328 2400 21358
rect 2901 21355 2967 21358
rect 89933 21418 89999 21421
rect 91400 21418 92200 21448
rect 89933 21416 92200 21418
rect 89933 21360 89938 21416
rect 89994 21360 92200 21416
rect 89933 21358 92200 21360
rect 89933 21355 89999 21358
rect 91400 21328 92200 21358
rect 7133 21282 7199 21285
rect 84321 21282 84387 21285
rect 7133 21280 9634 21282
rect 6686 21248 7002 21249
rect 6686 21184 6692 21248
rect 6756 21184 6772 21248
rect 6836 21184 6852 21248
rect 6916 21184 6932 21248
rect 6996 21184 7002 21248
rect 7133 21224 7138 21280
rect 7194 21250 9634 21280
rect 83940 21280 84387 21282
rect 7194 21224 10156 21250
rect 7133 21222 10156 21224
rect 83940 21224 84326 21280
rect 84382 21224 84387 21280
rect 83940 21222 84387 21224
rect 7133 21219 7199 21222
rect 9574 21190 10156 21222
rect 84321 21219 84387 21222
rect 87830 21248 88146 21249
rect 6686 21183 7002 21184
rect 87830 21184 87836 21248
rect 87900 21184 87916 21248
rect 87980 21184 87996 21248
rect 88060 21184 88076 21248
rect 88140 21184 88146 21248
rect 87830 21183 88146 21184
rect 5950 20704 6266 20705
rect 5950 20640 5956 20704
rect 6020 20640 6036 20704
rect 6100 20640 6116 20704
rect 6180 20640 6196 20704
rect 6260 20640 6266 20704
rect 5950 20639 6266 20640
rect 87094 20704 87410 20705
rect 87094 20640 87100 20704
rect 87164 20640 87180 20704
rect 87244 20640 87260 20704
rect 87324 20640 87340 20704
rect 87404 20640 87410 20704
rect 87094 20639 87410 20640
rect 7133 20194 7199 20197
rect 84321 20194 84387 20197
rect 7133 20192 9634 20194
rect 6686 20160 7002 20161
rect 6686 20096 6692 20160
rect 6756 20096 6772 20160
rect 6836 20096 6852 20160
rect 6916 20096 6932 20160
rect 6996 20096 7002 20160
rect 7133 20136 7138 20192
rect 7194 20162 9634 20192
rect 83940 20192 84387 20194
rect 7194 20136 10156 20162
rect 7133 20134 10156 20136
rect 83940 20136 84326 20192
rect 84382 20136 84387 20192
rect 83940 20134 84387 20136
rect 7133 20131 7199 20134
rect 9574 20102 10156 20134
rect 84321 20131 84387 20134
rect 87830 20160 88146 20161
rect 6686 20095 7002 20096
rect 87830 20096 87836 20160
rect 87900 20096 87916 20160
rect 87980 20096 87996 20160
rect 88060 20096 88076 20160
rect 88140 20096 88146 20160
rect 87830 20095 88146 20096
rect 1600 20058 2400 20088
rect 2901 20058 2967 20061
rect 1600 20056 2967 20058
rect 1600 20000 2906 20056
rect 2962 20000 2967 20056
rect 1600 19998 2967 20000
rect 1600 19968 2400 19998
rect 2901 19995 2967 19998
rect 89933 20058 89999 20061
rect 91400 20058 92200 20088
rect 89933 20056 92200 20058
rect 89933 20000 89938 20056
rect 89994 20000 92200 20056
rect 89933 19998 92200 20000
rect 89933 19995 89999 19998
rect 91400 19968 92200 19998
rect 5950 19616 6266 19617
rect 5950 19552 5956 19616
rect 6020 19552 6036 19616
rect 6100 19552 6116 19616
rect 6180 19552 6196 19616
rect 6260 19552 6266 19616
rect 5950 19551 6266 19552
rect 87094 19616 87410 19617
rect 87094 19552 87100 19616
rect 87164 19552 87180 19616
rect 87244 19552 87260 19616
rect 87324 19552 87340 19616
rect 87404 19552 87410 19616
rect 87094 19551 87410 19552
rect 1600 19378 2400 19408
rect 4925 19378 4991 19381
rect 88369 19378 88435 19381
rect 1600 19376 4991 19378
rect 1600 19320 4930 19376
rect 4986 19320 4991 19376
rect 1600 19318 4991 19320
rect 1600 19288 2400 19318
rect 4925 19315 4991 19318
rect 83910 19376 88435 19378
rect 83910 19320 88374 19376
rect 88430 19320 88435 19376
rect 83910 19318 88435 19320
rect 9617 19074 9683 19077
rect 83910 19076 83970 19318
rect 88369 19315 88435 19318
rect 90025 19378 90091 19381
rect 91400 19378 92200 19408
rect 90025 19376 92200 19378
rect 90025 19320 90030 19376
rect 90086 19320 92200 19376
rect 90025 19318 92200 19320
rect 90025 19315 90091 19318
rect 91400 19288 92200 19318
rect 6686 19072 7002 19073
rect 6686 19008 6692 19072
rect 6756 19008 6772 19072
rect 6836 19008 6852 19072
rect 6916 19008 6932 19072
rect 6996 19008 7002 19072
rect 9617 19072 10156 19074
rect 9617 19016 9622 19072
rect 9678 19016 10156 19072
rect 9617 19014 10156 19016
rect 87830 19072 88146 19073
rect 9617 19011 9683 19014
rect 6686 19007 7002 19008
rect 87830 19008 87836 19072
rect 87900 19008 87916 19072
rect 87980 19008 87996 19072
rect 88060 19008 88076 19072
rect 88140 19008 88146 19072
rect 87830 19007 88146 19008
rect 5950 18528 6266 18529
rect 5950 18464 5956 18528
rect 6020 18464 6036 18528
rect 6100 18464 6116 18528
rect 6180 18464 6196 18528
rect 6260 18464 6266 18528
rect 5950 18463 6266 18464
rect 87094 18528 87410 18529
rect 87094 18464 87100 18528
rect 87164 18464 87180 18528
rect 87244 18464 87260 18528
rect 87324 18464 87340 18528
rect 87404 18464 87410 18528
rect 87094 18463 87410 18464
rect 88185 18154 88251 18157
rect 83910 18152 88251 18154
rect 83910 18096 88190 18152
rect 88246 18096 88251 18152
rect 83910 18094 88251 18096
rect 1600 18018 2400 18048
rect 5109 18018 5175 18021
rect 1600 18016 5175 18018
rect 1600 17960 5114 18016
rect 5170 17960 5175 18016
rect 9617 17986 9683 17989
rect 83910 17988 83970 18094
rect 88185 18091 88251 18094
rect 89933 18018 89999 18021
rect 91400 18018 92200 18048
rect 89933 18016 92200 18018
rect 1600 17958 5175 17960
rect 1600 17928 2400 17958
rect 5109 17955 5175 17958
rect 6686 17984 7002 17985
rect 6686 17920 6692 17984
rect 6756 17920 6772 17984
rect 6836 17920 6852 17984
rect 6916 17920 6932 17984
rect 6996 17920 7002 17984
rect 9617 17984 10156 17986
rect 9617 17928 9622 17984
rect 9678 17928 10156 17984
rect 9617 17926 10156 17928
rect 87830 17984 88146 17985
rect 9617 17923 9683 17926
rect 6686 17919 7002 17920
rect 87830 17920 87836 17984
rect 87900 17920 87916 17984
rect 87980 17920 87996 17984
rect 88060 17920 88076 17984
rect 88140 17920 88146 17984
rect 89933 17960 89938 18016
rect 89994 17960 92200 18016
rect 89933 17958 92200 17960
rect 89933 17955 89999 17958
rect 91400 17928 92200 17958
rect 87830 17919 88146 17920
rect 5950 17440 6266 17441
rect 5950 17376 5956 17440
rect 6020 17376 6036 17440
rect 6100 17376 6116 17440
rect 6180 17376 6196 17440
rect 6260 17376 6266 17440
rect 5950 17375 6266 17376
rect 87094 17440 87410 17441
rect 87094 17376 87100 17440
rect 87164 17376 87180 17440
rect 87244 17376 87260 17440
rect 87324 17376 87340 17440
rect 87404 17376 87410 17440
rect 87094 17375 87410 17376
rect 7133 16930 7199 16933
rect 84321 16930 84387 16933
rect 7133 16928 9634 16930
rect 6686 16896 7002 16897
rect 6686 16832 6692 16896
rect 6756 16832 6772 16896
rect 6836 16832 6852 16896
rect 6916 16832 6932 16896
rect 6996 16832 7002 16896
rect 7133 16872 7138 16928
rect 7194 16898 9634 16928
rect 83940 16928 84387 16930
rect 7194 16872 10156 16898
rect 7133 16870 10156 16872
rect 83940 16872 84326 16928
rect 84382 16872 84387 16928
rect 83940 16870 84387 16872
rect 7133 16867 7199 16870
rect 9574 16838 10156 16870
rect 84321 16867 84387 16870
rect 87830 16896 88146 16897
rect 6686 16831 7002 16832
rect 87830 16832 87836 16896
rect 87900 16832 87916 16896
rect 87980 16832 87996 16896
rect 88060 16832 88076 16896
rect 88140 16832 88146 16896
rect 87830 16831 88146 16832
rect 1600 16658 2400 16688
rect 5201 16658 5267 16661
rect 1600 16656 5267 16658
rect 1600 16600 5206 16656
rect 5262 16600 5267 16656
rect 1600 16598 5267 16600
rect 1600 16568 2400 16598
rect 5201 16595 5267 16598
rect 89933 16658 89999 16661
rect 91400 16658 92200 16688
rect 89933 16656 92200 16658
rect 89933 16600 89938 16656
rect 89994 16600 92200 16656
rect 89933 16598 92200 16600
rect 89933 16595 89999 16598
rect 91400 16568 92200 16598
rect 5950 16352 6266 16353
rect 5950 16288 5956 16352
rect 6020 16288 6036 16352
rect 6100 16288 6116 16352
rect 6180 16288 6196 16352
rect 6260 16288 6266 16352
rect 5950 16287 6266 16288
rect 87094 16352 87410 16353
rect 87094 16288 87100 16352
rect 87164 16288 87180 16352
rect 87244 16288 87260 16352
rect 87324 16288 87340 16352
rect 87404 16288 87410 16352
rect 87094 16287 87410 16288
rect 1600 15978 2400 16008
rect 2901 15978 2967 15981
rect 1600 15976 2967 15978
rect 1600 15920 2906 15976
rect 2962 15920 2967 15976
rect 1600 15918 2967 15920
rect 1600 15888 2400 15918
rect 2901 15915 2967 15918
rect 89933 15978 89999 15981
rect 91400 15978 92200 16008
rect 89933 15976 92200 15978
rect 89933 15920 89938 15976
rect 89994 15920 92200 15976
rect 89933 15918 92200 15920
rect 89933 15915 89999 15918
rect 91400 15888 92200 15918
rect 7593 15842 7659 15845
rect 84321 15842 84387 15845
rect 7593 15840 9634 15842
rect 6686 15808 7002 15809
rect 6686 15744 6692 15808
rect 6756 15744 6772 15808
rect 6836 15744 6852 15808
rect 6916 15744 6932 15808
rect 6996 15744 7002 15808
rect 7593 15784 7598 15840
rect 7654 15810 9634 15840
rect 83940 15840 84387 15842
rect 7654 15784 10156 15810
rect 7593 15782 10156 15784
rect 83940 15784 84326 15840
rect 84382 15784 84387 15840
rect 83940 15782 84387 15784
rect 7593 15779 7659 15782
rect 9574 15750 10156 15782
rect 84321 15779 84387 15782
rect 87830 15808 88146 15809
rect 6686 15743 7002 15744
rect 87830 15744 87836 15808
rect 87900 15744 87916 15808
rect 87980 15744 87996 15808
rect 88060 15744 88076 15808
rect 88140 15744 88146 15808
rect 87830 15743 88146 15744
rect 5950 15264 6266 15265
rect 5950 15200 5956 15264
rect 6020 15200 6036 15264
rect 6100 15200 6116 15264
rect 6180 15200 6196 15264
rect 6260 15200 6266 15264
rect 5950 15199 6266 15200
rect 87094 15264 87410 15265
rect 87094 15200 87100 15264
rect 87164 15200 87180 15264
rect 87244 15200 87260 15264
rect 87324 15200 87340 15264
rect 87404 15200 87410 15264
rect 87094 15199 87410 15200
rect 7593 14754 7659 14757
rect 84321 14754 84387 14757
rect 7593 14752 9634 14754
rect 6686 14720 7002 14721
rect 6686 14656 6692 14720
rect 6756 14656 6772 14720
rect 6836 14656 6852 14720
rect 6916 14656 6932 14720
rect 6996 14656 7002 14720
rect 7593 14696 7598 14752
rect 7654 14722 9634 14752
rect 83940 14752 84387 14754
rect 7654 14696 10156 14722
rect 7593 14694 10156 14696
rect 83940 14696 84326 14752
rect 84382 14696 84387 14752
rect 83940 14694 84387 14696
rect 7593 14691 7659 14694
rect 9574 14662 10156 14694
rect 84321 14691 84387 14694
rect 87830 14720 88146 14721
rect 6686 14655 7002 14656
rect 87830 14656 87836 14720
rect 87900 14656 87916 14720
rect 87980 14656 87996 14720
rect 88060 14656 88076 14720
rect 88140 14656 88146 14720
rect 87830 14655 88146 14656
rect 1600 14618 2400 14648
rect 2901 14618 2967 14621
rect 1600 14616 2967 14618
rect 1600 14560 2906 14616
rect 2962 14560 2967 14616
rect 1600 14558 2967 14560
rect 1600 14528 2400 14558
rect 2901 14555 2967 14558
rect 89933 14618 89999 14621
rect 91400 14618 92200 14648
rect 89933 14616 92200 14618
rect 89933 14560 89938 14616
rect 89994 14560 92200 14616
rect 89933 14558 92200 14560
rect 89933 14555 89999 14558
rect 91400 14528 92200 14558
rect 5950 14176 6266 14177
rect 5950 14112 5956 14176
rect 6020 14112 6036 14176
rect 6100 14112 6116 14176
rect 6180 14112 6196 14176
rect 6260 14112 6266 14176
rect 5950 14111 6266 14112
rect 87094 14176 87410 14177
rect 87094 14112 87100 14176
rect 87164 14112 87180 14176
rect 87244 14112 87260 14176
rect 87324 14112 87340 14176
rect 87404 14112 87410 14176
rect 87094 14111 87410 14112
rect 1600 13938 2400 13968
rect 4925 13938 4991 13941
rect 88369 13938 88435 13941
rect 1600 13936 4991 13938
rect 1600 13880 4930 13936
rect 4986 13880 4991 13936
rect 1600 13878 4991 13880
rect 1600 13848 2400 13878
rect 4925 13875 4991 13878
rect 83910 13936 88435 13938
rect 83910 13880 88374 13936
rect 88430 13880 88435 13936
rect 83910 13878 88435 13880
rect 5661 13802 5727 13805
rect 5661 13800 9634 13802
rect 5661 13744 5666 13800
rect 5722 13744 9634 13800
rect 5661 13742 9634 13744
rect 5661 13739 5727 13742
rect 9574 13634 9634 13742
rect 83910 13636 83970 13878
rect 88369 13875 88435 13878
rect 89933 13938 89999 13941
rect 91400 13938 92200 13968
rect 89933 13936 92200 13938
rect 89933 13880 89938 13936
rect 89994 13880 92200 13936
rect 89933 13878 92200 13880
rect 89933 13875 89999 13878
rect 91400 13848 92200 13878
rect 6686 13632 7002 13633
rect 6686 13568 6692 13632
rect 6756 13568 6772 13632
rect 6836 13568 6852 13632
rect 6916 13568 6932 13632
rect 6996 13568 7002 13632
rect 9574 13574 10156 13634
rect 87830 13632 88146 13633
rect 6686 13567 7002 13568
rect 87830 13568 87836 13632
rect 87900 13568 87916 13632
rect 87980 13568 87996 13632
rect 88060 13568 88076 13632
rect 88140 13568 88146 13632
rect 87830 13567 88146 13568
rect 5950 13088 6266 13089
rect 5950 13024 5956 13088
rect 6020 13024 6036 13088
rect 6100 13024 6116 13088
rect 6180 13024 6196 13088
rect 6260 13024 6266 13088
rect 5950 13023 6266 13024
rect 87094 13088 87410 13089
rect 87094 13024 87100 13088
rect 87164 13024 87180 13088
rect 87244 13024 87260 13088
rect 87324 13024 87340 13088
rect 87404 13024 87410 13088
rect 87094 13023 87410 13024
rect 6686 12544 7002 12545
rect 6686 12480 6692 12544
rect 6756 12480 6772 12544
rect 6836 12480 6852 12544
rect 6916 12480 6932 12544
rect 6996 12480 7002 12544
rect 6686 12479 7002 12480
rect 87830 12544 88146 12545
rect 87830 12480 87836 12544
rect 87900 12480 87916 12544
rect 87980 12480 87996 12544
rect 88060 12480 88076 12544
rect 88140 12480 88146 12544
rect 87830 12479 88146 12480
rect 5950 12000 6266 12001
rect 5950 11936 5956 12000
rect 6020 11936 6036 12000
rect 6100 11936 6116 12000
rect 6180 11936 6196 12000
rect 6260 11936 6266 12000
rect 5950 11935 6266 11936
rect 87094 12000 87410 12001
rect 87094 11936 87100 12000
rect 87164 11936 87180 12000
rect 87244 11936 87260 12000
rect 87324 11936 87340 12000
rect 87404 11936 87410 12000
rect 87094 11935 87410 11936
rect 6686 11456 7002 11457
rect 6686 11392 6692 11456
rect 6756 11392 6772 11456
rect 6836 11392 6852 11456
rect 6916 11392 6932 11456
rect 6996 11392 7002 11456
rect 6686 11391 7002 11392
rect 87830 11456 88146 11457
rect 87830 11392 87836 11456
rect 87900 11392 87916 11456
rect 87980 11392 87996 11456
rect 88060 11392 88076 11456
rect 88140 11392 88146 11456
rect 87830 11391 88146 11392
rect 5950 10912 6266 10913
rect 5950 10848 5956 10912
rect 6020 10848 6036 10912
rect 6100 10848 6116 10912
rect 6180 10848 6196 10912
rect 6260 10848 6266 10912
rect 5950 10847 6266 10848
rect 87094 10912 87410 10913
rect 87094 10848 87100 10912
rect 87164 10848 87180 10912
rect 87244 10848 87260 10912
rect 87324 10848 87340 10912
rect 87404 10848 87410 10912
rect 87094 10847 87410 10848
rect 9801 10674 9867 10677
rect 11117 10674 11183 10677
rect 9801 10672 11183 10674
rect 9801 10616 9806 10672
rect 9862 10616 11122 10672
rect 11178 10616 11183 10672
rect 9801 10614 11183 10616
rect 9801 10611 9867 10614
rect 11117 10611 11183 10614
rect 7869 10538 7935 10541
rect 12221 10538 12287 10541
rect 7869 10536 18190 10538
rect 7869 10480 7874 10536
rect 7930 10480 12226 10536
rect 12282 10480 18190 10536
rect 7869 10478 18190 10480
rect 7869 10475 7935 10478
rect 12221 10475 12287 10478
rect 8329 10402 8395 10405
rect 13325 10402 13391 10405
rect 18130 10402 18190 10478
rect 46693 10402 46759 10405
rect 8329 10400 15522 10402
rect 6686 10368 7002 10369
rect 6686 10304 6692 10368
rect 6756 10304 6772 10368
rect 6836 10304 6852 10368
rect 6916 10304 6932 10368
rect 6996 10304 7002 10368
rect 8329 10344 8334 10400
rect 8390 10344 13330 10400
rect 13386 10344 15522 10400
rect 8329 10342 15522 10344
rect 18130 10400 46759 10402
rect 18130 10344 46698 10400
rect 46754 10344 46759 10400
rect 18130 10342 46759 10344
rect 8329 10339 8395 10342
rect 13325 10339 13391 10342
rect 6686 10303 7002 10304
rect 8145 10266 8211 10269
rect 14429 10266 14495 10269
rect 15462 10266 15522 10342
rect 46693 10339 46759 10342
rect 87830 10368 88146 10369
rect 87830 10304 87836 10368
rect 87900 10304 87916 10368
rect 87980 10304 87996 10368
rect 88060 10304 88076 10368
rect 88140 10304 88146 10368
rect 87830 10303 88146 10304
rect 84413 10266 84479 10269
rect 8145 10264 15338 10266
rect 8145 10208 8150 10264
rect 8206 10208 14434 10264
rect 14490 10208 15338 10264
rect 8145 10206 15338 10208
rect 15462 10206 49746 10266
rect 8145 10203 8211 10206
rect 14429 10203 14495 10206
rect 12221 10130 12287 10133
rect 13325 10130 13391 10133
rect 15278 10130 15338 10206
rect 12221 10128 12578 10130
rect 12221 10072 12226 10128
rect 12282 10072 12578 10128
rect 12221 10070 12578 10072
rect 12221 10067 12287 10070
rect 12518 9994 12578 10070
rect 13325 10128 14602 10130
rect 13325 10072 13330 10128
rect 13386 10072 14602 10128
rect 13325 10070 14602 10072
rect 13325 10067 13391 10070
rect 12653 9994 12719 9997
rect 12518 9992 12719 9994
rect 12518 9936 12658 9992
rect 12714 9936 12719 9992
rect 12518 9934 12719 9936
rect 14542 9994 14602 10070
rect 15278 10070 49378 10130
rect 14677 9994 14743 9997
rect 14542 9992 14743 9994
rect 14542 9936 14682 9992
rect 14738 9936 14743 9992
rect 14542 9934 14743 9936
rect 15278 9994 15338 10070
rect 15413 9994 15479 9997
rect 15278 9992 15479 9994
rect 15278 9936 15418 9992
rect 15474 9936 15479 9992
rect 15278 9934 15479 9936
rect 12653 9931 12719 9934
rect 14677 9931 14743 9934
rect 15413 9931 15479 9934
rect 46693 9994 46759 9997
rect 49085 9994 49151 9997
rect 46693 9992 49151 9994
rect 46693 9936 46698 9992
rect 46754 9936 49090 9992
rect 49146 9936 49151 9992
rect 46693 9934 49151 9936
rect 46693 9931 46759 9934
rect 49085 9931 49151 9934
rect 49318 9858 49378 10070
rect 49686 9994 49746 10206
rect 56770 10264 84479 10266
rect 56770 10208 84418 10264
rect 84474 10208 84479 10264
rect 56770 10206 84479 10208
rect 50189 9994 50255 9997
rect 51569 9994 51635 9997
rect 56770 9994 56830 10206
rect 84413 10203 84479 10206
rect 49686 9992 50255 9994
rect 49686 9936 50194 9992
rect 50250 9936 50255 9992
rect 49686 9934 50255 9936
rect 50189 9931 50255 9934
rect 50422 9992 56830 9994
rect 50422 9936 51574 9992
rect 51630 9936 56830 9992
rect 50422 9934 56830 9936
rect 50422 9858 50482 9934
rect 51569 9931 51635 9934
rect 5950 9824 6266 9825
rect 5950 9760 5956 9824
rect 6020 9760 6036 9824
rect 6100 9760 6116 9824
rect 6180 9760 6196 9824
rect 6260 9760 6266 9824
rect 49318 9798 50482 9858
rect 87094 9824 87410 9825
rect 5950 9759 6266 9760
rect 87094 9760 87100 9824
rect 87164 9760 87180 9824
rect 87244 9760 87260 9824
rect 87324 9760 87340 9824
rect 87404 9760 87410 9824
rect 87094 9759 87410 9760
rect 6686 9280 7002 9281
rect 6686 9216 6692 9280
rect 6756 9216 6772 9280
rect 6836 9216 6852 9280
rect 6916 9216 6932 9280
rect 6996 9216 7002 9280
rect 6686 9215 7002 9216
rect 87830 9280 88146 9281
rect 87830 9216 87836 9280
rect 87900 9216 87916 9280
rect 87980 9216 87996 9280
rect 88060 9216 88076 9280
rect 88140 9216 88146 9280
rect 87830 9215 88146 9216
rect 5950 8736 6266 8737
rect 5950 8672 5956 8736
rect 6020 8672 6036 8736
rect 6100 8672 6116 8736
rect 6180 8672 6196 8736
rect 6260 8672 6266 8736
rect 5950 8671 6266 8672
rect 87094 8736 87410 8737
rect 87094 8672 87100 8736
rect 87164 8672 87180 8736
rect 87244 8672 87260 8736
rect 87324 8672 87340 8736
rect 87404 8672 87410 8736
rect 87094 8671 87410 8672
rect 8421 8498 8487 8501
rect 48073 8498 48139 8501
rect 8421 8496 48139 8498
rect 8421 8440 8426 8496
rect 8482 8440 48078 8496
rect 48134 8440 48139 8496
rect 8421 8438 48139 8440
rect 8421 8435 8487 8438
rect 48073 8435 48139 8438
rect 6686 8192 7002 8193
rect 6686 8128 6692 8192
rect 6756 8128 6772 8192
rect 6836 8128 6852 8192
rect 6916 8128 6932 8192
rect 6996 8128 7002 8192
rect 6686 8127 7002 8128
rect 87830 8192 88146 8193
rect 87830 8128 87836 8192
rect 87900 8128 87916 8192
rect 87980 8128 87996 8192
rect 88060 8128 88076 8192
rect 88140 8128 88146 8192
rect 87830 8127 88146 8128
rect 5950 7648 6266 7649
rect 5950 7584 5956 7648
rect 6020 7584 6036 7648
rect 6100 7584 6116 7648
rect 6180 7584 6196 7648
rect 6260 7584 6266 7648
rect 5950 7583 6266 7584
rect 18718 7648 19034 7649
rect 18718 7584 18724 7648
rect 18788 7584 18804 7648
rect 18868 7584 18884 7648
rect 18948 7584 18964 7648
rect 19028 7584 19034 7648
rect 18718 7583 19034 7584
rect 37718 7648 38034 7649
rect 37718 7584 37724 7648
rect 37788 7584 37804 7648
rect 37868 7584 37884 7648
rect 37948 7584 37964 7648
rect 38028 7584 38034 7648
rect 37718 7583 38034 7584
rect 56718 7648 57034 7649
rect 56718 7584 56724 7648
rect 56788 7584 56804 7648
rect 56868 7584 56884 7648
rect 56948 7584 56964 7648
rect 57028 7584 57034 7648
rect 56718 7583 57034 7584
rect 75718 7648 76034 7649
rect 75718 7584 75724 7648
rect 75788 7584 75804 7648
rect 75868 7584 75884 7648
rect 75948 7584 75964 7648
rect 76028 7584 76034 7648
rect 75718 7583 76034 7584
rect 87094 7648 87410 7649
rect 87094 7584 87100 7648
rect 87164 7584 87180 7648
rect 87244 7584 87260 7648
rect 87324 7584 87340 7648
rect 87404 7584 87410 7648
rect 87094 7583 87410 7584
rect 6686 7104 7002 7105
rect 6686 7040 6692 7104
rect 6756 7040 6772 7104
rect 6836 7040 6852 7104
rect 6916 7040 6932 7104
rect 6996 7040 7002 7104
rect 6686 7039 7002 7040
rect 19378 7104 19694 7105
rect 19378 7040 19384 7104
rect 19448 7040 19464 7104
rect 19528 7040 19544 7104
rect 19608 7040 19624 7104
rect 19688 7040 19694 7104
rect 19378 7039 19694 7040
rect 38378 7104 38694 7105
rect 38378 7040 38384 7104
rect 38448 7040 38464 7104
rect 38528 7040 38544 7104
rect 38608 7040 38624 7104
rect 38688 7040 38694 7104
rect 38378 7039 38694 7040
rect 57378 7104 57694 7105
rect 57378 7040 57384 7104
rect 57448 7040 57464 7104
rect 57528 7040 57544 7104
rect 57608 7040 57624 7104
rect 57688 7040 57694 7104
rect 57378 7039 57694 7040
rect 76378 7104 76694 7105
rect 76378 7040 76384 7104
rect 76448 7040 76464 7104
rect 76528 7040 76544 7104
rect 76608 7040 76624 7104
rect 76688 7040 76694 7104
rect 76378 7039 76694 7040
rect 87830 7104 88146 7105
rect 87830 7040 87836 7104
rect 87900 7040 87916 7104
rect 87980 7040 87996 7104
rect 88060 7040 88076 7104
rect 88140 7040 88146 7104
rect 87830 7039 88146 7040
rect 18718 6560 19034 6561
rect 18718 6496 18724 6560
rect 18788 6496 18804 6560
rect 18868 6496 18884 6560
rect 18948 6496 18964 6560
rect 19028 6496 19034 6560
rect 18718 6495 19034 6496
rect 37718 6560 38034 6561
rect 37718 6496 37724 6560
rect 37788 6496 37804 6560
rect 37868 6496 37884 6560
rect 37948 6496 37964 6560
rect 38028 6496 38034 6560
rect 37718 6495 38034 6496
rect 56718 6560 57034 6561
rect 56718 6496 56724 6560
rect 56788 6496 56804 6560
rect 56868 6496 56884 6560
rect 56948 6496 56964 6560
rect 57028 6496 57034 6560
rect 56718 6495 57034 6496
rect 75718 6560 76034 6561
rect 75718 6496 75724 6560
rect 75788 6496 75804 6560
rect 75868 6496 75884 6560
rect 75948 6496 75964 6560
rect 76028 6496 76034 6560
rect 75718 6495 76034 6496
rect 19378 6016 19694 6017
rect 19378 5952 19384 6016
rect 19448 5952 19464 6016
rect 19528 5952 19544 6016
rect 19608 5952 19624 6016
rect 19688 5952 19694 6016
rect 19378 5951 19694 5952
rect 38378 6016 38694 6017
rect 38378 5952 38384 6016
rect 38448 5952 38464 6016
rect 38528 5952 38544 6016
rect 38608 5952 38624 6016
rect 38688 5952 38694 6016
rect 38378 5951 38694 5952
rect 57378 6016 57694 6017
rect 57378 5952 57384 6016
rect 57448 5952 57464 6016
rect 57528 5952 57544 6016
rect 57608 5952 57624 6016
rect 57688 5952 57694 6016
rect 57378 5951 57694 5952
rect 76378 6016 76694 6017
rect 76378 5952 76384 6016
rect 76448 5952 76464 6016
rect 76528 5952 76544 6016
rect 76608 5952 76624 6016
rect 76688 5952 76694 6016
rect 76378 5951 76694 5952
rect 18718 5472 19034 5473
rect 18718 5408 18724 5472
rect 18788 5408 18804 5472
rect 18868 5408 18884 5472
rect 18948 5408 18964 5472
rect 19028 5408 19034 5472
rect 18718 5407 19034 5408
rect 37718 5472 38034 5473
rect 37718 5408 37724 5472
rect 37788 5408 37804 5472
rect 37868 5408 37884 5472
rect 37948 5408 37964 5472
rect 38028 5408 38034 5472
rect 37718 5407 38034 5408
rect 56718 5472 57034 5473
rect 56718 5408 56724 5472
rect 56788 5408 56804 5472
rect 56868 5408 56884 5472
rect 56948 5408 56964 5472
rect 57028 5408 57034 5472
rect 56718 5407 57034 5408
rect 75718 5472 76034 5473
rect 75718 5408 75724 5472
rect 75788 5408 75804 5472
rect 75868 5408 75884 5472
rect 75948 5408 75964 5472
rect 76028 5408 76034 5472
rect 75718 5407 76034 5408
rect 19378 4928 19694 4929
rect 19378 4864 19384 4928
rect 19448 4864 19464 4928
rect 19528 4864 19544 4928
rect 19608 4864 19624 4928
rect 19688 4864 19694 4928
rect 19378 4863 19694 4864
rect 38378 4928 38694 4929
rect 38378 4864 38384 4928
rect 38448 4864 38464 4928
rect 38528 4864 38544 4928
rect 38608 4864 38624 4928
rect 38688 4864 38694 4928
rect 38378 4863 38694 4864
rect 57378 4928 57694 4929
rect 57378 4864 57384 4928
rect 57448 4864 57464 4928
rect 57528 4864 57544 4928
rect 57608 4864 57624 4928
rect 57688 4864 57694 4928
rect 57378 4863 57694 4864
rect 76378 4928 76694 4929
rect 76378 4864 76384 4928
rect 76448 4864 76464 4928
rect 76528 4864 76544 4928
rect 76608 4864 76624 4928
rect 76688 4864 76694 4928
rect 76378 4863 76694 4864
<< via3 >>
rect 18724 89244 18788 89248
rect 18724 89188 18728 89244
rect 18728 89188 18784 89244
rect 18784 89188 18788 89244
rect 18724 89184 18788 89188
rect 18804 89244 18868 89248
rect 18804 89188 18808 89244
rect 18808 89188 18864 89244
rect 18864 89188 18868 89244
rect 18804 89184 18868 89188
rect 18884 89244 18948 89248
rect 18884 89188 18888 89244
rect 18888 89188 18944 89244
rect 18944 89188 18948 89244
rect 18884 89184 18948 89188
rect 18964 89244 19028 89248
rect 18964 89188 18968 89244
rect 18968 89188 19024 89244
rect 19024 89188 19028 89244
rect 18964 89184 19028 89188
rect 37724 89244 37788 89248
rect 37724 89188 37728 89244
rect 37728 89188 37784 89244
rect 37784 89188 37788 89244
rect 37724 89184 37788 89188
rect 37804 89244 37868 89248
rect 37804 89188 37808 89244
rect 37808 89188 37864 89244
rect 37864 89188 37868 89244
rect 37804 89184 37868 89188
rect 37884 89244 37948 89248
rect 37884 89188 37888 89244
rect 37888 89188 37944 89244
rect 37944 89188 37948 89244
rect 37884 89184 37948 89188
rect 37964 89244 38028 89248
rect 37964 89188 37968 89244
rect 37968 89188 38024 89244
rect 38024 89188 38028 89244
rect 37964 89184 38028 89188
rect 56724 89244 56788 89248
rect 56724 89188 56728 89244
rect 56728 89188 56784 89244
rect 56784 89188 56788 89244
rect 56724 89184 56788 89188
rect 56804 89244 56868 89248
rect 56804 89188 56808 89244
rect 56808 89188 56864 89244
rect 56864 89188 56868 89244
rect 56804 89184 56868 89188
rect 56884 89244 56948 89248
rect 56884 89188 56888 89244
rect 56888 89188 56944 89244
rect 56944 89188 56948 89244
rect 56884 89184 56948 89188
rect 56964 89244 57028 89248
rect 56964 89188 56968 89244
rect 56968 89188 57024 89244
rect 57024 89188 57028 89244
rect 56964 89184 57028 89188
rect 75724 89244 75788 89248
rect 75724 89188 75728 89244
rect 75728 89188 75784 89244
rect 75784 89188 75788 89244
rect 75724 89184 75788 89188
rect 75804 89244 75868 89248
rect 75804 89188 75808 89244
rect 75808 89188 75864 89244
rect 75864 89188 75868 89244
rect 75804 89184 75868 89188
rect 75884 89244 75948 89248
rect 75884 89188 75888 89244
rect 75888 89188 75944 89244
rect 75944 89188 75948 89244
rect 75884 89184 75948 89188
rect 75964 89244 76028 89248
rect 75964 89188 75968 89244
rect 75968 89188 76024 89244
rect 76024 89188 76028 89244
rect 75964 89184 76028 89188
rect 19384 88700 19448 88704
rect 19384 88644 19388 88700
rect 19388 88644 19444 88700
rect 19444 88644 19448 88700
rect 19384 88640 19448 88644
rect 19464 88700 19528 88704
rect 19464 88644 19468 88700
rect 19468 88644 19524 88700
rect 19524 88644 19528 88700
rect 19464 88640 19528 88644
rect 19544 88700 19608 88704
rect 19544 88644 19548 88700
rect 19548 88644 19604 88700
rect 19604 88644 19608 88700
rect 19544 88640 19608 88644
rect 19624 88700 19688 88704
rect 19624 88644 19628 88700
rect 19628 88644 19684 88700
rect 19684 88644 19688 88700
rect 19624 88640 19688 88644
rect 38384 88700 38448 88704
rect 38384 88644 38388 88700
rect 38388 88644 38444 88700
rect 38444 88644 38448 88700
rect 38384 88640 38448 88644
rect 38464 88700 38528 88704
rect 38464 88644 38468 88700
rect 38468 88644 38524 88700
rect 38524 88644 38528 88700
rect 38464 88640 38528 88644
rect 38544 88700 38608 88704
rect 38544 88644 38548 88700
rect 38548 88644 38604 88700
rect 38604 88644 38608 88700
rect 38544 88640 38608 88644
rect 38624 88700 38688 88704
rect 38624 88644 38628 88700
rect 38628 88644 38684 88700
rect 38684 88644 38688 88700
rect 38624 88640 38688 88644
rect 57384 88700 57448 88704
rect 57384 88644 57388 88700
rect 57388 88644 57444 88700
rect 57444 88644 57448 88700
rect 57384 88640 57448 88644
rect 57464 88700 57528 88704
rect 57464 88644 57468 88700
rect 57468 88644 57524 88700
rect 57524 88644 57528 88700
rect 57464 88640 57528 88644
rect 57544 88700 57608 88704
rect 57544 88644 57548 88700
rect 57548 88644 57604 88700
rect 57604 88644 57608 88700
rect 57544 88640 57608 88644
rect 57624 88700 57688 88704
rect 57624 88644 57628 88700
rect 57628 88644 57684 88700
rect 57684 88644 57688 88700
rect 57624 88640 57688 88644
rect 76384 88700 76448 88704
rect 76384 88644 76388 88700
rect 76388 88644 76444 88700
rect 76444 88644 76448 88700
rect 76384 88640 76448 88644
rect 76464 88700 76528 88704
rect 76464 88644 76468 88700
rect 76468 88644 76524 88700
rect 76524 88644 76528 88700
rect 76464 88640 76528 88644
rect 76544 88700 76608 88704
rect 76544 88644 76548 88700
rect 76548 88644 76604 88700
rect 76604 88644 76608 88700
rect 76544 88640 76608 88644
rect 76624 88700 76688 88704
rect 76624 88644 76628 88700
rect 76628 88644 76684 88700
rect 76684 88644 76688 88700
rect 76624 88640 76688 88644
rect 18724 88156 18788 88160
rect 18724 88100 18728 88156
rect 18728 88100 18784 88156
rect 18784 88100 18788 88156
rect 18724 88096 18788 88100
rect 18804 88156 18868 88160
rect 18804 88100 18808 88156
rect 18808 88100 18864 88156
rect 18864 88100 18868 88156
rect 18804 88096 18868 88100
rect 18884 88156 18948 88160
rect 18884 88100 18888 88156
rect 18888 88100 18944 88156
rect 18944 88100 18948 88156
rect 18884 88096 18948 88100
rect 18964 88156 19028 88160
rect 18964 88100 18968 88156
rect 18968 88100 19024 88156
rect 19024 88100 19028 88156
rect 18964 88096 19028 88100
rect 37724 88156 37788 88160
rect 37724 88100 37728 88156
rect 37728 88100 37784 88156
rect 37784 88100 37788 88156
rect 37724 88096 37788 88100
rect 37804 88156 37868 88160
rect 37804 88100 37808 88156
rect 37808 88100 37864 88156
rect 37864 88100 37868 88156
rect 37804 88096 37868 88100
rect 37884 88156 37948 88160
rect 37884 88100 37888 88156
rect 37888 88100 37944 88156
rect 37944 88100 37948 88156
rect 37884 88096 37948 88100
rect 37964 88156 38028 88160
rect 37964 88100 37968 88156
rect 37968 88100 38024 88156
rect 38024 88100 38028 88156
rect 37964 88096 38028 88100
rect 56724 88156 56788 88160
rect 56724 88100 56728 88156
rect 56728 88100 56784 88156
rect 56784 88100 56788 88156
rect 56724 88096 56788 88100
rect 56804 88156 56868 88160
rect 56804 88100 56808 88156
rect 56808 88100 56864 88156
rect 56864 88100 56868 88156
rect 56804 88096 56868 88100
rect 56884 88156 56948 88160
rect 56884 88100 56888 88156
rect 56888 88100 56944 88156
rect 56944 88100 56948 88156
rect 56884 88096 56948 88100
rect 56964 88156 57028 88160
rect 56964 88100 56968 88156
rect 56968 88100 57024 88156
rect 57024 88100 57028 88156
rect 56964 88096 57028 88100
rect 75724 88156 75788 88160
rect 75724 88100 75728 88156
rect 75728 88100 75784 88156
rect 75784 88100 75788 88156
rect 75724 88096 75788 88100
rect 75804 88156 75868 88160
rect 75804 88100 75808 88156
rect 75808 88100 75864 88156
rect 75864 88100 75868 88156
rect 75804 88096 75868 88100
rect 75884 88156 75948 88160
rect 75884 88100 75888 88156
rect 75888 88100 75944 88156
rect 75944 88100 75948 88156
rect 75884 88096 75948 88100
rect 75964 88156 76028 88160
rect 75964 88100 75968 88156
rect 75968 88100 76024 88156
rect 76024 88100 76028 88156
rect 75964 88096 76028 88100
rect 19384 87612 19448 87616
rect 19384 87556 19388 87612
rect 19388 87556 19444 87612
rect 19444 87556 19448 87612
rect 19384 87552 19448 87556
rect 19464 87612 19528 87616
rect 19464 87556 19468 87612
rect 19468 87556 19524 87612
rect 19524 87556 19528 87612
rect 19464 87552 19528 87556
rect 19544 87612 19608 87616
rect 19544 87556 19548 87612
rect 19548 87556 19604 87612
rect 19604 87556 19608 87612
rect 19544 87552 19608 87556
rect 19624 87612 19688 87616
rect 19624 87556 19628 87612
rect 19628 87556 19684 87612
rect 19684 87556 19688 87612
rect 19624 87552 19688 87556
rect 38384 87612 38448 87616
rect 38384 87556 38388 87612
rect 38388 87556 38444 87612
rect 38444 87556 38448 87612
rect 38384 87552 38448 87556
rect 38464 87612 38528 87616
rect 38464 87556 38468 87612
rect 38468 87556 38524 87612
rect 38524 87556 38528 87612
rect 38464 87552 38528 87556
rect 38544 87612 38608 87616
rect 38544 87556 38548 87612
rect 38548 87556 38604 87612
rect 38604 87556 38608 87612
rect 38544 87552 38608 87556
rect 38624 87612 38688 87616
rect 38624 87556 38628 87612
rect 38628 87556 38684 87612
rect 38684 87556 38688 87612
rect 38624 87552 38688 87556
rect 57384 87612 57448 87616
rect 57384 87556 57388 87612
rect 57388 87556 57444 87612
rect 57444 87556 57448 87612
rect 57384 87552 57448 87556
rect 57464 87612 57528 87616
rect 57464 87556 57468 87612
rect 57468 87556 57524 87612
rect 57524 87556 57528 87612
rect 57464 87552 57528 87556
rect 57544 87612 57608 87616
rect 57544 87556 57548 87612
rect 57548 87556 57604 87612
rect 57604 87556 57608 87612
rect 57544 87552 57608 87556
rect 57624 87612 57688 87616
rect 57624 87556 57628 87612
rect 57628 87556 57684 87612
rect 57684 87556 57688 87612
rect 57624 87552 57688 87556
rect 76384 87612 76448 87616
rect 76384 87556 76388 87612
rect 76388 87556 76444 87612
rect 76444 87556 76448 87612
rect 76384 87552 76448 87556
rect 76464 87612 76528 87616
rect 76464 87556 76468 87612
rect 76468 87556 76524 87612
rect 76524 87556 76528 87612
rect 76464 87552 76528 87556
rect 76544 87612 76608 87616
rect 76544 87556 76548 87612
rect 76548 87556 76604 87612
rect 76604 87556 76608 87612
rect 76544 87552 76608 87556
rect 76624 87612 76688 87616
rect 76624 87556 76628 87612
rect 76628 87556 76684 87612
rect 76684 87556 76688 87612
rect 76624 87552 76688 87556
rect 5956 87068 6020 87072
rect 5956 87012 5960 87068
rect 5960 87012 6016 87068
rect 6016 87012 6020 87068
rect 5956 87008 6020 87012
rect 6036 87068 6100 87072
rect 6036 87012 6040 87068
rect 6040 87012 6096 87068
rect 6096 87012 6100 87068
rect 6036 87008 6100 87012
rect 6116 87068 6180 87072
rect 6116 87012 6120 87068
rect 6120 87012 6176 87068
rect 6176 87012 6180 87068
rect 6116 87008 6180 87012
rect 6196 87068 6260 87072
rect 6196 87012 6200 87068
rect 6200 87012 6256 87068
rect 6256 87012 6260 87068
rect 6196 87008 6260 87012
rect 18724 87068 18788 87072
rect 18724 87012 18728 87068
rect 18728 87012 18784 87068
rect 18784 87012 18788 87068
rect 18724 87008 18788 87012
rect 18804 87068 18868 87072
rect 18804 87012 18808 87068
rect 18808 87012 18864 87068
rect 18864 87012 18868 87068
rect 18804 87008 18868 87012
rect 18884 87068 18948 87072
rect 18884 87012 18888 87068
rect 18888 87012 18944 87068
rect 18944 87012 18948 87068
rect 18884 87008 18948 87012
rect 18964 87068 19028 87072
rect 18964 87012 18968 87068
rect 18968 87012 19024 87068
rect 19024 87012 19028 87068
rect 18964 87008 19028 87012
rect 37724 87068 37788 87072
rect 37724 87012 37728 87068
rect 37728 87012 37784 87068
rect 37784 87012 37788 87068
rect 37724 87008 37788 87012
rect 37804 87068 37868 87072
rect 37804 87012 37808 87068
rect 37808 87012 37864 87068
rect 37864 87012 37868 87068
rect 37804 87008 37868 87012
rect 37884 87068 37948 87072
rect 37884 87012 37888 87068
rect 37888 87012 37944 87068
rect 37944 87012 37948 87068
rect 37884 87008 37948 87012
rect 37964 87068 38028 87072
rect 37964 87012 37968 87068
rect 37968 87012 38024 87068
rect 38024 87012 38028 87068
rect 37964 87008 38028 87012
rect 56724 87068 56788 87072
rect 56724 87012 56728 87068
rect 56728 87012 56784 87068
rect 56784 87012 56788 87068
rect 56724 87008 56788 87012
rect 56804 87068 56868 87072
rect 56804 87012 56808 87068
rect 56808 87012 56864 87068
rect 56864 87012 56868 87068
rect 56804 87008 56868 87012
rect 56884 87068 56948 87072
rect 56884 87012 56888 87068
rect 56888 87012 56944 87068
rect 56944 87012 56948 87068
rect 56884 87008 56948 87012
rect 56964 87068 57028 87072
rect 56964 87012 56968 87068
rect 56968 87012 57024 87068
rect 57024 87012 57028 87068
rect 56964 87008 57028 87012
rect 75724 87068 75788 87072
rect 75724 87012 75728 87068
rect 75728 87012 75784 87068
rect 75784 87012 75788 87068
rect 75724 87008 75788 87012
rect 75804 87068 75868 87072
rect 75804 87012 75808 87068
rect 75808 87012 75864 87068
rect 75864 87012 75868 87068
rect 75804 87008 75868 87012
rect 75884 87068 75948 87072
rect 75884 87012 75888 87068
rect 75888 87012 75944 87068
rect 75944 87012 75948 87068
rect 75884 87008 75948 87012
rect 75964 87068 76028 87072
rect 75964 87012 75968 87068
rect 75968 87012 76024 87068
rect 76024 87012 76028 87068
rect 75964 87008 76028 87012
rect 87100 87068 87164 87072
rect 87100 87012 87104 87068
rect 87104 87012 87160 87068
rect 87160 87012 87164 87068
rect 87100 87008 87164 87012
rect 87180 87068 87244 87072
rect 87180 87012 87184 87068
rect 87184 87012 87240 87068
rect 87240 87012 87244 87068
rect 87180 87008 87244 87012
rect 87260 87068 87324 87072
rect 87260 87012 87264 87068
rect 87264 87012 87320 87068
rect 87320 87012 87324 87068
rect 87260 87008 87324 87012
rect 87340 87068 87404 87072
rect 87340 87012 87344 87068
rect 87344 87012 87400 87068
rect 87400 87012 87404 87068
rect 87340 87008 87404 87012
rect 6692 86524 6756 86528
rect 6692 86468 6696 86524
rect 6696 86468 6752 86524
rect 6752 86468 6756 86524
rect 6692 86464 6756 86468
rect 6772 86524 6836 86528
rect 6772 86468 6776 86524
rect 6776 86468 6832 86524
rect 6832 86468 6836 86524
rect 6772 86464 6836 86468
rect 6852 86524 6916 86528
rect 6852 86468 6856 86524
rect 6856 86468 6912 86524
rect 6912 86468 6916 86524
rect 6852 86464 6916 86468
rect 6932 86524 6996 86528
rect 6932 86468 6936 86524
rect 6936 86468 6992 86524
rect 6992 86468 6996 86524
rect 6932 86464 6996 86468
rect 19384 86524 19448 86528
rect 19384 86468 19388 86524
rect 19388 86468 19444 86524
rect 19444 86468 19448 86524
rect 19384 86464 19448 86468
rect 19464 86524 19528 86528
rect 19464 86468 19468 86524
rect 19468 86468 19524 86524
rect 19524 86468 19528 86524
rect 19464 86464 19528 86468
rect 19544 86524 19608 86528
rect 19544 86468 19548 86524
rect 19548 86468 19604 86524
rect 19604 86468 19608 86524
rect 19544 86464 19608 86468
rect 19624 86524 19688 86528
rect 19624 86468 19628 86524
rect 19628 86468 19684 86524
rect 19684 86468 19688 86524
rect 19624 86464 19688 86468
rect 38384 86524 38448 86528
rect 38384 86468 38388 86524
rect 38388 86468 38444 86524
rect 38444 86468 38448 86524
rect 38384 86464 38448 86468
rect 38464 86524 38528 86528
rect 38464 86468 38468 86524
rect 38468 86468 38524 86524
rect 38524 86468 38528 86524
rect 38464 86464 38528 86468
rect 38544 86524 38608 86528
rect 38544 86468 38548 86524
rect 38548 86468 38604 86524
rect 38604 86468 38608 86524
rect 38544 86464 38608 86468
rect 38624 86524 38688 86528
rect 38624 86468 38628 86524
rect 38628 86468 38684 86524
rect 38684 86468 38688 86524
rect 38624 86464 38688 86468
rect 57384 86524 57448 86528
rect 57384 86468 57388 86524
rect 57388 86468 57444 86524
rect 57444 86468 57448 86524
rect 57384 86464 57448 86468
rect 57464 86524 57528 86528
rect 57464 86468 57468 86524
rect 57468 86468 57524 86524
rect 57524 86468 57528 86524
rect 57464 86464 57528 86468
rect 57544 86524 57608 86528
rect 57544 86468 57548 86524
rect 57548 86468 57604 86524
rect 57604 86468 57608 86524
rect 57544 86464 57608 86468
rect 57624 86524 57688 86528
rect 57624 86468 57628 86524
rect 57628 86468 57684 86524
rect 57684 86468 57688 86524
rect 57624 86464 57688 86468
rect 76384 86524 76448 86528
rect 76384 86468 76388 86524
rect 76388 86468 76444 86524
rect 76444 86468 76448 86524
rect 76384 86464 76448 86468
rect 76464 86524 76528 86528
rect 76464 86468 76468 86524
rect 76468 86468 76524 86524
rect 76524 86468 76528 86524
rect 76464 86464 76528 86468
rect 76544 86524 76608 86528
rect 76544 86468 76548 86524
rect 76548 86468 76604 86524
rect 76604 86468 76608 86524
rect 76544 86464 76608 86468
rect 76624 86524 76688 86528
rect 76624 86468 76628 86524
rect 76628 86468 76684 86524
rect 76684 86468 76688 86524
rect 76624 86464 76688 86468
rect 87836 86524 87900 86528
rect 87836 86468 87840 86524
rect 87840 86468 87896 86524
rect 87896 86468 87900 86524
rect 87836 86464 87900 86468
rect 87916 86524 87980 86528
rect 87916 86468 87920 86524
rect 87920 86468 87976 86524
rect 87976 86468 87980 86524
rect 87916 86464 87980 86468
rect 87996 86524 88060 86528
rect 87996 86468 88000 86524
rect 88000 86468 88056 86524
rect 88056 86468 88060 86524
rect 87996 86464 88060 86468
rect 88076 86524 88140 86528
rect 88076 86468 88080 86524
rect 88080 86468 88136 86524
rect 88136 86468 88140 86524
rect 88076 86464 88140 86468
rect 5956 85980 6020 85984
rect 5956 85924 5960 85980
rect 5960 85924 6016 85980
rect 6016 85924 6020 85980
rect 5956 85920 6020 85924
rect 6036 85980 6100 85984
rect 6036 85924 6040 85980
rect 6040 85924 6096 85980
rect 6096 85924 6100 85980
rect 6036 85920 6100 85924
rect 6116 85980 6180 85984
rect 6116 85924 6120 85980
rect 6120 85924 6176 85980
rect 6176 85924 6180 85980
rect 6116 85920 6180 85924
rect 6196 85980 6260 85984
rect 6196 85924 6200 85980
rect 6200 85924 6256 85980
rect 6256 85924 6260 85980
rect 6196 85920 6260 85924
rect 87100 85980 87164 85984
rect 87100 85924 87104 85980
rect 87104 85924 87160 85980
rect 87160 85924 87164 85980
rect 87100 85920 87164 85924
rect 87180 85980 87244 85984
rect 87180 85924 87184 85980
rect 87184 85924 87240 85980
rect 87240 85924 87244 85980
rect 87180 85920 87244 85924
rect 87260 85980 87324 85984
rect 87260 85924 87264 85980
rect 87264 85924 87320 85980
rect 87320 85924 87324 85980
rect 87260 85920 87324 85924
rect 87340 85980 87404 85984
rect 87340 85924 87344 85980
rect 87344 85924 87400 85980
rect 87400 85924 87404 85980
rect 87340 85920 87404 85924
rect 6692 85436 6756 85440
rect 6692 85380 6696 85436
rect 6696 85380 6752 85436
rect 6752 85380 6756 85436
rect 6692 85376 6756 85380
rect 6772 85436 6836 85440
rect 6772 85380 6776 85436
rect 6776 85380 6832 85436
rect 6832 85380 6836 85436
rect 6772 85376 6836 85380
rect 6852 85436 6916 85440
rect 6852 85380 6856 85436
rect 6856 85380 6912 85436
rect 6912 85380 6916 85436
rect 6852 85376 6916 85380
rect 6932 85436 6996 85440
rect 6932 85380 6936 85436
rect 6936 85380 6992 85436
rect 6992 85380 6996 85436
rect 6932 85376 6996 85380
rect 87836 85436 87900 85440
rect 87836 85380 87840 85436
rect 87840 85380 87896 85436
rect 87896 85380 87900 85436
rect 87836 85376 87900 85380
rect 87916 85436 87980 85440
rect 87916 85380 87920 85436
rect 87920 85380 87976 85436
rect 87976 85380 87980 85436
rect 87916 85376 87980 85380
rect 87996 85436 88060 85440
rect 87996 85380 88000 85436
rect 88000 85380 88056 85436
rect 88056 85380 88060 85436
rect 87996 85376 88060 85380
rect 88076 85436 88140 85440
rect 88076 85380 88080 85436
rect 88080 85380 88136 85436
rect 88136 85380 88140 85436
rect 88076 85376 88140 85380
rect 5956 84892 6020 84896
rect 5956 84836 5960 84892
rect 5960 84836 6016 84892
rect 6016 84836 6020 84892
rect 5956 84832 6020 84836
rect 6036 84892 6100 84896
rect 6036 84836 6040 84892
rect 6040 84836 6096 84892
rect 6096 84836 6100 84892
rect 6036 84832 6100 84836
rect 6116 84892 6180 84896
rect 6116 84836 6120 84892
rect 6120 84836 6176 84892
rect 6176 84836 6180 84892
rect 6116 84832 6180 84836
rect 6196 84892 6260 84896
rect 6196 84836 6200 84892
rect 6200 84836 6256 84892
rect 6256 84836 6260 84892
rect 6196 84832 6260 84836
rect 87100 84892 87164 84896
rect 87100 84836 87104 84892
rect 87104 84836 87160 84892
rect 87160 84836 87164 84892
rect 87100 84832 87164 84836
rect 87180 84892 87244 84896
rect 87180 84836 87184 84892
rect 87184 84836 87240 84892
rect 87240 84836 87244 84892
rect 87180 84832 87244 84836
rect 87260 84892 87324 84896
rect 87260 84836 87264 84892
rect 87264 84836 87320 84892
rect 87320 84836 87324 84892
rect 87260 84832 87324 84836
rect 87340 84892 87404 84896
rect 87340 84836 87344 84892
rect 87344 84836 87400 84892
rect 87400 84836 87404 84892
rect 87340 84832 87404 84836
rect 6692 84348 6756 84352
rect 6692 84292 6696 84348
rect 6696 84292 6752 84348
rect 6752 84292 6756 84348
rect 6692 84288 6756 84292
rect 6772 84348 6836 84352
rect 6772 84292 6776 84348
rect 6776 84292 6832 84348
rect 6832 84292 6836 84348
rect 6772 84288 6836 84292
rect 6852 84348 6916 84352
rect 6852 84292 6856 84348
rect 6856 84292 6912 84348
rect 6912 84292 6916 84348
rect 6852 84288 6916 84292
rect 6932 84348 6996 84352
rect 6932 84292 6936 84348
rect 6936 84292 6992 84348
rect 6992 84292 6996 84348
rect 6932 84288 6996 84292
rect 87836 84348 87900 84352
rect 87836 84292 87840 84348
rect 87840 84292 87896 84348
rect 87896 84292 87900 84348
rect 87836 84288 87900 84292
rect 87916 84348 87980 84352
rect 87916 84292 87920 84348
rect 87920 84292 87976 84348
rect 87976 84292 87980 84348
rect 87916 84288 87980 84292
rect 87996 84348 88060 84352
rect 87996 84292 88000 84348
rect 88000 84292 88056 84348
rect 88056 84292 88060 84348
rect 87996 84288 88060 84292
rect 88076 84348 88140 84352
rect 88076 84292 88080 84348
rect 88080 84292 88136 84348
rect 88136 84292 88140 84348
rect 88076 84288 88140 84292
rect 5956 83804 6020 83808
rect 5956 83748 5960 83804
rect 5960 83748 6016 83804
rect 6016 83748 6020 83804
rect 5956 83744 6020 83748
rect 6036 83804 6100 83808
rect 6036 83748 6040 83804
rect 6040 83748 6096 83804
rect 6096 83748 6100 83804
rect 6036 83744 6100 83748
rect 6116 83804 6180 83808
rect 6116 83748 6120 83804
rect 6120 83748 6176 83804
rect 6176 83748 6180 83804
rect 6116 83744 6180 83748
rect 6196 83804 6260 83808
rect 6196 83748 6200 83804
rect 6200 83748 6256 83804
rect 6256 83748 6260 83804
rect 6196 83744 6260 83748
rect 87100 83804 87164 83808
rect 87100 83748 87104 83804
rect 87104 83748 87160 83804
rect 87160 83748 87164 83804
rect 87100 83744 87164 83748
rect 87180 83804 87244 83808
rect 87180 83748 87184 83804
rect 87184 83748 87240 83804
rect 87240 83748 87244 83804
rect 87180 83744 87244 83748
rect 87260 83804 87324 83808
rect 87260 83748 87264 83804
rect 87264 83748 87320 83804
rect 87320 83748 87324 83804
rect 87260 83744 87324 83748
rect 87340 83804 87404 83808
rect 87340 83748 87344 83804
rect 87344 83748 87400 83804
rect 87400 83748 87404 83804
rect 87340 83744 87404 83748
rect 6692 83260 6756 83264
rect 6692 83204 6696 83260
rect 6696 83204 6752 83260
rect 6752 83204 6756 83260
rect 6692 83200 6756 83204
rect 6772 83260 6836 83264
rect 6772 83204 6776 83260
rect 6776 83204 6832 83260
rect 6832 83204 6836 83260
rect 6772 83200 6836 83204
rect 6852 83260 6916 83264
rect 6852 83204 6856 83260
rect 6856 83204 6912 83260
rect 6912 83204 6916 83260
rect 6852 83200 6916 83204
rect 6932 83260 6996 83264
rect 6932 83204 6936 83260
rect 6936 83204 6992 83260
rect 6992 83204 6996 83260
rect 6932 83200 6996 83204
rect 87836 83260 87900 83264
rect 87836 83204 87840 83260
rect 87840 83204 87896 83260
rect 87896 83204 87900 83260
rect 87836 83200 87900 83204
rect 87916 83260 87980 83264
rect 87916 83204 87920 83260
rect 87920 83204 87976 83260
rect 87976 83204 87980 83260
rect 87916 83200 87980 83204
rect 87996 83260 88060 83264
rect 87996 83204 88000 83260
rect 88000 83204 88056 83260
rect 88056 83204 88060 83260
rect 87996 83200 88060 83204
rect 88076 83260 88140 83264
rect 88076 83204 88080 83260
rect 88080 83204 88136 83260
rect 88136 83204 88140 83260
rect 88076 83200 88140 83204
rect 5956 82716 6020 82720
rect 5956 82660 5960 82716
rect 5960 82660 6016 82716
rect 6016 82660 6020 82716
rect 5956 82656 6020 82660
rect 6036 82716 6100 82720
rect 6036 82660 6040 82716
rect 6040 82660 6096 82716
rect 6096 82660 6100 82716
rect 6036 82656 6100 82660
rect 6116 82716 6180 82720
rect 6116 82660 6120 82716
rect 6120 82660 6176 82716
rect 6176 82660 6180 82716
rect 6116 82656 6180 82660
rect 6196 82716 6260 82720
rect 6196 82660 6200 82716
rect 6200 82660 6256 82716
rect 6256 82660 6260 82716
rect 6196 82656 6260 82660
rect 87100 82716 87164 82720
rect 87100 82660 87104 82716
rect 87104 82660 87160 82716
rect 87160 82660 87164 82716
rect 87100 82656 87164 82660
rect 87180 82716 87244 82720
rect 87180 82660 87184 82716
rect 87184 82660 87240 82716
rect 87240 82660 87244 82716
rect 87180 82656 87244 82660
rect 87260 82716 87324 82720
rect 87260 82660 87264 82716
rect 87264 82660 87320 82716
rect 87320 82660 87324 82716
rect 87260 82656 87324 82660
rect 87340 82716 87404 82720
rect 87340 82660 87344 82716
rect 87344 82660 87400 82716
rect 87400 82660 87404 82716
rect 87340 82656 87404 82660
rect 6692 82172 6756 82176
rect 6692 82116 6696 82172
rect 6696 82116 6752 82172
rect 6752 82116 6756 82172
rect 6692 82112 6756 82116
rect 6772 82172 6836 82176
rect 6772 82116 6776 82172
rect 6776 82116 6832 82172
rect 6832 82116 6836 82172
rect 6772 82112 6836 82116
rect 6852 82172 6916 82176
rect 6852 82116 6856 82172
rect 6856 82116 6912 82172
rect 6912 82116 6916 82172
rect 6852 82112 6916 82116
rect 6932 82172 6996 82176
rect 6932 82116 6936 82172
rect 6936 82116 6992 82172
rect 6992 82116 6996 82172
rect 6932 82112 6996 82116
rect 87836 82172 87900 82176
rect 87836 82116 87840 82172
rect 87840 82116 87896 82172
rect 87896 82116 87900 82172
rect 87836 82112 87900 82116
rect 87916 82172 87980 82176
rect 87916 82116 87920 82172
rect 87920 82116 87976 82172
rect 87976 82116 87980 82172
rect 87916 82112 87980 82116
rect 87996 82172 88060 82176
rect 87996 82116 88000 82172
rect 88000 82116 88056 82172
rect 88056 82116 88060 82172
rect 87996 82112 88060 82116
rect 88076 82172 88140 82176
rect 88076 82116 88080 82172
rect 88080 82116 88136 82172
rect 88136 82116 88140 82172
rect 88076 82112 88140 82116
rect 5956 81628 6020 81632
rect 5956 81572 5960 81628
rect 5960 81572 6016 81628
rect 6016 81572 6020 81628
rect 5956 81568 6020 81572
rect 6036 81628 6100 81632
rect 6036 81572 6040 81628
rect 6040 81572 6096 81628
rect 6096 81572 6100 81628
rect 6036 81568 6100 81572
rect 6116 81628 6180 81632
rect 6116 81572 6120 81628
rect 6120 81572 6176 81628
rect 6176 81572 6180 81628
rect 6116 81568 6180 81572
rect 6196 81628 6260 81632
rect 6196 81572 6200 81628
rect 6200 81572 6256 81628
rect 6256 81572 6260 81628
rect 6196 81568 6260 81572
rect 87100 81628 87164 81632
rect 87100 81572 87104 81628
rect 87104 81572 87160 81628
rect 87160 81572 87164 81628
rect 87100 81568 87164 81572
rect 87180 81628 87244 81632
rect 87180 81572 87184 81628
rect 87184 81572 87240 81628
rect 87240 81572 87244 81628
rect 87180 81568 87244 81572
rect 87260 81628 87324 81632
rect 87260 81572 87264 81628
rect 87264 81572 87320 81628
rect 87320 81572 87324 81628
rect 87260 81568 87324 81572
rect 87340 81628 87404 81632
rect 87340 81572 87344 81628
rect 87344 81572 87400 81628
rect 87400 81572 87404 81628
rect 87340 81568 87404 81572
rect 6692 81084 6756 81088
rect 6692 81028 6696 81084
rect 6696 81028 6752 81084
rect 6752 81028 6756 81084
rect 6692 81024 6756 81028
rect 6772 81084 6836 81088
rect 6772 81028 6776 81084
rect 6776 81028 6832 81084
rect 6832 81028 6836 81084
rect 6772 81024 6836 81028
rect 6852 81084 6916 81088
rect 6852 81028 6856 81084
rect 6856 81028 6912 81084
rect 6912 81028 6916 81084
rect 6852 81024 6916 81028
rect 6932 81084 6996 81088
rect 6932 81028 6936 81084
rect 6936 81028 6992 81084
rect 6992 81028 6996 81084
rect 6932 81024 6996 81028
rect 87836 81084 87900 81088
rect 87836 81028 87840 81084
rect 87840 81028 87896 81084
rect 87896 81028 87900 81084
rect 87836 81024 87900 81028
rect 87916 81084 87980 81088
rect 87916 81028 87920 81084
rect 87920 81028 87976 81084
rect 87976 81028 87980 81084
rect 87916 81024 87980 81028
rect 87996 81084 88060 81088
rect 87996 81028 88000 81084
rect 88000 81028 88056 81084
rect 88056 81028 88060 81084
rect 87996 81024 88060 81028
rect 88076 81084 88140 81088
rect 88076 81028 88080 81084
rect 88080 81028 88136 81084
rect 88136 81028 88140 81084
rect 88076 81024 88140 81028
rect 5956 80540 6020 80544
rect 5956 80484 5960 80540
rect 5960 80484 6016 80540
rect 6016 80484 6020 80540
rect 5956 80480 6020 80484
rect 6036 80540 6100 80544
rect 6036 80484 6040 80540
rect 6040 80484 6096 80540
rect 6096 80484 6100 80540
rect 6036 80480 6100 80484
rect 6116 80540 6180 80544
rect 6116 80484 6120 80540
rect 6120 80484 6176 80540
rect 6176 80484 6180 80540
rect 6116 80480 6180 80484
rect 6196 80540 6260 80544
rect 6196 80484 6200 80540
rect 6200 80484 6256 80540
rect 6256 80484 6260 80540
rect 6196 80480 6260 80484
rect 87100 80540 87164 80544
rect 87100 80484 87104 80540
rect 87104 80484 87160 80540
rect 87160 80484 87164 80540
rect 87100 80480 87164 80484
rect 87180 80540 87244 80544
rect 87180 80484 87184 80540
rect 87184 80484 87240 80540
rect 87240 80484 87244 80540
rect 87180 80480 87244 80484
rect 87260 80540 87324 80544
rect 87260 80484 87264 80540
rect 87264 80484 87320 80540
rect 87320 80484 87324 80540
rect 87260 80480 87324 80484
rect 87340 80540 87404 80544
rect 87340 80484 87344 80540
rect 87344 80484 87400 80540
rect 87400 80484 87404 80540
rect 87340 80480 87404 80484
rect 6692 79996 6756 80000
rect 6692 79940 6696 79996
rect 6696 79940 6752 79996
rect 6752 79940 6756 79996
rect 6692 79936 6756 79940
rect 6772 79996 6836 80000
rect 6772 79940 6776 79996
rect 6776 79940 6832 79996
rect 6832 79940 6836 79996
rect 6772 79936 6836 79940
rect 6852 79996 6916 80000
rect 6852 79940 6856 79996
rect 6856 79940 6912 79996
rect 6912 79940 6916 79996
rect 6852 79936 6916 79940
rect 6932 79996 6996 80000
rect 6932 79940 6936 79996
rect 6936 79940 6992 79996
rect 6992 79940 6996 79996
rect 6932 79936 6996 79940
rect 87836 79996 87900 80000
rect 87836 79940 87840 79996
rect 87840 79940 87896 79996
rect 87896 79940 87900 79996
rect 87836 79936 87900 79940
rect 87916 79996 87980 80000
rect 87916 79940 87920 79996
rect 87920 79940 87976 79996
rect 87976 79940 87980 79996
rect 87916 79936 87980 79940
rect 87996 79996 88060 80000
rect 87996 79940 88000 79996
rect 88000 79940 88056 79996
rect 88056 79940 88060 79996
rect 87996 79936 88060 79940
rect 88076 79996 88140 80000
rect 88076 79940 88080 79996
rect 88080 79940 88136 79996
rect 88136 79940 88140 79996
rect 88076 79936 88140 79940
rect 5956 79452 6020 79456
rect 5956 79396 5960 79452
rect 5960 79396 6016 79452
rect 6016 79396 6020 79452
rect 5956 79392 6020 79396
rect 6036 79452 6100 79456
rect 6036 79396 6040 79452
rect 6040 79396 6096 79452
rect 6096 79396 6100 79452
rect 6036 79392 6100 79396
rect 6116 79452 6180 79456
rect 6116 79396 6120 79452
rect 6120 79396 6176 79452
rect 6176 79396 6180 79452
rect 6116 79392 6180 79396
rect 6196 79452 6260 79456
rect 6196 79396 6200 79452
rect 6200 79396 6256 79452
rect 6256 79396 6260 79452
rect 6196 79392 6260 79396
rect 87100 79452 87164 79456
rect 87100 79396 87104 79452
rect 87104 79396 87160 79452
rect 87160 79396 87164 79452
rect 87100 79392 87164 79396
rect 87180 79452 87244 79456
rect 87180 79396 87184 79452
rect 87184 79396 87240 79452
rect 87240 79396 87244 79452
rect 87180 79392 87244 79396
rect 87260 79452 87324 79456
rect 87260 79396 87264 79452
rect 87264 79396 87320 79452
rect 87320 79396 87324 79452
rect 87260 79392 87324 79396
rect 87340 79452 87404 79456
rect 87340 79396 87344 79452
rect 87344 79396 87400 79452
rect 87400 79396 87404 79452
rect 87340 79392 87404 79396
rect 6692 78908 6756 78912
rect 6692 78852 6696 78908
rect 6696 78852 6752 78908
rect 6752 78852 6756 78908
rect 6692 78848 6756 78852
rect 6772 78908 6836 78912
rect 6772 78852 6776 78908
rect 6776 78852 6832 78908
rect 6832 78852 6836 78908
rect 6772 78848 6836 78852
rect 6852 78908 6916 78912
rect 6852 78852 6856 78908
rect 6856 78852 6912 78908
rect 6912 78852 6916 78908
rect 6852 78848 6916 78852
rect 6932 78908 6996 78912
rect 6932 78852 6936 78908
rect 6936 78852 6992 78908
rect 6992 78852 6996 78908
rect 6932 78848 6996 78852
rect 87836 78908 87900 78912
rect 87836 78852 87840 78908
rect 87840 78852 87896 78908
rect 87896 78852 87900 78908
rect 87836 78848 87900 78852
rect 87916 78908 87980 78912
rect 87916 78852 87920 78908
rect 87920 78852 87976 78908
rect 87976 78852 87980 78908
rect 87916 78848 87980 78852
rect 87996 78908 88060 78912
rect 87996 78852 88000 78908
rect 88000 78852 88056 78908
rect 88056 78852 88060 78908
rect 87996 78848 88060 78852
rect 88076 78908 88140 78912
rect 88076 78852 88080 78908
rect 88080 78852 88136 78908
rect 88136 78852 88140 78908
rect 88076 78848 88140 78852
rect 5956 78364 6020 78368
rect 5956 78308 5960 78364
rect 5960 78308 6016 78364
rect 6016 78308 6020 78364
rect 5956 78304 6020 78308
rect 6036 78364 6100 78368
rect 6036 78308 6040 78364
rect 6040 78308 6096 78364
rect 6096 78308 6100 78364
rect 6036 78304 6100 78308
rect 6116 78364 6180 78368
rect 6116 78308 6120 78364
rect 6120 78308 6176 78364
rect 6176 78308 6180 78364
rect 6116 78304 6180 78308
rect 6196 78364 6260 78368
rect 6196 78308 6200 78364
rect 6200 78308 6256 78364
rect 6256 78308 6260 78364
rect 6196 78304 6260 78308
rect 87100 78364 87164 78368
rect 87100 78308 87104 78364
rect 87104 78308 87160 78364
rect 87160 78308 87164 78364
rect 87100 78304 87164 78308
rect 87180 78364 87244 78368
rect 87180 78308 87184 78364
rect 87184 78308 87240 78364
rect 87240 78308 87244 78364
rect 87180 78304 87244 78308
rect 87260 78364 87324 78368
rect 87260 78308 87264 78364
rect 87264 78308 87320 78364
rect 87320 78308 87324 78364
rect 87260 78304 87324 78308
rect 87340 78364 87404 78368
rect 87340 78308 87344 78364
rect 87344 78308 87400 78364
rect 87400 78308 87404 78364
rect 87340 78304 87404 78308
rect 6692 77820 6756 77824
rect 6692 77764 6696 77820
rect 6696 77764 6752 77820
rect 6752 77764 6756 77820
rect 6692 77760 6756 77764
rect 6772 77820 6836 77824
rect 6772 77764 6776 77820
rect 6776 77764 6832 77820
rect 6832 77764 6836 77820
rect 6772 77760 6836 77764
rect 6852 77820 6916 77824
rect 6852 77764 6856 77820
rect 6856 77764 6912 77820
rect 6912 77764 6916 77820
rect 6852 77760 6916 77764
rect 6932 77820 6996 77824
rect 6932 77764 6936 77820
rect 6936 77764 6992 77820
rect 6992 77764 6996 77820
rect 6932 77760 6996 77764
rect 87836 77820 87900 77824
rect 87836 77764 87840 77820
rect 87840 77764 87896 77820
rect 87896 77764 87900 77820
rect 87836 77760 87900 77764
rect 87916 77820 87980 77824
rect 87916 77764 87920 77820
rect 87920 77764 87976 77820
rect 87976 77764 87980 77820
rect 87916 77760 87980 77764
rect 87996 77820 88060 77824
rect 87996 77764 88000 77820
rect 88000 77764 88056 77820
rect 88056 77764 88060 77820
rect 87996 77760 88060 77764
rect 88076 77820 88140 77824
rect 88076 77764 88080 77820
rect 88080 77764 88136 77820
rect 88136 77764 88140 77820
rect 88076 77760 88140 77764
rect 5956 77276 6020 77280
rect 5956 77220 5960 77276
rect 5960 77220 6016 77276
rect 6016 77220 6020 77276
rect 5956 77216 6020 77220
rect 6036 77276 6100 77280
rect 6036 77220 6040 77276
rect 6040 77220 6096 77276
rect 6096 77220 6100 77276
rect 6036 77216 6100 77220
rect 6116 77276 6180 77280
rect 6116 77220 6120 77276
rect 6120 77220 6176 77276
rect 6176 77220 6180 77276
rect 6116 77216 6180 77220
rect 6196 77276 6260 77280
rect 6196 77220 6200 77276
rect 6200 77220 6256 77276
rect 6256 77220 6260 77276
rect 6196 77216 6260 77220
rect 87100 77276 87164 77280
rect 87100 77220 87104 77276
rect 87104 77220 87160 77276
rect 87160 77220 87164 77276
rect 87100 77216 87164 77220
rect 87180 77276 87244 77280
rect 87180 77220 87184 77276
rect 87184 77220 87240 77276
rect 87240 77220 87244 77276
rect 87180 77216 87244 77220
rect 87260 77276 87324 77280
rect 87260 77220 87264 77276
rect 87264 77220 87320 77276
rect 87320 77220 87324 77276
rect 87260 77216 87324 77220
rect 87340 77276 87404 77280
rect 87340 77220 87344 77276
rect 87344 77220 87400 77276
rect 87400 77220 87404 77276
rect 87340 77216 87404 77220
rect 6692 76732 6756 76736
rect 6692 76676 6696 76732
rect 6696 76676 6752 76732
rect 6752 76676 6756 76732
rect 6692 76672 6756 76676
rect 6772 76732 6836 76736
rect 6772 76676 6776 76732
rect 6776 76676 6832 76732
rect 6832 76676 6836 76732
rect 6772 76672 6836 76676
rect 6852 76732 6916 76736
rect 6852 76676 6856 76732
rect 6856 76676 6912 76732
rect 6912 76676 6916 76732
rect 6852 76672 6916 76676
rect 6932 76732 6996 76736
rect 6932 76676 6936 76732
rect 6936 76676 6992 76732
rect 6992 76676 6996 76732
rect 6932 76672 6996 76676
rect 87836 76732 87900 76736
rect 87836 76676 87840 76732
rect 87840 76676 87896 76732
rect 87896 76676 87900 76732
rect 87836 76672 87900 76676
rect 87916 76732 87980 76736
rect 87916 76676 87920 76732
rect 87920 76676 87976 76732
rect 87976 76676 87980 76732
rect 87916 76672 87980 76676
rect 87996 76732 88060 76736
rect 87996 76676 88000 76732
rect 88000 76676 88056 76732
rect 88056 76676 88060 76732
rect 87996 76672 88060 76676
rect 88076 76732 88140 76736
rect 88076 76676 88080 76732
rect 88080 76676 88136 76732
rect 88136 76676 88140 76732
rect 88076 76672 88140 76676
rect 5956 76188 6020 76192
rect 5956 76132 5960 76188
rect 5960 76132 6016 76188
rect 6016 76132 6020 76188
rect 5956 76128 6020 76132
rect 6036 76188 6100 76192
rect 6036 76132 6040 76188
rect 6040 76132 6096 76188
rect 6096 76132 6100 76188
rect 6036 76128 6100 76132
rect 6116 76188 6180 76192
rect 6116 76132 6120 76188
rect 6120 76132 6176 76188
rect 6176 76132 6180 76188
rect 6116 76128 6180 76132
rect 6196 76188 6260 76192
rect 6196 76132 6200 76188
rect 6200 76132 6256 76188
rect 6256 76132 6260 76188
rect 6196 76128 6260 76132
rect 87100 76188 87164 76192
rect 87100 76132 87104 76188
rect 87104 76132 87160 76188
rect 87160 76132 87164 76188
rect 87100 76128 87164 76132
rect 87180 76188 87244 76192
rect 87180 76132 87184 76188
rect 87184 76132 87240 76188
rect 87240 76132 87244 76188
rect 87180 76128 87244 76132
rect 87260 76188 87324 76192
rect 87260 76132 87264 76188
rect 87264 76132 87320 76188
rect 87320 76132 87324 76188
rect 87260 76128 87324 76132
rect 87340 76188 87404 76192
rect 87340 76132 87344 76188
rect 87344 76132 87400 76188
rect 87400 76132 87404 76188
rect 87340 76128 87404 76132
rect 6692 75644 6756 75648
rect 6692 75588 6696 75644
rect 6696 75588 6752 75644
rect 6752 75588 6756 75644
rect 6692 75584 6756 75588
rect 6772 75644 6836 75648
rect 6772 75588 6776 75644
rect 6776 75588 6832 75644
rect 6832 75588 6836 75644
rect 6772 75584 6836 75588
rect 6852 75644 6916 75648
rect 6852 75588 6856 75644
rect 6856 75588 6912 75644
rect 6912 75588 6916 75644
rect 6852 75584 6916 75588
rect 6932 75644 6996 75648
rect 6932 75588 6936 75644
rect 6936 75588 6992 75644
rect 6992 75588 6996 75644
rect 6932 75584 6996 75588
rect 87836 75644 87900 75648
rect 87836 75588 87840 75644
rect 87840 75588 87896 75644
rect 87896 75588 87900 75644
rect 87836 75584 87900 75588
rect 87916 75644 87980 75648
rect 87916 75588 87920 75644
rect 87920 75588 87976 75644
rect 87976 75588 87980 75644
rect 87916 75584 87980 75588
rect 87996 75644 88060 75648
rect 87996 75588 88000 75644
rect 88000 75588 88056 75644
rect 88056 75588 88060 75644
rect 87996 75584 88060 75588
rect 88076 75644 88140 75648
rect 88076 75588 88080 75644
rect 88080 75588 88136 75644
rect 88136 75588 88140 75644
rect 88076 75584 88140 75588
rect 5956 75100 6020 75104
rect 5956 75044 5960 75100
rect 5960 75044 6016 75100
rect 6016 75044 6020 75100
rect 5956 75040 6020 75044
rect 6036 75100 6100 75104
rect 6036 75044 6040 75100
rect 6040 75044 6096 75100
rect 6096 75044 6100 75100
rect 6036 75040 6100 75044
rect 6116 75100 6180 75104
rect 6116 75044 6120 75100
rect 6120 75044 6176 75100
rect 6176 75044 6180 75100
rect 6116 75040 6180 75044
rect 6196 75100 6260 75104
rect 6196 75044 6200 75100
rect 6200 75044 6256 75100
rect 6256 75044 6260 75100
rect 6196 75040 6260 75044
rect 87100 75100 87164 75104
rect 87100 75044 87104 75100
rect 87104 75044 87160 75100
rect 87160 75044 87164 75100
rect 87100 75040 87164 75044
rect 87180 75100 87244 75104
rect 87180 75044 87184 75100
rect 87184 75044 87240 75100
rect 87240 75044 87244 75100
rect 87180 75040 87244 75044
rect 87260 75100 87324 75104
rect 87260 75044 87264 75100
rect 87264 75044 87320 75100
rect 87320 75044 87324 75100
rect 87260 75040 87324 75044
rect 87340 75100 87404 75104
rect 87340 75044 87344 75100
rect 87344 75044 87400 75100
rect 87400 75044 87404 75100
rect 87340 75040 87404 75044
rect 6692 74556 6756 74560
rect 6692 74500 6696 74556
rect 6696 74500 6752 74556
rect 6752 74500 6756 74556
rect 6692 74496 6756 74500
rect 6772 74556 6836 74560
rect 6772 74500 6776 74556
rect 6776 74500 6832 74556
rect 6832 74500 6836 74556
rect 6772 74496 6836 74500
rect 6852 74556 6916 74560
rect 6852 74500 6856 74556
rect 6856 74500 6912 74556
rect 6912 74500 6916 74556
rect 6852 74496 6916 74500
rect 6932 74556 6996 74560
rect 6932 74500 6936 74556
rect 6936 74500 6992 74556
rect 6992 74500 6996 74556
rect 6932 74496 6996 74500
rect 87836 74556 87900 74560
rect 87836 74500 87840 74556
rect 87840 74500 87896 74556
rect 87896 74500 87900 74556
rect 87836 74496 87900 74500
rect 87916 74556 87980 74560
rect 87916 74500 87920 74556
rect 87920 74500 87976 74556
rect 87976 74500 87980 74556
rect 87916 74496 87980 74500
rect 87996 74556 88060 74560
rect 87996 74500 88000 74556
rect 88000 74500 88056 74556
rect 88056 74500 88060 74556
rect 87996 74496 88060 74500
rect 88076 74556 88140 74560
rect 88076 74500 88080 74556
rect 88080 74500 88136 74556
rect 88136 74500 88140 74556
rect 88076 74496 88140 74500
rect 5956 74012 6020 74016
rect 5956 73956 5960 74012
rect 5960 73956 6016 74012
rect 6016 73956 6020 74012
rect 5956 73952 6020 73956
rect 6036 74012 6100 74016
rect 6036 73956 6040 74012
rect 6040 73956 6096 74012
rect 6096 73956 6100 74012
rect 6036 73952 6100 73956
rect 6116 74012 6180 74016
rect 6116 73956 6120 74012
rect 6120 73956 6176 74012
rect 6176 73956 6180 74012
rect 6116 73952 6180 73956
rect 6196 74012 6260 74016
rect 6196 73956 6200 74012
rect 6200 73956 6256 74012
rect 6256 73956 6260 74012
rect 6196 73952 6260 73956
rect 87100 74012 87164 74016
rect 87100 73956 87104 74012
rect 87104 73956 87160 74012
rect 87160 73956 87164 74012
rect 87100 73952 87164 73956
rect 87180 74012 87244 74016
rect 87180 73956 87184 74012
rect 87184 73956 87240 74012
rect 87240 73956 87244 74012
rect 87180 73952 87244 73956
rect 87260 74012 87324 74016
rect 87260 73956 87264 74012
rect 87264 73956 87320 74012
rect 87320 73956 87324 74012
rect 87260 73952 87324 73956
rect 87340 74012 87404 74016
rect 87340 73956 87344 74012
rect 87344 73956 87400 74012
rect 87400 73956 87404 74012
rect 87340 73952 87404 73956
rect 6692 73468 6756 73472
rect 6692 73412 6696 73468
rect 6696 73412 6752 73468
rect 6752 73412 6756 73468
rect 6692 73408 6756 73412
rect 6772 73468 6836 73472
rect 6772 73412 6776 73468
rect 6776 73412 6832 73468
rect 6832 73412 6836 73468
rect 6772 73408 6836 73412
rect 6852 73468 6916 73472
rect 6852 73412 6856 73468
rect 6856 73412 6912 73468
rect 6912 73412 6916 73468
rect 6852 73408 6916 73412
rect 6932 73468 6996 73472
rect 6932 73412 6936 73468
rect 6936 73412 6992 73468
rect 6992 73412 6996 73468
rect 6932 73408 6996 73412
rect 87836 73468 87900 73472
rect 87836 73412 87840 73468
rect 87840 73412 87896 73468
rect 87896 73412 87900 73468
rect 87836 73408 87900 73412
rect 87916 73468 87980 73472
rect 87916 73412 87920 73468
rect 87920 73412 87976 73468
rect 87976 73412 87980 73468
rect 87916 73408 87980 73412
rect 87996 73468 88060 73472
rect 87996 73412 88000 73468
rect 88000 73412 88056 73468
rect 88056 73412 88060 73468
rect 87996 73408 88060 73412
rect 88076 73468 88140 73472
rect 88076 73412 88080 73468
rect 88080 73412 88136 73468
rect 88136 73412 88140 73468
rect 88076 73408 88140 73412
rect 5956 72924 6020 72928
rect 5956 72868 5960 72924
rect 5960 72868 6016 72924
rect 6016 72868 6020 72924
rect 5956 72864 6020 72868
rect 6036 72924 6100 72928
rect 6036 72868 6040 72924
rect 6040 72868 6096 72924
rect 6096 72868 6100 72924
rect 6036 72864 6100 72868
rect 6116 72924 6180 72928
rect 6116 72868 6120 72924
rect 6120 72868 6176 72924
rect 6176 72868 6180 72924
rect 6116 72864 6180 72868
rect 6196 72924 6260 72928
rect 6196 72868 6200 72924
rect 6200 72868 6256 72924
rect 6256 72868 6260 72924
rect 6196 72864 6260 72868
rect 87100 72924 87164 72928
rect 87100 72868 87104 72924
rect 87104 72868 87160 72924
rect 87160 72868 87164 72924
rect 87100 72864 87164 72868
rect 87180 72924 87244 72928
rect 87180 72868 87184 72924
rect 87184 72868 87240 72924
rect 87240 72868 87244 72924
rect 87180 72864 87244 72868
rect 87260 72924 87324 72928
rect 87260 72868 87264 72924
rect 87264 72868 87320 72924
rect 87320 72868 87324 72924
rect 87260 72864 87324 72868
rect 87340 72924 87404 72928
rect 87340 72868 87344 72924
rect 87344 72868 87400 72924
rect 87400 72868 87404 72924
rect 87340 72864 87404 72868
rect 6692 72380 6756 72384
rect 6692 72324 6696 72380
rect 6696 72324 6752 72380
rect 6752 72324 6756 72380
rect 6692 72320 6756 72324
rect 6772 72380 6836 72384
rect 6772 72324 6776 72380
rect 6776 72324 6832 72380
rect 6832 72324 6836 72380
rect 6772 72320 6836 72324
rect 6852 72380 6916 72384
rect 6852 72324 6856 72380
rect 6856 72324 6912 72380
rect 6912 72324 6916 72380
rect 6852 72320 6916 72324
rect 6932 72380 6996 72384
rect 6932 72324 6936 72380
rect 6936 72324 6992 72380
rect 6992 72324 6996 72380
rect 6932 72320 6996 72324
rect 87836 72380 87900 72384
rect 87836 72324 87840 72380
rect 87840 72324 87896 72380
rect 87896 72324 87900 72380
rect 87836 72320 87900 72324
rect 87916 72380 87980 72384
rect 87916 72324 87920 72380
rect 87920 72324 87976 72380
rect 87976 72324 87980 72380
rect 87916 72320 87980 72324
rect 87996 72380 88060 72384
rect 87996 72324 88000 72380
rect 88000 72324 88056 72380
rect 88056 72324 88060 72380
rect 87996 72320 88060 72324
rect 88076 72380 88140 72384
rect 88076 72324 88080 72380
rect 88080 72324 88136 72380
rect 88136 72324 88140 72380
rect 88076 72320 88140 72324
rect 5956 71836 6020 71840
rect 5956 71780 5960 71836
rect 5960 71780 6016 71836
rect 6016 71780 6020 71836
rect 5956 71776 6020 71780
rect 6036 71836 6100 71840
rect 6036 71780 6040 71836
rect 6040 71780 6096 71836
rect 6096 71780 6100 71836
rect 6036 71776 6100 71780
rect 6116 71836 6180 71840
rect 6116 71780 6120 71836
rect 6120 71780 6176 71836
rect 6176 71780 6180 71836
rect 6116 71776 6180 71780
rect 6196 71836 6260 71840
rect 6196 71780 6200 71836
rect 6200 71780 6256 71836
rect 6256 71780 6260 71836
rect 6196 71776 6260 71780
rect 87100 71836 87164 71840
rect 87100 71780 87104 71836
rect 87104 71780 87160 71836
rect 87160 71780 87164 71836
rect 87100 71776 87164 71780
rect 87180 71836 87244 71840
rect 87180 71780 87184 71836
rect 87184 71780 87240 71836
rect 87240 71780 87244 71836
rect 87180 71776 87244 71780
rect 87260 71836 87324 71840
rect 87260 71780 87264 71836
rect 87264 71780 87320 71836
rect 87320 71780 87324 71836
rect 87260 71776 87324 71780
rect 87340 71836 87404 71840
rect 87340 71780 87344 71836
rect 87344 71780 87400 71836
rect 87400 71780 87404 71836
rect 87340 71776 87404 71780
rect 6692 71292 6756 71296
rect 6692 71236 6696 71292
rect 6696 71236 6752 71292
rect 6752 71236 6756 71292
rect 6692 71232 6756 71236
rect 6772 71292 6836 71296
rect 6772 71236 6776 71292
rect 6776 71236 6832 71292
rect 6832 71236 6836 71292
rect 6772 71232 6836 71236
rect 6852 71292 6916 71296
rect 6852 71236 6856 71292
rect 6856 71236 6912 71292
rect 6912 71236 6916 71292
rect 6852 71232 6916 71236
rect 6932 71292 6996 71296
rect 6932 71236 6936 71292
rect 6936 71236 6992 71292
rect 6992 71236 6996 71292
rect 6932 71232 6996 71236
rect 87836 71292 87900 71296
rect 87836 71236 87840 71292
rect 87840 71236 87896 71292
rect 87896 71236 87900 71292
rect 87836 71232 87900 71236
rect 87916 71292 87980 71296
rect 87916 71236 87920 71292
rect 87920 71236 87976 71292
rect 87976 71236 87980 71292
rect 87916 71232 87980 71236
rect 87996 71292 88060 71296
rect 87996 71236 88000 71292
rect 88000 71236 88056 71292
rect 88056 71236 88060 71292
rect 87996 71232 88060 71236
rect 88076 71292 88140 71296
rect 88076 71236 88080 71292
rect 88080 71236 88136 71292
rect 88136 71236 88140 71292
rect 88076 71232 88140 71236
rect 5956 70748 6020 70752
rect 5956 70692 5960 70748
rect 5960 70692 6016 70748
rect 6016 70692 6020 70748
rect 5956 70688 6020 70692
rect 6036 70748 6100 70752
rect 6036 70692 6040 70748
rect 6040 70692 6096 70748
rect 6096 70692 6100 70748
rect 6036 70688 6100 70692
rect 6116 70748 6180 70752
rect 6116 70692 6120 70748
rect 6120 70692 6176 70748
rect 6176 70692 6180 70748
rect 6116 70688 6180 70692
rect 6196 70748 6260 70752
rect 6196 70692 6200 70748
rect 6200 70692 6256 70748
rect 6256 70692 6260 70748
rect 6196 70688 6260 70692
rect 87100 70748 87164 70752
rect 87100 70692 87104 70748
rect 87104 70692 87160 70748
rect 87160 70692 87164 70748
rect 87100 70688 87164 70692
rect 87180 70748 87244 70752
rect 87180 70692 87184 70748
rect 87184 70692 87240 70748
rect 87240 70692 87244 70748
rect 87180 70688 87244 70692
rect 87260 70748 87324 70752
rect 87260 70692 87264 70748
rect 87264 70692 87320 70748
rect 87320 70692 87324 70748
rect 87260 70688 87324 70692
rect 87340 70748 87404 70752
rect 87340 70692 87344 70748
rect 87344 70692 87400 70748
rect 87400 70692 87404 70748
rect 87340 70688 87404 70692
rect 6692 70204 6756 70208
rect 6692 70148 6696 70204
rect 6696 70148 6752 70204
rect 6752 70148 6756 70204
rect 6692 70144 6756 70148
rect 6772 70204 6836 70208
rect 6772 70148 6776 70204
rect 6776 70148 6832 70204
rect 6832 70148 6836 70204
rect 6772 70144 6836 70148
rect 6852 70204 6916 70208
rect 6852 70148 6856 70204
rect 6856 70148 6912 70204
rect 6912 70148 6916 70204
rect 6852 70144 6916 70148
rect 6932 70204 6996 70208
rect 6932 70148 6936 70204
rect 6936 70148 6992 70204
rect 6992 70148 6996 70204
rect 6932 70144 6996 70148
rect 87836 70204 87900 70208
rect 87836 70148 87840 70204
rect 87840 70148 87896 70204
rect 87896 70148 87900 70204
rect 87836 70144 87900 70148
rect 87916 70204 87980 70208
rect 87916 70148 87920 70204
rect 87920 70148 87976 70204
rect 87976 70148 87980 70204
rect 87916 70144 87980 70148
rect 87996 70204 88060 70208
rect 87996 70148 88000 70204
rect 88000 70148 88056 70204
rect 88056 70148 88060 70204
rect 87996 70144 88060 70148
rect 88076 70204 88140 70208
rect 88076 70148 88080 70204
rect 88080 70148 88136 70204
rect 88136 70148 88140 70204
rect 88076 70144 88140 70148
rect 5956 69660 6020 69664
rect 5956 69604 5960 69660
rect 5960 69604 6016 69660
rect 6016 69604 6020 69660
rect 5956 69600 6020 69604
rect 6036 69660 6100 69664
rect 6036 69604 6040 69660
rect 6040 69604 6096 69660
rect 6096 69604 6100 69660
rect 6036 69600 6100 69604
rect 6116 69660 6180 69664
rect 6116 69604 6120 69660
rect 6120 69604 6176 69660
rect 6176 69604 6180 69660
rect 6116 69600 6180 69604
rect 6196 69660 6260 69664
rect 6196 69604 6200 69660
rect 6200 69604 6256 69660
rect 6256 69604 6260 69660
rect 6196 69600 6260 69604
rect 87100 69660 87164 69664
rect 87100 69604 87104 69660
rect 87104 69604 87160 69660
rect 87160 69604 87164 69660
rect 87100 69600 87164 69604
rect 87180 69660 87244 69664
rect 87180 69604 87184 69660
rect 87184 69604 87240 69660
rect 87240 69604 87244 69660
rect 87180 69600 87244 69604
rect 87260 69660 87324 69664
rect 87260 69604 87264 69660
rect 87264 69604 87320 69660
rect 87320 69604 87324 69660
rect 87260 69600 87324 69604
rect 87340 69660 87404 69664
rect 87340 69604 87344 69660
rect 87344 69604 87400 69660
rect 87400 69604 87404 69660
rect 87340 69600 87404 69604
rect 6692 69116 6756 69120
rect 6692 69060 6696 69116
rect 6696 69060 6752 69116
rect 6752 69060 6756 69116
rect 6692 69056 6756 69060
rect 6772 69116 6836 69120
rect 6772 69060 6776 69116
rect 6776 69060 6832 69116
rect 6832 69060 6836 69116
rect 6772 69056 6836 69060
rect 6852 69116 6916 69120
rect 6852 69060 6856 69116
rect 6856 69060 6912 69116
rect 6912 69060 6916 69116
rect 6852 69056 6916 69060
rect 6932 69116 6996 69120
rect 6932 69060 6936 69116
rect 6936 69060 6992 69116
rect 6992 69060 6996 69116
rect 6932 69056 6996 69060
rect 87836 69116 87900 69120
rect 87836 69060 87840 69116
rect 87840 69060 87896 69116
rect 87896 69060 87900 69116
rect 87836 69056 87900 69060
rect 87916 69116 87980 69120
rect 87916 69060 87920 69116
rect 87920 69060 87976 69116
rect 87976 69060 87980 69116
rect 87916 69056 87980 69060
rect 87996 69116 88060 69120
rect 87996 69060 88000 69116
rect 88000 69060 88056 69116
rect 88056 69060 88060 69116
rect 87996 69056 88060 69060
rect 88076 69116 88140 69120
rect 88076 69060 88080 69116
rect 88080 69060 88136 69116
rect 88136 69060 88140 69116
rect 88076 69056 88140 69060
rect 5956 68572 6020 68576
rect 5956 68516 5960 68572
rect 5960 68516 6016 68572
rect 6016 68516 6020 68572
rect 5956 68512 6020 68516
rect 6036 68572 6100 68576
rect 6036 68516 6040 68572
rect 6040 68516 6096 68572
rect 6096 68516 6100 68572
rect 6036 68512 6100 68516
rect 6116 68572 6180 68576
rect 6116 68516 6120 68572
rect 6120 68516 6176 68572
rect 6176 68516 6180 68572
rect 6116 68512 6180 68516
rect 6196 68572 6260 68576
rect 6196 68516 6200 68572
rect 6200 68516 6256 68572
rect 6256 68516 6260 68572
rect 6196 68512 6260 68516
rect 87100 68572 87164 68576
rect 87100 68516 87104 68572
rect 87104 68516 87160 68572
rect 87160 68516 87164 68572
rect 87100 68512 87164 68516
rect 87180 68572 87244 68576
rect 87180 68516 87184 68572
rect 87184 68516 87240 68572
rect 87240 68516 87244 68572
rect 87180 68512 87244 68516
rect 87260 68572 87324 68576
rect 87260 68516 87264 68572
rect 87264 68516 87320 68572
rect 87320 68516 87324 68572
rect 87260 68512 87324 68516
rect 87340 68572 87404 68576
rect 87340 68516 87344 68572
rect 87344 68516 87400 68572
rect 87400 68516 87404 68572
rect 87340 68512 87404 68516
rect 6692 68028 6756 68032
rect 6692 67972 6696 68028
rect 6696 67972 6752 68028
rect 6752 67972 6756 68028
rect 6692 67968 6756 67972
rect 6772 68028 6836 68032
rect 6772 67972 6776 68028
rect 6776 67972 6832 68028
rect 6832 67972 6836 68028
rect 6772 67968 6836 67972
rect 6852 68028 6916 68032
rect 6852 67972 6856 68028
rect 6856 67972 6912 68028
rect 6912 67972 6916 68028
rect 6852 67968 6916 67972
rect 6932 68028 6996 68032
rect 6932 67972 6936 68028
rect 6936 67972 6992 68028
rect 6992 67972 6996 68028
rect 6932 67968 6996 67972
rect 87836 68028 87900 68032
rect 87836 67972 87840 68028
rect 87840 67972 87896 68028
rect 87896 67972 87900 68028
rect 87836 67968 87900 67972
rect 87916 68028 87980 68032
rect 87916 67972 87920 68028
rect 87920 67972 87976 68028
rect 87976 67972 87980 68028
rect 87916 67968 87980 67972
rect 87996 68028 88060 68032
rect 87996 67972 88000 68028
rect 88000 67972 88056 68028
rect 88056 67972 88060 68028
rect 87996 67968 88060 67972
rect 88076 68028 88140 68032
rect 88076 67972 88080 68028
rect 88080 67972 88136 68028
rect 88136 67972 88140 68028
rect 88076 67968 88140 67972
rect 5956 67484 6020 67488
rect 5956 67428 5960 67484
rect 5960 67428 6016 67484
rect 6016 67428 6020 67484
rect 5956 67424 6020 67428
rect 6036 67484 6100 67488
rect 6036 67428 6040 67484
rect 6040 67428 6096 67484
rect 6096 67428 6100 67484
rect 6036 67424 6100 67428
rect 6116 67484 6180 67488
rect 6116 67428 6120 67484
rect 6120 67428 6176 67484
rect 6176 67428 6180 67484
rect 6116 67424 6180 67428
rect 6196 67484 6260 67488
rect 6196 67428 6200 67484
rect 6200 67428 6256 67484
rect 6256 67428 6260 67484
rect 6196 67424 6260 67428
rect 87100 67484 87164 67488
rect 87100 67428 87104 67484
rect 87104 67428 87160 67484
rect 87160 67428 87164 67484
rect 87100 67424 87164 67428
rect 87180 67484 87244 67488
rect 87180 67428 87184 67484
rect 87184 67428 87240 67484
rect 87240 67428 87244 67484
rect 87180 67424 87244 67428
rect 87260 67484 87324 67488
rect 87260 67428 87264 67484
rect 87264 67428 87320 67484
rect 87320 67428 87324 67484
rect 87260 67424 87324 67428
rect 87340 67484 87404 67488
rect 87340 67428 87344 67484
rect 87344 67428 87400 67484
rect 87400 67428 87404 67484
rect 87340 67424 87404 67428
rect 6692 66940 6756 66944
rect 6692 66884 6696 66940
rect 6696 66884 6752 66940
rect 6752 66884 6756 66940
rect 6692 66880 6756 66884
rect 6772 66940 6836 66944
rect 6772 66884 6776 66940
rect 6776 66884 6832 66940
rect 6832 66884 6836 66940
rect 6772 66880 6836 66884
rect 6852 66940 6916 66944
rect 6852 66884 6856 66940
rect 6856 66884 6912 66940
rect 6912 66884 6916 66940
rect 6852 66880 6916 66884
rect 6932 66940 6996 66944
rect 6932 66884 6936 66940
rect 6936 66884 6992 66940
rect 6992 66884 6996 66940
rect 6932 66880 6996 66884
rect 87836 66940 87900 66944
rect 87836 66884 87840 66940
rect 87840 66884 87896 66940
rect 87896 66884 87900 66940
rect 87836 66880 87900 66884
rect 87916 66940 87980 66944
rect 87916 66884 87920 66940
rect 87920 66884 87976 66940
rect 87976 66884 87980 66940
rect 87916 66880 87980 66884
rect 87996 66940 88060 66944
rect 87996 66884 88000 66940
rect 88000 66884 88056 66940
rect 88056 66884 88060 66940
rect 87996 66880 88060 66884
rect 88076 66940 88140 66944
rect 88076 66884 88080 66940
rect 88080 66884 88136 66940
rect 88136 66884 88140 66940
rect 88076 66880 88140 66884
rect 5956 66396 6020 66400
rect 5956 66340 5960 66396
rect 5960 66340 6016 66396
rect 6016 66340 6020 66396
rect 5956 66336 6020 66340
rect 6036 66396 6100 66400
rect 6036 66340 6040 66396
rect 6040 66340 6096 66396
rect 6096 66340 6100 66396
rect 6036 66336 6100 66340
rect 6116 66396 6180 66400
rect 6116 66340 6120 66396
rect 6120 66340 6176 66396
rect 6176 66340 6180 66396
rect 6116 66336 6180 66340
rect 6196 66396 6260 66400
rect 6196 66340 6200 66396
rect 6200 66340 6256 66396
rect 6256 66340 6260 66396
rect 6196 66336 6260 66340
rect 87100 66396 87164 66400
rect 87100 66340 87104 66396
rect 87104 66340 87160 66396
rect 87160 66340 87164 66396
rect 87100 66336 87164 66340
rect 87180 66396 87244 66400
rect 87180 66340 87184 66396
rect 87184 66340 87240 66396
rect 87240 66340 87244 66396
rect 87180 66336 87244 66340
rect 87260 66396 87324 66400
rect 87260 66340 87264 66396
rect 87264 66340 87320 66396
rect 87320 66340 87324 66396
rect 87260 66336 87324 66340
rect 87340 66396 87404 66400
rect 87340 66340 87344 66396
rect 87344 66340 87400 66396
rect 87400 66340 87404 66396
rect 87340 66336 87404 66340
rect 6692 65852 6756 65856
rect 6692 65796 6696 65852
rect 6696 65796 6752 65852
rect 6752 65796 6756 65852
rect 6692 65792 6756 65796
rect 6772 65852 6836 65856
rect 6772 65796 6776 65852
rect 6776 65796 6832 65852
rect 6832 65796 6836 65852
rect 6772 65792 6836 65796
rect 6852 65852 6916 65856
rect 6852 65796 6856 65852
rect 6856 65796 6912 65852
rect 6912 65796 6916 65852
rect 6852 65792 6916 65796
rect 6932 65852 6996 65856
rect 6932 65796 6936 65852
rect 6936 65796 6992 65852
rect 6992 65796 6996 65852
rect 6932 65792 6996 65796
rect 87836 65852 87900 65856
rect 87836 65796 87840 65852
rect 87840 65796 87896 65852
rect 87896 65796 87900 65852
rect 87836 65792 87900 65796
rect 87916 65852 87980 65856
rect 87916 65796 87920 65852
rect 87920 65796 87976 65852
rect 87976 65796 87980 65852
rect 87916 65792 87980 65796
rect 87996 65852 88060 65856
rect 87996 65796 88000 65852
rect 88000 65796 88056 65852
rect 88056 65796 88060 65852
rect 87996 65792 88060 65796
rect 88076 65852 88140 65856
rect 88076 65796 88080 65852
rect 88080 65796 88136 65852
rect 88136 65796 88140 65852
rect 88076 65792 88140 65796
rect 5956 65308 6020 65312
rect 5956 65252 5960 65308
rect 5960 65252 6016 65308
rect 6016 65252 6020 65308
rect 5956 65248 6020 65252
rect 6036 65308 6100 65312
rect 6036 65252 6040 65308
rect 6040 65252 6096 65308
rect 6096 65252 6100 65308
rect 6036 65248 6100 65252
rect 6116 65308 6180 65312
rect 6116 65252 6120 65308
rect 6120 65252 6176 65308
rect 6176 65252 6180 65308
rect 6116 65248 6180 65252
rect 6196 65308 6260 65312
rect 6196 65252 6200 65308
rect 6200 65252 6256 65308
rect 6256 65252 6260 65308
rect 6196 65248 6260 65252
rect 87100 65308 87164 65312
rect 87100 65252 87104 65308
rect 87104 65252 87160 65308
rect 87160 65252 87164 65308
rect 87100 65248 87164 65252
rect 87180 65308 87244 65312
rect 87180 65252 87184 65308
rect 87184 65252 87240 65308
rect 87240 65252 87244 65308
rect 87180 65248 87244 65252
rect 87260 65308 87324 65312
rect 87260 65252 87264 65308
rect 87264 65252 87320 65308
rect 87320 65252 87324 65308
rect 87260 65248 87324 65252
rect 87340 65308 87404 65312
rect 87340 65252 87344 65308
rect 87344 65252 87400 65308
rect 87400 65252 87404 65308
rect 87340 65248 87404 65252
rect 6692 64764 6756 64768
rect 6692 64708 6696 64764
rect 6696 64708 6752 64764
rect 6752 64708 6756 64764
rect 6692 64704 6756 64708
rect 6772 64764 6836 64768
rect 6772 64708 6776 64764
rect 6776 64708 6832 64764
rect 6832 64708 6836 64764
rect 6772 64704 6836 64708
rect 6852 64764 6916 64768
rect 6852 64708 6856 64764
rect 6856 64708 6912 64764
rect 6912 64708 6916 64764
rect 6852 64704 6916 64708
rect 6932 64764 6996 64768
rect 6932 64708 6936 64764
rect 6936 64708 6992 64764
rect 6992 64708 6996 64764
rect 6932 64704 6996 64708
rect 87836 64764 87900 64768
rect 87836 64708 87840 64764
rect 87840 64708 87896 64764
rect 87896 64708 87900 64764
rect 87836 64704 87900 64708
rect 87916 64764 87980 64768
rect 87916 64708 87920 64764
rect 87920 64708 87976 64764
rect 87976 64708 87980 64764
rect 87916 64704 87980 64708
rect 87996 64764 88060 64768
rect 87996 64708 88000 64764
rect 88000 64708 88056 64764
rect 88056 64708 88060 64764
rect 87996 64704 88060 64708
rect 88076 64764 88140 64768
rect 88076 64708 88080 64764
rect 88080 64708 88136 64764
rect 88136 64708 88140 64764
rect 88076 64704 88140 64708
rect 5956 64220 6020 64224
rect 5956 64164 5960 64220
rect 5960 64164 6016 64220
rect 6016 64164 6020 64220
rect 5956 64160 6020 64164
rect 6036 64220 6100 64224
rect 6036 64164 6040 64220
rect 6040 64164 6096 64220
rect 6096 64164 6100 64220
rect 6036 64160 6100 64164
rect 6116 64220 6180 64224
rect 6116 64164 6120 64220
rect 6120 64164 6176 64220
rect 6176 64164 6180 64220
rect 6116 64160 6180 64164
rect 6196 64220 6260 64224
rect 6196 64164 6200 64220
rect 6200 64164 6256 64220
rect 6256 64164 6260 64220
rect 6196 64160 6260 64164
rect 87100 64220 87164 64224
rect 87100 64164 87104 64220
rect 87104 64164 87160 64220
rect 87160 64164 87164 64220
rect 87100 64160 87164 64164
rect 87180 64220 87244 64224
rect 87180 64164 87184 64220
rect 87184 64164 87240 64220
rect 87240 64164 87244 64220
rect 87180 64160 87244 64164
rect 87260 64220 87324 64224
rect 87260 64164 87264 64220
rect 87264 64164 87320 64220
rect 87320 64164 87324 64220
rect 87260 64160 87324 64164
rect 87340 64220 87404 64224
rect 87340 64164 87344 64220
rect 87344 64164 87400 64220
rect 87400 64164 87404 64220
rect 87340 64160 87404 64164
rect 6692 63676 6756 63680
rect 6692 63620 6696 63676
rect 6696 63620 6752 63676
rect 6752 63620 6756 63676
rect 6692 63616 6756 63620
rect 6772 63676 6836 63680
rect 6772 63620 6776 63676
rect 6776 63620 6832 63676
rect 6832 63620 6836 63676
rect 6772 63616 6836 63620
rect 6852 63676 6916 63680
rect 6852 63620 6856 63676
rect 6856 63620 6912 63676
rect 6912 63620 6916 63676
rect 6852 63616 6916 63620
rect 6932 63676 6996 63680
rect 6932 63620 6936 63676
rect 6936 63620 6992 63676
rect 6992 63620 6996 63676
rect 6932 63616 6996 63620
rect 87836 63676 87900 63680
rect 87836 63620 87840 63676
rect 87840 63620 87896 63676
rect 87896 63620 87900 63676
rect 87836 63616 87900 63620
rect 87916 63676 87980 63680
rect 87916 63620 87920 63676
rect 87920 63620 87976 63676
rect 87976 63620 87980 63676
rect 87916 63616 87980 63620
rect 87996 63676 88060 63680
rect 87996 63620 88000 63676
rect 88000 63620 88056 63676
rect 88056 63620 88060 63676
rect 87996 63616 88060 63620
rect 88076 63676 88140 63680
rect 88076 63620 88080 63676
rect 88080 63620 88136 63676
rect 88136 63620 88140 63676
rect 88076 63616 88140 63620
rect 5956 63132 6020 63136
rect 5956 63076 5960 63132
rect 5960 63076 6016 63132
rect 6016 63076 6020 63132
rect 5956 63072 6020 63076
rect 6036 63132 6100 63136
rect 6036 63076 6040 63132
rect 6040 63076 6096 63132
rect 6096 63076 6100 63132
rect 6036 63072 6100 63076
rect 6116 63132 6180 63136
rect 6116 63076 6120 63132
rect 6120 63076 6176 63132
rect 6176 63076 6180 63132
rect 6116 63072 6180 63076
rect 6196 63132 6260 63136
rect 6196 63076 6200 63132
rect 6200 63076 6256 63132
rect 6256 63076 6260 63132
rect 6196 63072 6260 63076
rect 87100 63132 87164 63136
rect 87100 63076 87104 63132
rect 87104 63076 87160 63132
rect 87160 63076 87164 63132
rect 87100 63072 87164 63076
rect 87180 63132 87244 63136
rect 87180 63076 87184 63132
rect 87184 63076 87240 63132
rect 87240 63076 87244 63132
rect 87180 63072 87244 63076
rect 87260 63132 87324 63136
rect 87260 63076 87264 63132
rect 87264 63076 87320 63132
rect 87320 63076 87324 63132
rect 87260 63072 87324 63076
rect 87340 63132 87404 63136
rect 87340 63076 87344 63132
rect 87344 63076 87400 63132
rect 87400 63076 87404 63132
rect 87340 63072 87404 63076
rect 6692 62588 6756 62592
rect 6692 62532 6696 62588
rect 6696 62532 6752 62588
rect 6752 62532 6756 62588
rect 6692 62528 6756 62532
rect 6772 62588 6836 62592
rect 6772 62532 6776 62588
rect 6776 62532 6832 62588
rect 6832 62532 6836 62588
rect 6772 62528 6836 62532
rect 6852 62588 6916 62592
rect 6852 62532 6856 62588
rect 6856 62532 6912 62588
rect 6912 62532 6916 62588
rect 6852 62528 6916 62532
rect 6932 62588 6996 62592
rect 6932 62532 6936 62588
rect 6936 62532 6992 62588
rect 6992 62532 6996 62588
rect 6932 62528 6996 62532
rect 87836 62588 87900 62592
rect 87836 62532 87840 62588
rect 87840 62532 87896 62588
rect 87896 62532 87900 62588
rect 87836 62528 87900 62532
rect 87916 62588 87980 62592
rect 87916 62532 87920 62588
rect 87920 62532 87976 62588
rect 87976 62532 87980 62588
rect 87916 62528 87980 62532
rect 87996 62588 88060 62592
rect 87996 62532 88000 62588
rect 88000 62532 88056 62588
rect 88056 62532 88060 62588
rect 87996 62528 88060 62532
rect 88076 62588 88140 62592
rect 88076 62532 88080 62588
rect 88080 62532 88136 62588
rect 88136 62532 88140 62588
rect 88076 62528 88140 62532
rect 5956 62044 6020 62048
rect 5956 61988 5960 62044
rect 5960 61988 6016 62044
rect 6016 61988 6020 62044
rect 5956 61984 6020 61988
rect 6036 62044 6100 62048
rect 6036 61988 6040 62044
rect 6040 61988 6096 62044
rect 6096 61988 6100 62044
rect 6036 61984 6100 61988
rect 6116 62044 6180 62048
rect 6116 61988 6120 62044
rect 6120 61988 6176 62044
rect 6176 61988 6180 62044
rect 6116 61984 6180 61988
rect 6196 62044 6260 62048
rect 6196 61988 6200 62044
rect 6200 61988 6256 62044
rect 6256 61988 6260 62044
rect 6196 61984 6260 61988
rect 87100 62044 87164 62048
rect 87100 61988 87104 62044
rect 87104 61988 87160 62044
rect 87160 61988 87164 62044
rect 87100 61984 87164 61988
rect 87180 62044 87244 62048
rect 87180 61988 87184 62044
rect 87184 61988 87240 62044
rect 87240 61988 87244 62044
rect 87180 61984 87244 61988
rect 87260 62044 87324 62048
rect 87260 61988 87264 62044
rect 87264 61988 87320 62044
rect 87320 61988 87324 62044
rect 87260 61984 87324 61988
rect 87340 62044 87404 62048
rect 87340 61988 87344 62044
rect 87344 61988 87400 62044
rect 87400 61988 87404 62044
rect 87340 61984 87404 61988
rect 6692 61500 6756 61504
rect 6692 61444 6696 61500
rect 6696 61444 6752 61500
rect 6752 61444 6756 61500
rect 6692 61440 6756 61444
rect 6772 61500 6836 61504
rect 6772 61444 6776 61500
rect 6776 61444 6832 61500
rect 6832 61444 6836 61500
rect 6772 61440 6836 61444
rect 6852 61500 6916 61504
rect 6852 61444 6856 61500
rect 6856 61444 6912 61500
rect 6912 61444 6916 61500
rect 6852 61440 6916 61444
rect 6932 61500 6996 61504
rect 6932 61444 6936 61500
rect 6936 61444 6992 61500
rect 6992 61444 6996 61500
rect 6932 61440 6996 61444
rect 87836 61500 87900 61504
rect 87836 61444 87840 61500
rect 87840 61444 87896 61500
rect 87896 61444 87900 61500
rect 87836 61440 87900 61444
rect 87916 61500 87980 61504
rect 87916 61444 87920 61500
rect 87920 61444 87976 61500
rect 87976 61444 87980 61500
rect 87916 61440 87980 61444
rect 87996 61500 88060 61504
rect 87996 61444 88000 61500
rect 88000 61444 88056 61500
rect 88056 61444 88060 61500
rect 87996 61440 88060 61444
rect 88076 61500 88140 61504
rect 88076 61444 88080 61500
rect 88080 61444 88136 61500
rect 88136 61444 88140 61500
rect 88076 61440 88140 61444
rect 5956 60956 6020 60960
rect 5956 60900 5960 60956
rect 5960 60900 6016 60956
rect 6016 60900 6020 60956
rect 5956 60896 6020 60900
rect 6036 60956 6100 60960
rect 6036 60900 6040 60956
rect 6040 60900 6096 60956
rect 6096 60900 6100 60956
rect 6036 60896 6100 60900
rect 6116 60956 6180 60960
rect 6116 60900 6120 60956
rect 6120 60900 6176 60956
rect 6176 60900 6180 60956
rect 6116 60896 6180 60900
rect 6196 60956 6260 60960
rect 6196 60900 6200 60956
rect 6200 60900 6256 60956
rect 6256 60900 6260 60956
rect 6196 60896 6260 60900
rect 87100 60956 87164 60960
rect 87100 60900 87104 60956
rect 87104 60900 87160 60956
rect 87160 60900 87164 60956
rect 87100 60896 87164 60900
rect 87180 60956 87244 60960
rect 87180 60900 87184 60956
rect 87184 60900 87240 60956
rect 87240 60900 87244 60956
rect 87180 60896 87244 60900
rect 87260 60956 87324 60960
rect 87260 60900 87264 60956
rect 87264 60900 87320 60956
rect 87320 60900 87324 60956
rect 87260 60896 87324 60900
rect 87340 60956 87404 60960
rect 87340 60900 87344 60956
rect 87344 60900 87400 60956
rect 87400 60900 87404 60956
rect 87340 60896 87404 60900
rect 6692 60412 6756 60416
rect 6692 60356 6696 60412
rect 6696 60356 6752 60412
rect 6752 60356 6756 60412
rect 6692 60352 6756 60356
rect 6772 60412 6836 60416
rect 6772 60356 6776 60412
rect 6776 60356 6832 60412
rect 6832 60356 6836 60412
rect 6772 60352 6836 60356
rect 6852 60412 6916 60416
rect 6852 60356 6856 60412
rect 6856 60356 6912 60412
rect 6912 60356 6916 60412
rect 6852 60352 6916 60356
rect 6932 60412 6996 60416
rect 6932 60356 6936 60412
rect 6936 60356 6992 60412
rect 6992 60356 6996 60412
rect 6932 60352 6996 60356
rect 87836 60412 87900 60416
rect 87836 60356 87840 60412
rect 87840 60356 87896 60412
rect 87896 60356 87900 60412
rect 87836 60352 87900 60356
rect 87916 60412 87980 60416
rect 87916 60356 87920 60412
rect 87920 60356 87976 60412
rect 87976 60356 87980 60412
rect 87916 60352 87980 60356
rect 87996 60412 88060 60416
rect 87996 60356 88000 60412
rect 88000 60356 88056 60412
rect 88056 60356 88060 60412
rect 87996 60352 88060 60356
rect 88076 60412 88140 60416
rect 88076 60356 88080 60412
rect 88080 60356 88136 60412
rect 88136 60356 88140 60412
rect 88076 60352 88140 60356
rect 5956 59868 6020 59872
rect 5956 59812 5960 59868
rect 5960 59812 6016 59868
rect 6016 59812 6020 59868
rect 5956 59808 6020 59812
rect 6036 59868 6100 59872
rect 6036 59812 6040 59868
rect 6040 59812 6096 59868
rect 6096 59812 6100 59868
rect 6036 59808 6100 59812
rect 6116 59868 6180 59872
rect 6116 59812 6120 59868
rect 6120 59812 6176 59868
rect 6176 59812 6180 59868
rect 6116 59808 6180 59812
rect 6196 59868 6260 59872
rect 6196 59812 6200 59868
rect 6200 59812 6256 59868
rect 6256 59812 6260 59868
rect 6196 59808 6260 59812
rect 87100 59868 87164 59872
rect 87100 59812 87104 59868
rect 87104 59812 87160 59868
rect 87160 59812 87164 59868
rect 87100 59808 87164 59812
rect 87180 59868 87244 59872
rect 87180 59812 87184 59868
rect 87184 59812 87240 59868
rect 87240 59812 87244 59868
rect 87180 59808 87244 59812
rect 87260 59868 87324 59872
rect 87260 59812 87264 59868
rect 87264 59812 87320 59868
rect 87320 59812 87324 59868
rect 87260 59808 87324 59812
rect 87340 59868 87404 59872
rect 87340 59812 87344 59868
rect 87344 59812 87400 59868
rect 87400 59812 87404 59868
rect 87340 59808 87404 59812
rect 6692 59324 6756 59328
rect 6692 59268 6696 59324
rect 6696 59268 6752 59324
rect 6752 59268 6756 59324
rect 6692 59264 6756 59268
rect 6772 59324 6836 59328
rect 6772 59268 6776 59324
rect 6776 59268 6832 59324
rect 6832 59268 6836 59324
rect 6772 59264 6836 59268
rect 6852 59324 6916 59328
rect 6852 59268 6856 59324
rect 6856 59268 6912 59324
rect 6912 59268 6916 59324
rect 6852 59264 6916 59268
rect 6932 59324 6996 59328
rect 6932 59268 6936 59324
rect 6936 59268 6992 59324
rect 6992 59268 6996 59324
rect 6932 59264 6996 59268
rect 87836 59324 87900 59328
rect 87836 59268 87840 59324
rect 87840 59268 87896 59324
rect 87896 59268 87900 59324
rect 87836 59264 87900 59268
rect 87916 59324 87980 59328
rect 87916 59268 87920 59324
rect 87920 59268 87976 59324
rect 87976 59268 87980 59324
rect 87916 59264 87980 59268
rect 87996 59324 88060 59328
rect 87996 59268 88000 59324
rect 88000 59268 88056 59324
rect 88056 59268 88060 59324
rect 87996 59264 88060 59268
rect 88076 59324 88140 59328
rect 88076 59268 88080 59324
rect 88080 59268 88136 59324
rect 88136 59268 88140 59324
rect 88076 59264 88140 59268
rect 5956 58780 6020 58784
rect 5956 58724 5960 58780
rect 5960 58724 6016 58780
rect 6016 58724 6020 58780
rect 5956 58720 6020 58724
rect 6036 58780 6100 58784
rect 6036 58724 6040 58780
rect 6040 58724 6096 58780
rect 6096 58724 6100 58780
rect 6036 58720 6100 58724
rect 6116 58780 6180 58784
rect 6116 58724 6120 58780
rect 6120 58724 6176 58780
rect 6176 58724 6180 58780
rect 6116 58720 6180 58724
rect 6196 58780 6260 58784
rect 6196 58724 6200 58780
rect 6200 58724 6256 58780
rect 6256 58724 6260 58780
rect 6196 58720 6260 58724
rect 87100 58780 87164 58784
rect 87100 58724 87104 58780
rect 87104 58724 87160 58780
rect 87160 58724 87164 58780
rect 87100 58720 87164 58724
rect 87180 58780 87244 58784
rect 87180 58724 87184 58780
rect 87184 58724 87240 58780
rect 87240 58724 87244 58780
rect 87180 58720 87244 58724
rect 87260 58780 87324 58784
rect 87260 58724 87264 58780
rect 87264 58724 87320 58780
rect 87320 58724 87324 58780
rect 87260 58720 87324 58724
rect 87340 58780 87404 58784
rect 87340 58724 87344 58780
rect 87344 58724 87400 58780
rect 87400 58724 87404 58780
rect 87340 58720 87404 58724
rect 6692 58236 6756 58240
rect 6692 58180 6696 58236
rect 6696 58180 6752 58236
rect 6752 58180 6756 58236
rect 6692 58176 6756 58180
rect 6772 58236 6836 58240
rect 6772 58180 6776 58236
rect 6776 58180 6832 58236
rect 6832 58180 6836 58236
rect 6772 58176 6836 58180
rect 6852 58236 6916 58240
rect 6852 58180 6856 58236
rect 6856 58180 6912 58236
rect 6912 58180 6916 58236
rect 6852 58176 6916 58180
rect 6932 58236 6996 58240
rect 6932 58180 6936 58236
rect 6936 58180 6992 58236
rect 6992 58180 6996 58236
rect 6932 58176 6996 58180
rect 87836 58236 87900 58240
rect 87836 58180 87840 58236
rect 87840 58180 87896 58236
rect 87896 58180 87900 58236
rect 87836 58176 87900 58180
rect 87916 58236 87980 58240
rect 87916 58180 87920 58236
rect 87920 58180 87976 58236
rect 87976 58180 87980 58236
rect 87916 58176 87980 58180
rect 87996 58236 88060 58240
rect 87996 58180 88000 58236
rect 88000 58180 88056 58236
rect 88056 58180 88060 58236
rect 87996 58176 88060 58180
rect 88076 58236 88140 58240
rect 88076 58180 88080 58236
rect 88080 58180 88136 58236
rect 88136 58180 88140 58236
rect 88076 58176 88140 58180
rect 5956 57692 6020 57696
rect 5956 57636 5960 57692
rect 5960 57636 6016 57692
rect 6016 57636 6020 57692
rect 5956 57632 6020 57636
rect 6036 57692 6100 57696
rect 6036 57636 6040 57692
rect 6040 57636 6096 57692
rect 6096 57636 6100 57692
rect 6036 57632 6100 57636
rect 6116 57692 6180 57696
rect 6116 57636 6120 57692
rect 6120 57636 6176 57692
rect 6176 57636 6180 57692
rect 6116 57632 6180 57636
rect 6196 57692 6260 57696
rect 6196 57636 6200 57692
rect 6200 57636 6256 57692
rect 6256 57636 6260 57692
rect 6196 57632 6260 57636
rect 87100 57692 87164 57696
rect 87100 57636 87104 57692
rect 87104 57636 87160 57692
rect 87160 57636 87164 57692
rect 87100 57632 87164 57636
rect 87180 57692 87244 57696
rect 87180 57636 87184 57692
rect 87184 57636 87240 57692
rect 87240 57636 87244 57692
rect 87180 57632 87244 57636
rect 87260 57692 87324 57696
rect 87260 57636 87264 57692
rect 87264 57636 87320 57692
rect 87320 57636 87324 57692
rect 87260 57632 87324 57636
rect 87340 57692 87404 57696
rect 87340 57636 87344 57692
rect 87344 57636 87400 57692
rect 87400 57636 87404 57692
rect 87340 57632 87404 57636
rect 6692 57148 6756 57152
rect 6692 57092 6696 57148
rect 6696 57092 6752 57148
rect 6752 57092 6756 57148
rect 6692 57088 6756 57092
rect 6772 57148 6836 57152
rect 6772 57092 6776 57148
rect 6776 57092 6832 57148
rect 6832 57092 6836 57148
rect 6772 57088 6836 57092
rect 6852 57148 6916 57152
rect 6852 57092 6856 57148
rect 6856 57092 6912 57148
rect 6912 57092 6916 57148
rect 6852 57088 6916 57092
rect 6932 57148 6996 57152
rect 6932 57092 6936 57148
rect 6936 57092 6992 57148
rect 6992 57092 6996 57148
rect 6932 57088 6996 57092
rect 87836 57148 87900 57152
rect 87836 57092 87840 57148
rect 87840 57092 87896 57148
rect 87896 57092 87900 57148
rect 87836 57088 87900 57092
rect 87916 57148 87980 57152
rect 87916 57092 87920 57148
rect 87920 57092 87976 57148
rect 87976 57092 87980 57148
rect 87916 57088 87980 57092
rect 87996 57148 88060 57152
rect 87996 57092 88000 57148
rect 88000 57092 88056 57148
rect 88056 57092 88060 57148
rect 87996 57088 88060 57092
rect 88076 57148 88140 57152
rect 88076 57092 88080 57148
rect 88080 57092 88136 57148
rect 88136 57092 88140 57148
rect 88076 57088 88140 57092
rect 5956 56604 6020 56608
rect 5956 56548 5960 56604
rect 5960 56548 6016 56604
rect 6016 56548 6020 56604
rect 5956 56544 6020 56548
rect 6036 56604 6100 56608
rect 6036 56548 6040 56604
rect 6040 56548 6096 56604
rect 6096 56548 6100 56604
rect 6036 56544 6100 56548
rect 6116 56604 6180 56608
rect 6116 56548 6120 56604
rect 6120 56548 6176 56604
rect 6176 56548 6180 56604
rect 6116 56544 6180 56548
rect 6196 56604 6260 56608
rect 6196 56548 6200 56604
rect 6200 56548 6256 56604
rect 6256 56548 6260 56604
rect 6196 56544 6260 56548
rect 87100 56604 87164 56608
rect 87100 56548 87104 56604
rect 87104 56548 87160 56604
rect 87160 56548 87164 56604
rect 87100 56544 87164 56548
rect 87180 56604 87244 56608
rect 87180 56548 87184 56604
rect 87184 56548 87240 56604
rect 87240 56548 87244 56604
rect 87180 56544 87244 56548
rect 87260 56604 87324 56608
rect 87260 56548 87264 56604
rect 87264 56548 87320 56604
rect 87320 56548 87324 56604
rect 87260 56544 87324 56548
rect 87340 56604 87404 56608
rect 87340 56548 87344 56604
rect 87344 56548 87400 56604
rect 87400 56548 87404 56604
rect 87340 56544 87404 56548
rect 6692 56060 6756 56064
rect 6692 56004 6696 56060
rect 6696 56004 6752 56060
rect 6752 56004 6756 56060
rect 6692 56000 6756 56004
rect 6772 56060 6836 56064
rect 6772 56004 6776 56060
rect 6776 56004 6832 56060
rect 6832 56004 6836 56060
rect 6772 56000 6836 56004
rect 6852 56060 6916 56064
rect 6852 56004 6856 56060
rect 6856 56004 6912 56060
rect 6912 56004 6916 56060
rect 6852 56000 6916 56004
rect 6932 56060 6996 56064
rect 6932 56004 6936 56060
rect 6936 56004 6992 56060
rect 6992 56004 6996 56060
rect 6932 56000 6996 56004
rect 87836 56060 87900 56064
rect 87836 56004 87840 56060
rect 87840 56004 87896 56060
rect 87896 56004 87900 56060
rect 87836 56000 87900 56004
rect 87916 56060 87980 56064
rect 87916 56004 87920 56060
rect 87920 56004 87976 56060
rect 87976 56004 87980 56060
rect 87916 56000 87980 56004
rect 87996 56060 88060 56064
rect 87996 56004 88000 56060
rect 88000 56004 88056 56060
rect 88056 56004 88060 56060
rect 87996 56000 88060 56004
rect 88076 56060 88140 56064
rect 88076 56004 88080 56060
rect 88080 56004 88136 56060
rect 88136 56004 88140 56060
rect 88076 56000 88140 56004
rect 5956 55516 6020 55520
rect 5956 55460 5960 55516
rect 5960 55460 6016 55516
rect 6016 55460 6020 55516
rect 5956 55456 6020 55460
rect 6036 55516 6100 55520
rect 6036 55460 6040 55516
rect 6040 55460 6096 55516
rect 6096 55460 6100 55516
rect 6036 55456 6100 55460
rect 6116 55516 6180 55520
rect 6116 55460 6120 55516
rect 6120 55460 6176 55516
rect 6176 55460 6180 55516
rect 6116 55456 6180 55460
rect 6196 55516 6260 55520
rect 6196 55460 6200 55516
rect 6200 55460 6256 55516
rect 6256 55460 6260 55516
rect 6196 55456 6260 55460
rect 87100 55516 87164 55520
rect 87100 55460 87104 55516
rect 87104 55460 87160 55516
rect 87160 55460 87164 55516
rect 87100 55456 87164 55460
rect 87180 55516 87244 55520
rect 87180 55460 87184 55516
rect 87184 55460 87240 55516
rect 87240 55460 87244 55516
rect 87180 55456 87244 55460
rect 87260 55516 87324 55520
rect 87260 55460 87264 55516
rect 87264 55460 87320 55516
rect 87320 55460 87324 55516
rect 87260 55456 87324 55460
rect 87340 55516 87404 55520
rect 87340 55460 87344 55516
rect 87344 55460 87400 55516
rect 87400 55460 87404 55516
rect 87340 55456 87404 55460
rect 6692 54972 6756 54976
rect 6692 54916 6696 54972
rect 6696 54916 6752 54972
rect 6752 54916 6756 54972
rect 6692 54912 6756 54916
rect 6772 54972 6836 54976
rect 6772 54916 6776 54972
rect 6776 54916 6832 54972
rect 6832 54916 6836 54972
rect 6772 54912 6836 54916
rect 6852 54972 6916 54976
rect 6852 54916 6856 54972
rect 6856 54916 6912 54972
rect 6912 54916 6916 54972
rect 6852 54912 6916 54916
rect 6932 54972 6996 54976
rect 6932 54916 6936 54972
rect 6936 54916 6992 54972
rect 6992 54916 6996 54972
rect 6932 54912 6996 54916
rect 87836 54972 87900 54976
rect 87836 54916 87840 54972
rect 87840 54916 87896 54972
rect 87896 54916 87900 54972
rect 87836 54912 87900 54916
rect 87916 54972 87980 54976
rect 87916 54916 87920 54972
rect 87920 54916 87976 54972
rect 87976 54916 87980 54972
rect 87916 54912 87980 54916
rect 87996 54972 88060 54976
rect 87996 54916 88000 54972
rect 88000 54916 88056 54972
rect 88056 54916 88060 54972
rect 87996 54912 88060 54916
rect 88076 54972 88140 54976
rect 88076 54916 88080 54972
rect 88080 54916 88136 54972
rect 88136 54916 88140 54972
rect 88076 54912 88140 54916
rect 5956 54428 6020 54432
rect 5956 54372 5960 54428
rect 5960 54372 6016 54428
rect 6016 54372 6020 54428
rect 5956 54368 6020 54372
rect 6036 54428 6100 54432
rect 6036 54372 6040 54428
rect 6040 54372 6096 54428
rect 6096 54372 6100 54428
rect 6036 54368 6100 54372
rect 6116 54428 6180 54432
rect 6116 54372 6120 54428
rect 6120 54372 6176 54428
rect 6176 54372 6180 54428
rect 6116 54368 6180 54372
rect 6196 54428 6260 54432
rect 6196 54372 6200 54428
rect 6200 54372 6256 54428
rect 6256 54372 6260 54428
rect 6196 54368 6260 54372
rect 87100 54428 87164 54432
rect 87100 54372 87104 54428
rect 87104 54372 87160 54428
rect 87160 54372 87164 54428
rect 87100 54368 87164 54372
rect 87180 54428 87244 54432
rect 87180 54372 87184 54428
rect 87184 54372 87240 54428
rect 87240 54372 87244 54428
rect 87180 54368 87244 54372
rect 87260 54428 87324 54432
rect 87260 54372 87264 54428
rect 87264 54372 87320 54428
rect 87320 54372 87324 54428
rect 87260 54368 87324 54372
rect 87340 54428 87404 54432
rect 87340 54372 87344 54428
rect 87344 54372 87400 54428
rect 87400 54372 87404 54428
rect 87340 54368 87404 54372
rect 6692 53884 6756 53888
rect 6692 53828 6696 53884
rect 6696 53828 6752 53884
rect 6752 53828 6756 53884
rect 6692 53824 6756 53828
rect 6772 53884 6836 53888
rect 6772 53828 6776 53884
rect 6776 53828 6832 53884
rect 6832 53828 6836 53884
rect 6772 53824 6836 53828
rect 6852 53884 6916 53888
rect 6852 53828 6856 53884
rect 6856 53828 6912 53884
rect 6912 53828 6916 53884
rect 6852 53824 6916 53828
rect 6932 53884 6996 53888
rect 6932 53828 6936 53884
rect 6936 53828 6992 53884
rect 6992 53828 6996 53884
rect 6932 53824 6996 53828
rect 87836 53884 87900 53888
rect 87836 53828 87840 53884
rect 87840 53828 87896 53884
rect 87896 53828 87900 53884
rect 87836 53824 87900 53828
rect 87916 53884 87980 53888
rect 87916 53828 87920 53884
rect 87920 53828 87976 53884
rect 87976 53828 87980 53884
rect 87916 53824 87980 53828
rect 87996 53884 88060 53888
rect 87996 53828 88000 53884
rect 88000 53828 88056 53884
rect 88056 53828 88060 53884
rect 87996 53824 88060 53828
rect 88076 53884 88140 53888
rect 88076 53828 88080 53884
rect 88080 53828 88136 53884
rect 88136 53828 88140 53884
rect 88076 53824 88140 53828
rect 5956 53340 6020 53344
rect 5956 53284 5960 53340
rect 5960 53284 6016 53340
rect 6016 53284 6020 53340
rect 5956 53280 6020 53284
rect 6036 53340 6100 53344
rect 6036 53284 6040 53340
rect 6040 53284 6096 53340
rect 6096 53284 6100 53340
rect 6036 53280 6100 53284
rect 6116 53340 6180 53344
rect 6116 53284 6120 53340
rect 6120 53284 6176 53340
rect 6176 53284 6180 53340
rect 6116 53280 6180 53284
rect 6196 53340 6260 53344
rect 6196 53284 6200 53340
rect 6200 53284 6256 53340
rect 6256 53284 6260 53340
rect 6196 53280 6260 53284
rect 87100 53340 87164 53344
rect 87100 53284 87104 53340
rect 87104 53284 87160 53340
rect 87160 53284 87164 53340
rect 87100 53280 87164 53284
rect 87180 53340 87244 53344
rect 87180 53284 87184 53340
rect 87184 53284 87240 53340
rect 87240 53284 87244 53340
rect 87180 53280 87244 53284
rect 87260 53340 87324 53344
rect 87260 53284 87264 53340
rect 87264 53284 87320 53340
rect 87320 53284 87324 53340
rect 87260 53280 87324 53284
rect 87340 53340 87404 53344
rect 87340 53284 87344 53340
rect 87344 53284 87400 53340
rect 87400 53284 87404 53340
rect 87340 53280 87404 53284
rect 6692 52796 6756 52800
rect 6692 52740 6696 52796
rect 6696 52740 6752 52796
rect 6752 52740 6756 52796
rect 6692 52736 6756 52740
rect 6772 52796 6836 52800
rect 6772 52740 6776 52796
rect 6776 52740 6832 52796
rect 6832 52740 6836 52796
rect 6772 52736 6836 52740
rect 6852 52796 6916 52800
rect 6852 52740 6856 52796
rect 6856 52740 6912 52796
rect 6912 52740 6916 52796
rect 6852 52736 6916 52740
rect 6932 52796 6996 52800
rect 6932 52740 6936 52796
rect 6936 52740 6992 52796
rect 6992 52740 6996 52796
rect 6932 52736 6996 52740
rect 87836 52796 87900 52800
rect 87836 52740 87840 52796
rect 87840 52740 87896 52796
rect 87896 52740 87900 52796
rect 87836 52736 87900 52740
rect 87916 52796 87980 52800
rect 87916 52740 87920 52796
rect 87920 52740 87976 52796
rect 87976 52740 87980 52796
rect 87916 52736 87980 52740
rect 87996 52796 88060 52800
rect 87996 52740 88000 52796
rect 88000 52740 88056 52796
rect 88056 52740 88060 52796
rect 87996 52736 88060 52740
rect 88076 52796 88140 52800
rect 88076 52740 88080 52796
rect 88080 52740 88136 52796
rect 88136 52740 88140 52796
rect 88076 52736 88140 52740
rect 5956 52252 6020 52256
rect 5956 52196 5960 52252
rect 5960 52196 6016 52252
rect 6016 52196 6020 52252
rect 5956 52192 6020 52196
rect 6036 52252 6100 52256
rect 6036 52196 6040 52252
rect 6040 52196 6096 52252
rect 6096 52196 6100 52252
rect 6036 52192 6100 52196
rect 6116 52252 6180 52256
rect 6116 52196 6120 52252
rect 6120 52196 6176 52252
rect 6176 52196 6180 52252
rect 6116 52192 6180 52196
rect 6196 52252 6260 52256
rect 6196 52196 6200 52252
rect 6200 52196 6256 52252
rect 6256 52196 6260 52252
rect 6196 52192 6260 52196
rect 87100 52252 87164 52256
rect 87100 52196 87104 52252
rect 87104 52196 87160 52252
rect 87160 52196 87164 52252
rect 87100 52192 87164 52196
rect 87180 52252 87244 52256
rect 87180 52196 87184 52252
rect 87184 52196 87240 52252
rect 87240 52196 87244 52252
rect 87180 52192 87244 52196
rect 87260 52252 87324 52256
rect 87260 52196 87264 52252
rect 87264 52196 87320 52252
rect 87320 52196 87324 52252
rect 87260 52192 87324 52196
rect 87340 52252 87404 52256
rect 87340 52196 87344 52252
rect 87344 52196 87400 52252
rect 87400 52196 87404 52252
rect 87340 52192 87404 52196
rect 6692 51708 6756 51712
rect 6692 51652 6696 51708
rect 6696 51652 6752 51708
rect 6752 51652 6756 51708
rect 6692 51648 6756 51652
rect 6772 51708 6836 51712
rect 6772 51652 6776 51708
rect 6776 51652 6832 51708
rect 6832 51652 6836 51708
rect 6772 51648 6836 51652
rect 6852 51708 6916 51712
rect 6852 51652 6856 51708
rect 6856 51652 6912 51708
rect 6912 51652 6916 51708
rect 6852 51648 6916 51652
rect 6932 51708 6996 51712
rect 6932 51652 6936 51708
rect 6936 51652 6992 51708
rect 6992 51652 6996 51708
rect 6932 51648 6996 51652
rect 87836 51708 87900 51712
rect 87836 51652 87840 51708
rect 87840 51652 87896 51708
rect 87896 51652 87900 51708
rect 87836 51648 87900 51652
rect 87916 51708 87980 51712
rect 87916 51652 87920 51708
rect 87920 51652 87976 51708
rect 87976 51652 87980 51708
rect 87916 51648 87980 51652
rect 87996 51708 88060 51712
rect 87996 51652 88000 51708
rect 88000 51652 88056 51708
rect 88056 51652 88060 51708
rect 87996 51648 88060 51652
rect 88076 51708 88140 51712
rect 88076 51652 88080 51708
rect 88080 51652 88136 51708
rect 88136 51652 88140 51708
rect 88076 51648 88140 51652
rect 5956 51164 6020 51168
rect 5956 51108 5960 51164
rect 5960 51108 6016 51164
rect 6016 51108 6020 51164
rect 5956 51104 6020 51108
rect 6036 51164 6100 51168
rect 6036 51108 6040 51164
rect 6040 51108 6096 51164
rect 6096 51108 6100 51164
rect 6036 51104 6100 51108
rect 6116 51164 6180 51168
rect 6116 51108 6120 51164
rect 6120 51108 6176 51164
rect 6176 51108 6180 51164
rect 6116 51104 6180 51108
rect 6196 51164 6260 51168
rect 6196 51108 6200 51164
rect 6200 51108 6256 51164
rect 6256 51108 6260 51164
rect 6196 51104 6260 51108
rect 87100 51164 87164 51168
rect 87100 51108 87104 51164
rect 87104 51108 87160 51164
rect 87160 51108 87164 51164
rect 87100 51104 87164 51108
rect 87180 51164 87244 51168
rect 87180 51108 87184 51164
rect 87184 51108 87240 51164
rect 87240 51108 87244 51164
rect 87180 51104 87244 51108
rect 87260 51164 87324 51168
rect 87260 51108 87264 51164
rect 87264 51108 87320 51164
rect 87320 51108 87324 51164
rect 87260 51104 87324 51108
rect 87340 51164 87404 51168
rect 87340 51108 87344 51164
rect 87344 51108 87400 51164
rect 87400 51108 87404 51164
rect 87340 51104 87404 51108
rect 6692 50620 6756 50624
rect 6692 50564 6696 50620
rect 6696 50564 6752 50620
rect 6752 50564 6756 50620
rect 6692 50560 6756 50564
rect 6772 50620 6836 50624
rect 6772 50564 6776 50620
rect 6776 50564 6832 50620
rect 6832 50564 6836 50620
rect 6772 50560 6836 50564
rect 6852 50620 6916 50624
rect 6852 50564 6856 50620
rect 6856 50564 6912 50620
rect 6912 50564 6916 50620
rect 6852 50560 6916 50564
rect 6932 50620 6996 50624
rect 6932 50564 6936 50620
rect 6936 50564 6992 50620
rect 6992 50564 6996 50620
rect 6932 50560 6996 50564
rect 87836 50620 87900 50624
rect 87836 50564 87840 50620
rect 87840 50564 87896 50620
rect 87896 50564 87900 50620
rect 87836 50560 87900 50564
rect 87916 50620 87980 50624
rect 87916 50564 87920 50620
rect 87920 50564 87976 50620
rect 87976 50564 87980 50620
rect 87916 50560 87980 50564
rect 87996 50620 88060 50624
rect 87996 50564 88000 50620
rect 88000 50564 88056 50620
rect 88056 50564 88060 50620
rect 87996 50560 88060 50564
rect 88076 50620 88140 50624
rect 88076 50564 88080 50620
rect 88080 50564 88136 50620
rect 88136 50564 88140 50620
rect 88076 50560 88140 50564
rect 5956 50076 6020 50080
rect 5956 50020 5960 50076
rect 5960 50020 6016 50076
rect 6016 50020 6020 50076
rect 5956 50016 6020 50020
rect 6036 50076 6100 50080
rect 6036 50020 6040 50076
rect 6040 50020 6096 50076
rect 6096 50020 6100 50076
rect 6036 50016 6100 50020
rect 6116 50076 6180 50080
rect 6116 50020 6120 50076
rect 6120 50020 6176 50076
rect 6176 50020 6180 50076
rect 6116 50016 6180 50020
rect 6196 50076 6260 50080
rect 6196 50020 6200 50076
rect 6200 50020 6256 50076
rect 6256 50020 6260 50076
rect 6196 50016 6260 50020
rect 87100 50076 87164 50080
rect 87100 50020 87104 50076
rect 87104 50020 87160 50076
rect 87160 50020 87164 50076
rect 87100 50016 87164 50020
rect 87180 50076 87244 50080
rect 87180 50020 87184 50076
rect 87184 50020 87240 50076
rect 87240 50020 87244 50076
rect 87180 50016 87244 50020
rect 87260 50076 87324 50080
rect 87260 50020 87264 50076
rect 87264 50020 87320 50076
rect 87320 50020 87324 50076
rect 87260 50016 87324 50020
rect 87340 50076 87404 50080
rect 87340 50020 87344 50076
rect 87344 50020 87400 50076
rect 87400 50020 87404 50076
rect 87340 50016 87404 50020
rect 6692 49532 6756 49536
rect 6692 49476 6696 49532
rect 6696 49476 6752 49532
rect 6752 49476 6756 49532
rect 6692 49472 6756 49476
rect 6772 49532 6836 49536
rect 6772 49476 6776 49532
rect 6776 49476 6832 49532
rect 6832 49476 6836 49532
rect 6772 49472 6836 49476
rect 6852 49532 6916 49536
rect 6852 49476 6856 49532
rect 6856 49476 6912 49532
rect 6912 49476 6916 49532
rect 6852 49472 6916 49476
rect 6932 49532 6996 49536
rect 6932 49476 6936 49532
rect 6936 49476 6992 49532
rect 6992 49476 6996 49532
rect 6932 49472 6996 49476
rect 87836 49532 87900 49536
rect 87836 49476 87840 49532
rect 87840 49476 87896 49532
rect 87896 49476 87900 49532
rect 87836 49472 87900 49476
rect 87916 49532 87980 49536
rect 87916 49476 87920 49532
rect 87920 49476 87976 49532
rect 87976 49476 87980 49532
rect 87916 49472 87980 49476
rect 87996 49532 88060 49536
rect 87996 49476 88000 49532
rect 88000 49476 88056 49532
rect 88056 49476 88060 49532
rect 87996 49472 88060 49476
rect 88076 49532 88140 49536
rect 88076 49476 88080 49532
rect 88080 49476 88136 49532
rect 88136 49476 88140 49532
rect 88076 49472 88140 49476
rect 5956 48988 6020 48992
rect 5956 48932 5960 48988
rect 5960 48932 6016 48988
rect 6016 48932 6020 48988
rect 5956 48928 6020 48932
rect 6036 48988 6100 48992
rect 6036 48932 6040 48988
rect 6040 48932 6096 48988
rect 6096 48932 6100 48988
rect 6036 48928 6100 48932
rect 6116 48988 6180 48992
rect 6116 48932 6120 48988
rect 6120 48932 6176 48988
rect 6176 48932 6180 48988
rect 6116 48928 6180 48932
rect 6196 48988 6260 48992
rect 6196 48932 6200 48988
rect 6200 48932 6256 48988
rect 6256 48932 6260 48988
rect 6196 48928 6260 48932
rect 87100 48988 87164 48992
rect 87100 48932 87104 48988
rect 87104 48932 87160 48988
rect 87160 48932 87164 48988
rect 87100 48928 87164 48932
rect 87180 48988 87244 48992
rect 87180 48932 87184 48988
rect 87184 48932 87240 48988
rect 87240 48932 87244 48988
rect 87180 48928 87244 48932
rect 87260 48988 87324 48992
rect 87260 48932 87264 48988
rect 87264 48932 87320 48988
rect 87320 48932 87324 48988
rect 87260 48928 87324 48932
rect 87340 48988 87404 48992
rect 87340 48932 87344 48988
rect 87344 48932 87400 48988
rect 87400 48932 87404 48988
rect 87340 48928 87404 48932
rect 6692 48444 6756 48448
rect 6692 48388 6696 48444
rect 6696 48388 6752 48444
rect 6752 48388 6756 48444
rect 6692 48384 6756 48388
rect 6772 48444 6836 48448
rect 6772 48388 6776 48444
rect 6776 48388 6832 48444
rect 6832 48388 6836 48444
rect 6772 48384 6836 48388
rect 6852 48444 6916 48448
rect 6852 48388 6856 48444
rect 6856 48388 6912 48444
rect 6912 48388 6916 48444
rect 6852 48384 6916 48388
rect 6932 48444 6996 48448
rect 6932 48388 6936 48444
rect 6936 48388 6992 48444
rect 6992 48388 6996 48444
rect 6932 48384 6996 48388
rect 87836 48444 87900 48448
rect 87836 48388 87840 48444
rect 87840 48388 87896 48444
rect 87896 48388 87900 48444
rect 87836 48384 87900 48388
rect 87916 48444 87980 48448
rect 87916 48388 87920 48444
rect 87920 48388 87976 48444
rect 87976 48388 87980 48444
rect 87916 48384 87980 48388
rect 87996 48444 88060 48448
rect 87996 48388 88000 48444
rect 88000 48388 88056 48444
rect 88056 48388 88060 48444
rect 87996 48384 88060 48388
rect 88076 48444 88140 48448
rect 88076 48388 88080 48444
rect 88080 48388 88136 48444
rect 88136 48388 88140 48444
rect 88076 48384 88140 48388
rect 5956 47900 6020 47904
rect 5956 47844 5960 47900
rect 5960 47844 6016 47900
rect 6016 47844 6020 47900
rect 5956 47840 6020 47844
rect 6036 47900 6100 47904
rect 6036 47844 6040 47900
rect 6040 47844 6096 47900
rect 6096 47844 6100 47900
rect 6036 47840 6100 47844
rect 6116 47900 6180 47904
rect 6116 47844 6120 47900
rect 6120 47844 6176 47900
rect 6176 47844 6180 47900
rect 6116 47840 6180 47844
rect 6196 47900 6260 47904
rect 6196 47844 6200 47900
rect 6200 47844 6256 47900
rect 6256 47844 6260 47900
rect 6196 47840 6260 47844
rect 87100 47900 87164 47904
rect 87100 47844 87104 47900
rect 87104 47844 87160 47900
rect 87160 47844 87164 47900
rect 87100 47840 87164 47844
rect 87180 47900 87244 47904
rect 87180 47844 87184 47900
rect 87184 47844 87240 47900
rect 87240 47844 87244 47900
rect 87180 47840 87244 47844
rect 87260 47900 87324 47904
rect 87260 47844 87264 47900
rect 87264 47844 87320 47900
rect 87320 47844 87324 47900
rect 87260 47840 87324 47844
rect 87340 47900 87404 47904
rect 87340 47844 87344 47900
rect 87344 47844 87400 47900
rect 87400 47844 87404 47900
rect 87340 47840 87404 47844
rect 6692 47356 6756 47360
rect 6692 47300 6696 47356
rect 6696 47300 6752 47356
rect 6752 47300 6756 47356
rect 6692 47296 6756 47300
rect 6772 47356 6836 47360
rect 6772 47300 6776 47356
rect 6776 47300 6832 47356
rect 6832 47300 6836 47356
rect 6772 47296 6836 47300
rect 6852 47356 6916 47360
rect 6852 47300 6856 47356
rect 6856 47300 6912 47356
rect 6912 47300 6916 47356
rect 6852 47296 6916 47300
rect 6932 47356 6996 47360
rect 6932 47300 6936 47356
rect 6936 47300 6992 47356
rect 6992 47300 6996 47356
rect 6932 47296 6996 47300
rect 87836 47356 87900 47360
rect 87836 47300 87840 47356
rect 87840 47300 87896 47356
rect 87896 47300 87900 47356
rect 87836 47296 87900 47300
rect 87916 47356 87980 47360
rect 87916 47300 87920 47356
rect 87920 47300 87976 47356
rect 87976 47300 87980 47356
rect 87916 47296 87980 47300
rect 87996 47356 88060 47360
rect 87996 47300 88000 47356
rect 88000 47300 88056 47356
rect 88056 47300 88060 47356
rect 87996 47296 88060 47300
rect 88076 47356 88140 47360
rect 88076 47300 88080 47356
rect 88080 47300 88136 47356
rect 88136 47300 88140 47356
rect 88076 47296 88140 47300
rect 5956 46812 6020 46816
rect 5956 46756 5960 46812
rect 5960 46756 6016 46812
rect 6016 46756 6020 46812
rect 5956 46752 6020 46756
rect 6036 46812 6100 46816
rect 6036 46756 6040 46812
rect 6040 46756 6096 46812
rect 6096 46756 6100 46812
rect 6036 46752 6100 46756
rect 6116 46812 6180 46816
rect 6116 46756 6120 46812
rect 6120 46756 6176 46812
rect 6176 46756 6180 46812
rect 6116 46752 6180 46756
rect 6196 46812 6260 46816
rect 6196 46756 6200 46812
rect 6200 46756 6256 46812
rect 6256 46756 6260 46812
rect 6196 46752 6260 46756
rect 87100 46812 87164 46816
rect 87100 46756 87104 46812
rect 87104 46756 87160 46812
rect 87160 46756 87164 46812
rect 87100 46752 87164 46756
rect 87180 46812 87244 46816
rect 87180 46756 87184 46812
rect 87184 46756 87240 46812
rect 87240 46756 87244 46812
rect 87180 46752 87244 46756
rect 87260 46812 87324 46816
rect 87260 46756 87264 46812
rect 87264 46756 87320 46812
rect 87320 46756 87324 46812
rect 87260 46752 87324 46756
rect 87340 46812 87404 46816
rect 87340 46756 87344 46812
rect 87344 46756 87400 46812
rect 87400 46756 87404 46812
rect 87340 46752 87404 46756
rect 6692 46268 6756 46272
rect 6692 46212 6696 46268
rect 6696 46212 6752 46268
rect 6752 46212 6756 46268
rect 6692 46208 6756 46212
rect 6772 46268 6836 46272
rect 6772 46212 6776 46268
rect 6776 46212 6832 46268
rect 6832 46212 6836 46268
rect 6772 46208 6836 46212
rect 6852 46268 6916 46272
rect 6852 46212 6856 46268
rect 6856 46212 6912 46268
rect 6912 46212 6916 46268
rect 6852 46208 6916 46212
rect 6932 46268 6996 46272
rect 6932 46212 6936 46268
rect 6936 46212 6992 46268
rect 6992 46212 6996 46268
rect 6932 46208 6996 46212
rect 87836 46268 87900 46272
rect 87836 46212 87840 46268
rect 87840 46212 87896 46268
rect 87896 46212 87900 46268
rect 87836 46208 87900 46212
rect 87916 46268 87980 46272
rect 87916 46212 87920 46268
rect 87920 46212 87976 46268
rect 87976 46212 87980 46268
rect 87916 46208 87980 46212
rect 87996 46268 88060 46272
rect 87996 46212 88000 46268
rect 88000 46212 88056 46268
rect 88056 46212 88060 46268
rect 87996 46208 88060 46212
rect 88076 46268 88140 46272
rect 88076 46212 88080 46268
rect 88080 46212 88136 46268
rect 88136 46212 88140 46268
rect 88076 46208 88140 46212
rect 5956 45724 6020 45728
rect 5956 45668 5960 45724
rect 5960 45668 6016 45724
rect 6016 45668 6020 45724
rect 5956 45664 6020 45668
rect 6036 45724 6100 45728
rect 6036 45668 6040 45724
rect 6040 45668 6096 45724
rect 6096 45668 6100 45724
rect 6036 45664 6100 45668
rect 6116 45724 6180 45728
rect 6116 45668 6120 45724
rect 6120 45668 6176 45724
rect 6176 45668 6180 45724
rect 6116 45664 6180 45668
rect 6196 45724 6260 45728
rect 6196 45668 6200 45724
rect 6200 45668 6256 45724
rect 6256 45668 6260 45724
rect 6196 45664 6260 45668
rect 87100 45724 87164 45728
rect 87100 45668 87104 45724
rect 87104 45668 87160 45724
rect 87160 45668 87164 45724
rect 87100 45664 87164 45668
rect 87180 45724 87244 45728
rect 87180 45668 87184 45724
rect 87184 45668 87240 45724
rect 87240 45668 87244 45724
rect 87180 45664 87244 45668
rect 87260 45724 87324 45728
rect 87260 45668 87264 45724
rect 87264 45668 87320 45724
rect 87320 45668 87324 45724
rect 87260 45664 87324 45668
rect 87340 45724 87404 45728
rect 87340 45668 87344 45724
rect 87344 45668 87400 45724
rect 87400 45668 87404 45724
rect 87340 45664 87404 45668
rect 6692 45180 6756 45184
rect 6692 45124 6696 45180
rect 6696 45124 6752 45180
rect 6752 45124 6756 45180
rect 6692 45120 6756 45124
rect 6772 45180 6836 45184
rect 6772 45124 6776 45180
rect 6776 45124 6832 45180
rect 6832 45124 6836 45180
rect 6772 45120 6836 45124
rect 6852 45180 6916 45184
rect 6852 45124 6856 45180
rect 6856 45124 6912 45180
rect 6912 45124 6916 45180
rect 6852 45120 6916 45124
rect 6932 45180 6996 45184
rect 6932 45124 6936 45180
rect 6936 45124 6992 45180
rect 6992 45124 6996 45180
rect 6932 45120 6996 45124
rect 87836 45180 87900 45184
rect 87836 45124 87840 45180
rect 87840 45124 87896 45180
rect 87896 45124 87900 45180
rect 87836 45120 87900 45124
rect 87916 45180 87980 45184
rect 87916 45124 87920 45180
rect 87920 45124 87976 45180
rect 87976 45124 87980 45180
rect 87916 45120 87980 45124
rect 87996 45180 88060 45184
rect 87996 45124 88000 45180
rect 88000 45124 88056 45180
rect 88056 45124 88060 45180
rect 87996 45120 88060 45124
rect 88076 45180 88140 45184
rect 88076 45124 88080 45180
rect 88080 45124 88136 45180
rect 88136 45124 88140 45180
rect 88076 45120 88140 45124
rect 5956 44636 6020 44640
rect 5956 44580 5960 44636
rect 5960 44580 6016 44636
rect 6016 44580 6020 44636
rect 5956 44576 6020 44580
rect 6036 44636 6100 44640
rect 6036 44580 6040 44636
rect 6040 44580 6096 44636
rect 6096 44580 6100 44636
rect 6036 44576 6100 44580
rect 6116 44636 6180 44640
rect 6116 44580 6120 44636
rect 6120 44580 6176 44636
rect 6176 44580 6180 44636
rect 6116 44576 6180 44580
rect 6196 44636 6260 44640
rect 6196 44580 6200 44636
rect 6200 44580 6256 44636
rect 6256 44580 6260 44636
rect 6196 44576 6260 44580
rect 87100 44636 87164 44640
rect 87100 44580 87104 44636
rect 87104 44580 87160 44636
rect 87160 44580 87164 44636
rect 87100 44576 87164 44580
rect 87180 44636 87244 44640
rect 87180 44580 87184 44636
rect 87184 44580 87240 44636
rect 87240 44580 87244 44636
rect 87180 44576 87244 44580
rect 87260 44636 87324 44640
rect 87260 44580 87264 44636
rect 87264 44580 87320 44636
rect 87320 44580 87324 44636
rect 87260 44576 87324 44580
rect 87340 44636 87404 44640
rect 87340 44580 87344 44636
rect 87344 44580 87400 44636
rect 87400 44580 87404 44636
rect 87340 44576 87404 44580
rect 6692 44092 6756 44096
rect 6692 44036 6696 44092
rect 6696 44036 6752 44092
rect 6752 44036 6756 44092
rect 6692 44032 6756 44036
rect 6772 44092 6836 44096
rect 6772 44036 6776 44092
rect 6776 44036 6832 44092
rect 6832 44036 6836 44092
rect 6772 44032 6836 44036
rect 6852 44092 6916 44096
rect 6852 44036 6856 44092
rect 6856 44036 6912 44092
rect 6912 44036 6916 44092
rect 6852 44032 6916 44036
rect 6932 44092 6996 44096
rect 6932 44036 6936 44092
rect 6936 44036 6992 44092
rect 6992 44036 6996 44092
rect 6932 44032 6996 44036
rect 87836 44092 87900 44096
rect 87836 44036 87840 44092
rect 87840 44036 87896 44092
rect 87896 44036 87900 44092
rect 87836 44032 87900 44036
rect 87916 44092 87980 44096
rect 87916 44036 87920 44092
rect 87920 44036 87976 44092
rect 87976 44036 87980 44092
rect 87916 44032 87980 44036
rect 87996 44092 88060 44096
rect 87996 44036 88000 44092
rect 88000 44036 88056 44092
rect 88056 44036 88060 44092
rect 87996 44032 88060 44036
rect 88076 44092 88140 44096
rect 88076 44036 88080 44092
rect 88080 44036 88136 44092
rect 88136 44036 88140 44092
rect 88076 44032 88140 44036
rect 5956 43548 6020 43552
rect 5956 43492 5960 43548
rect 5960 43492 6016 43548
rect 6016 43492 6020 43548
rect 5956 43488 6020 43492
rect 6036 43548 6100 43552
rect 6036 43492 6040 43548
rect 6040 43492 6096 43548
rect 6096 43492 6100 43548
rect 6036 43488 6100 43492
rect 6116 43548 6180 43552
rect 6116 43492 6120 43548
rect 6120 43492 6176 43548
rect 6176 43492 6180 43548
rect 6116 43488 6180 43492
rect 6196 43548 6260 43552
rect 6196 43492 6200 43548
rect 6200 43492 6256 43548
rect 6256 43492 6260 43548
rect 6196 43488 6260 43492
rect 87100 43548 87164 43552
rect 87100 43492 87104 43548
rect 87104 43492 87160 43548
rect 87160 43492 87164 43548
rect 87100 43488 87164 43492
rect 87180 43548 87244 43552
rect 87180 43492 87184 43548
rect 87184 43492 87240 43548
rect 87240 43492 87244 43548
rect 87180 43488 87244 43492
rect 87260 43548 87324 43552
rect 87260 43492 87264 43548
rect 87264 43492 87320 43548
rect 87320 43492 87324 43548
rect 87260 43488 87324 43492
rect 87340 43548 87404 43552
rect 87340 43492 87344 43548
rect 87344 43492 87400 43548
rect 87400 43492 87404 43548
rect 87340 43488 87404 43492
rect 6692 43004 6756 43008
rect 6692 42948 6696 43004
rect 6696 42948 6752 43004
rect 6752 42948 6756 43004
rect 6692 42944 6756 42948
rect 6772 43004 6836 43008
rect 6772 42948 6776 43004
rect 6776 42948 6832 43004
rect 6832 42948 6836 43004
rect 6772 42944 6836 42948
rect 6852 43004 6916 43008
rect 6852 42948 6856 43004
rect 6856 42948 6912 43004
rect 6912 42948 6916 43004
rect 6852 42944 6916 42948
rect 6932 43004 6996 43008
rect 6932 42948 6936 43004
rect 6936 42948 6992 43004
rect 6992 42948 6996 43004
rect 6932 42944 6996 42948
rect 87836 43004 87900 43008
rect 87836 42948 87840 43004
rect 87840 42948 87896 43004
rect 87896 42948 87900 43004
rect 87836 42944 87900 42948
rect 87916 43004 87980 43008
rect 87916 42948 87920 43004
rect 87920 42948 87976 43004
rect 87976 42948 87980 43004
rect 87916 42944 87980 42948
rect 87996 43004 88060 43008
rect 87996 42948 88000 43004
rect 88000 42948 88056 43004
rect 88056 42948 88060 43004
rect 87996 42944 88060 42948
rect 88076 43004 88140 43008
rect 88076 42948 88080 43004
rect 88080 42948 88136 43004
rect 88136 42948 88140 43004
rect 88076 42944 88140 42948
rect 5956 42460 6020 42464
rect 5956 42404 5960 42460
rect 5960 42404 6016 42460
rect 6016 42404 6020 42460
rect 5956 42400 6020 42404
rect 6036 42460 6100 42464
rect 6036 42404 6040 42460
rect 6040 42404 6096 42460
rect 6096 42404 6100 42460
rect 6036 42400 6100 42404
rect 6116 42460 6180 42464
rect 6116 42404 6120 42460
rect 6120 42404 6176 42460
rect 6176 42404 6180 42460
rect 6116 42400 6180 42404
rect 6196 42460 6260 42464
rect 6196 42404 6200 42460
rect 6200 42404 6256 42460
rect 6256 42404 6260 42460
rect 6196 42400 6260 42404
rect 87100 42460 87164 42464
rect 87100 42404 87104 42460
rect 87104 42404 87160 42460
rect 87160 42404 87164 42460
rect 87100 42400 87164 42404
rect 87180 42460 87244 42464
rect 87180 42404 87184 42460
rect 87184 42404 87240 42460
rect 87240 42404 87244 42460
rect 87180 42400 87244 42404
rect 87260 42460 87324 42464
rect 87260 42404 87264 42460
rect 87264 42404 87320 42460
rect 87320 42404 87324 42460
rect 87260 42400 87324 42404
rect 87340 42460 87404 42464
rect 87340 42404 87344 42460
rect 87344 42404 87400 42460
rect 87400 42404 87404 42460
rect 87340 42400 87404 42404
rect 6692 41916 6756 41920
rect 6692 41860 6696 41916
rect 6696 41860 6752 41916
rect 6752 41860 6756 41916
rect 6692 41856 6756 41860
rect 6772 41916 6836 41920
rect 6772 41860 6776 41916
rect 6776 41860 6832 41916
rect 6832 41860 6836 41916
rect 6772 41856 6836 41860
rect 6852 41916 6916 41920
rect 6852 41860 6856 41916
rect 6856 41860 6912 41916
rect 6912 41860 6916 41916
rect 6852 41856 6916 41860
rect 6932 41916 6996 41920
rect 6932 41860 6936 41916
rect 6936 41860 6992 41916
rect 6992 41860 6996 41916
rect 6932 41856 6996 41860
rect 87836 41916 87900 41920
rect 87836 41860 87840 41916
rect 87840 41860 87896 41916
rect 87896 41860 87900 41916
rect 87836 41856 87900 41860
rect 87916 41916 87980 41920
rect 87916 41860 87920 41916
rect 87920 41860 87976 41916
rect 87976 41860 87980 41916
rect 87916 41856 87980 41860
rect 87996 41916 88060 41920
rect 87996 41860 88000 41916
rect 88000 41860 88056 41916
rect 88056 41860 88060 41916
rect 87996 41856 88060 41860
rect 88076 41916 88140 41920
rect 88076 41860 88080 41916
rect 88080 41860 88136 41916
rect 88136 41860 88140 41916
rect 88076 41856 88140 41860
rect 5956 41372 6020 41376
rect 5956 41316 5960 41372
rect 5960 41316 6016 41372
rect 6016 41316 6020 41372
rect 5956 41312 6020 41316
rect 6036 41372 6100 41376
rect 6036 41316 6040 41372
rect 6040 41316 6096 41372
rect 6096 41316 6100 41372
rect 6036 41312 6100 41316
rect 6116 41372 6180 41376
rect 6116 41316 6120 41372
rect 6120 41316 6176 41372
rect 6176 41316 6180 41372
rect 6116 41312 6180 41316
rect 6196 41372 6260 41376
rect 6196 41316 6200 41372
rect 6200 41316 6256 41372
rect 6256 41316 6260 41372
rect 6196 41312 6260 41316
rect 87100 41372 87164 41376
rect 87100 41316 87104 41372
rect 87104 41316 87160 41372
rect 87160 41316 87164 41372
rect 87100 41312 87164 41316
rect 87180 41372 87244 41376
rect 87180 41316 87184 41372
rect 87184 41316 87240 41372
rect 87240 41316 87244 41372
rect 87180 41312 87244 41316
rect 87260 41372 87324 41376
rect 87260 41316 87264 41372
rect 87264 41316 87320 41372
rect 87320 41316 87324 41372
rect 87260 41312 87324 41316
rect 87340 41372 87404 41376
rect 87340 41316 87344 41372
rect 87344 41316 87400 41372
rect 87400 41316 87404 41372
rect 87340 41312 87404 41316
rect 6692 40828 6756 40832
rect 6692 40772 6696 40828
rect 6696 40772 6752 40828
rect 6752 40772 6756 40828
rect 6692 40768 6756 40772
rect 6772 40828 6836 40832
rect 6772 40772 6776 40828
rect 6776 40772 6832 40828
rect 6832 40772 6836 40828
rect 6772 40768 6836 40772
rect 6852 40828 6916 40832
rect 6852 40772 6856 40828
rect 6856 40772 6912 40828
rect 6912 40772 6916 40828
rect 6852 40768 6916 40772
rect 6932 40828 6996 40832
rect 6932 40772 6936 40828
rect 6936 40772 6992 40828
rect 6992 40772 6996 40828
rect 6932 40768 6996 40772
rect 87836 40828 87900 40832
rect 87836 40772 87840 40828
rect 87840 40772 87896 40828
rect 87896 40772 87900 40828
rect 87836 40768 87900 40772
rect 87916 40828 87980 40832
rect 87916 40772 87920 40828
rect 87920 40772 87976 40828
rect 87976 40772 87980 40828
rect 87916 40768 87980 40772
rect 87996 40828 88060 40832
rect 87996 40772 88000 40828
rect 88000 40772 88056 40828
rect 88056 40772 88060 40828
rect 87996 40768 88060 40772
rect 88076 40828 88140 40832
rect 88076 40772 88080 40828
rect 88080 40772 88136 40828
rect 88136 40772 88140 40828
rect 88076 40768 88140 40772
rect 5956 40284 6020 40288
rect 5956 40228 5960 40284
rect 5960 40228 6016 40284
rect 6016 40228 6020 40284
rect 5956 40224 6020 40228
rect 6036 40284 6100 40288
rect 6036 40228 6040 40284
rect 6040 40228 6096 40284
rect 6096 40228 6100 40284
rect 6036 40224 6100 40228
rect 6116 40284 6180 40288
rect 6116 40228 6120 40284
rect 6120 40228 6176 40284
rect 6176 40228 6180 40284
rect 6116 40224 6180 40228
rect 6196 40284 6260 40288
rect 6196 40228 6200 40284
rect 6200 40228 6256 40284
rect 6256 40228 6260 40284
rect 6196 40224 6260 40228
rect 87100 40284 87164 40288
rect 87100 40228 87104 40284
rect 87104 40228 87160 40284
rect 87160 40228 87164 40284
rect 87100 40224 87164 40228
rect 87180 40284 87244 40288
rect 87180 40228 87184 40284
rect 87184 40228 87240 40284
rect 87240 40228 87244 40284
rect 87180 40224 87244 40228
rect 87260 40284 87324 40288
rect 87260 40228 87264 40284
rect 87264 40228 87320 40284
rect 87320 40228 87324 40284
rect 87260 40224 87324 40228
rect 87340 40284 87404 40288
rect 87340 40228 87344 40284
rect 87344 40228 87400 40284
rect 87400 40228 87404 40284
rect 87340 40224 87404 40228
rect 6692 39740 6756 39744
rect 6692 39684 6696 39740
rect 6696 39684 6752 39740
rect 6752 39684 6756 39740
rect 6692 39680 6756 39684
rect 6772 39740 6836 39744
rect 6772 39684 6776 39740
rect 6776 39684 6832 39740
rect 6832 39684 6836 39740
rect 6772 39680 6836 39684
rect 6852 39740 6916 39744
rect 6852 39684 6856 39740
rect 6856 39684 6912 39740
rect 6912 39684 6916 39740
rect 6852 39680 6916 39684
rect 6932 39740 6996 39744
rect 6932 39684 6936 39740
rect 6936 39684 6992 39740
rect 6992 39684 6996 39740
rect 6932 39680 6996 39684
rect 87836 39740 87900 39744
rect 87836 39684 87840 39740
rect 87840 39684 87896 39740
rect 87896 39684 87900 39740
rect 87836 39680 87900 39684
rect 87916 39740 87980 39744
rect 87916 39684 87920 39740
rect 87920 39684 87976 39740
rect 87976 39684 87980 39740
rect 87916 39680 87980 39684
rect 87996 39740 88060 39744
rect 87996 39684 88000 39740
rect 88000 39684 88056 39740
rect 88056 39684 88060 39740
rect 87996 39680 88060 39684
rect 88076 39740 88140 39744
rect 88076 39684 88080 39740
rect 88080 39684 88136 39740
rect 88136 39684 88140 39740
rect 88076 39680 88140 39684
rect 5956 39196 6020 39200
rect 5956 39140 5960 39196
rect 5960 39140 6016 39196
rect 6016 39140 6020 39196
rect 5956 39136 6020 39140
rect 6036 39196 6100 39200
rect 6036 39140 6040 39196
rect 6040 39140 6096 39196
rect 6096 39140 6100 39196
rect 6036 39136 6100 39140
rect 6116 39196 6180 39200
rect 6116 39140 6120 39196
rect 6120 39140 6176 39196
rect 6176 39140 6180 39196
rect 6116 39136 6180 39140
rect 6196 39196 6260 39200
rect 6196 39140 6200 39196
rect 6200 39140 6256 39196
rect 6256 39140 6260 39196
rect 6196 39136 6260 39140
rect 87100 39196 87164 39200
rect 87100 39140 87104 39196
rect 87104 39140 87160 39196
rect 87160 39140 87164 39196
rect 87100 39136 87164 39140
rect 87180 39196 87244 39200
rect 87180 39140 87184 39196
rect 87184 39140 87240 39196
rect 87240 39140 87244 39196
rect 87180 39136 87244 39140
rect 87260 39196 87324 39200
rect 87260 39140 87264 39196
rect 87264 39140 87320 39196
rect 87320 39140 87324 39196
rect 87260 39136 87324 39140
rect 87340 39196 87404 39200
rect 87340 39140 87344 39196
rect 87344 39140 87400 39196
rect 87400 39140 87404 39196
rect 87340 39136 87404 39140
rect 6692 38652 6756 38656
rect 6692 38596 6696 38652
rect 6696 38596 6752 38652
rect 6752 38596 6756 38652
rect 6692 38592 6756 38596
rect 6772 38652 6836 38656
rect 6772 38596 6776 38652
rect 6776 38596 6832 38652
rect 6832 38596 6836 38652
rect 6772 38592 6836 38596
rect 6852 38652 6916 38656
rect 6852 38596 6856 38652
rect 6856 38596 6912 38652
rect 6912 38596 6916 38652
rect 6852 38592 6916 38596
rect 6932 38652 6996 38656
rect 6932 38596 6936 38652
rect 6936 38596 6992 38652
rect 6992 38596 6996 38652
rect 6932 38592 6996 38596
rect 87836 38652 87900 38656
rect 87836 38596 87840 38652
rect 87840 38596 87896 38652
rect 87896 38596 87900 38652
rect 87836 38592 87900 38596
rect 87916 38652 87980 38656
rect 87916 38596 87920 38652
rect 87920 38596 87976 38652
rect 87976 38596 87980 38652
rect 87916 38592 87980 38596
rect 87996 38652 88060 38656
rect 87996 38596 88000 38652
rect 88000 38596 88056 38652
rect 88056 38596 88060 38652
rect 87996 38592 88060 38596
rect 88076 38652 88140 38656
rect 88076 38596 88080 38652
rect 88080 38596 88136 38652
rect 88136 38596 88140 38652
rect 88076 38592 88140 38596
rect 5956 38108 6020 38112
rect 5956 38052 5960 38108
rect 5960 38052 6016 38108
rect 6016 38052 6020 38108
rect 5956 38048 6020 38052
rect 6036 38108 6100 38112
rect 6036 38052 6040 38108
rect 6040 38052 6096 38108
rect 6096 38052 6100 38108
rect 6036 38048 6100 38052
rect 6116 38108 6180 38112
rect 6116 38052 6120 38108
rect 6120 38052 6176 38108
rect 6176 38052 6180 38108
rect 6116 38048 6180 38052
rect 6196 38108 6260 38112
rect 6196 38052 6200 38108
rect 6200 38052 6256 38108
rect 6256 38052 6260 38108
rect 6196 38048 6260 38052
rect 87100 38108 87164 38112
rect 87100 38052 87104 38108
rect 87104 38052 87160 38108
rect 87160 38052 87164 38108
rect 87100 38048 87164 38052
rect 87180 38108 87244 38112
rect 87180 38052 87184 38108
rect 87184 38052 87240 38108
rect 87240 38052 87244 38108
rect 87180 38048 87244 38052
rect 87260 38108 87324 38112
rect 87260 38052 87264 38108
rect 87264 38052 87320 38108
rect 87320 38052 87324 38108
rect 87260 38048 87324 38052
rect 87340 38108 87404 38112
rect 87340 38052 87344 38108
rect 87344 38052 87400 38108
rect 87400 38052 87404 38108
rect 87340 38048 87404 38052
rect 6692 37564 6756 37568
rect 6692 37508 6696 37564
rect 6696 37508 6752 37564
rect 6752 37508 6756 37564
rect 6692 37504 6756 37508
rect 6772 37564 6836 37568
rect 6772 37508 6776 37564
rect 6776 37508 6832 37564
rect 6832 37508 6836 37564
rect 6772 37504 6836 37508
rect 6852 37564 6916 37568
rect 6852 37508 6856 37564
rect 6856 37508 6912 37564
rect 6912 37508 6916 37564
rect 6852 37504 6916 37508
rect 6932 37564 6996 37568
rect 6932 37508 6936 37564
rect 6936 37508 6992 37564
rect 6992 37508 6996 37564
rect 6932 37504 6996 37508
rect 87836 37564 87900 37568
rect 87836 37508 87840 37564
rect 87840 37508 87896 37564
rect 87896 37508 87900 37564
rect 87836 37504 87900 37508
rect 87916 37564 87980 37568
rect 87916 37508 87920 37564
rect 87920 37508 87976 37564
rect 87976 37508 87980 37564
rect 87916 37504 87980 37508
rect 87996 37564 88060 37568
rect 87996 37508 88000 37564
rect 88000 37508 88056 37564
rect 88056 37508 88060 37564
rect 87996 37504 88060 37508
rect 88076 37564 88140 37568
rect 88076 37508 88080 37564
rect 88080 37508 88136 37564
rect 88136 37508 88140 37564
rect 88076 37504 88140 37508
rect 5956 37020 6020 37024
rect 5956 36964 5960 37020
rect 5960 36964 6016 37020
rect 6016 36964 6020 37020
rect 5956 36960 6020 36964
rect 6036 37020 6100 37024
rect 6036 36964 6040 37020
rect 6040 36964 6096 37020
rect 6096 36964 6100 37020
rect 6036 36960 6100 36964
rect 6116 37020 6180 37024
rect 6116 36964 6120 37020
rect 6120 36964 6176 37020
rect 6176 36964 6180 37020
rect 6116 36960 6180 36964
rect 6196 37020 6260 37024
rect 6196 36964 6200 37020
rect 6200 36964 6256 37020
rect 6256 36964 6260 37020
rect 6196 36960 6260 36964
rect 87100 37020 87164 37024
rect 87100 36964 87104 37020
rect 87104 36964 87160 37020
rect 87160 36964 87164 37020
rect 87100 36960 87164 36964
rect 87180 37020 87244 37024
rect 87180 36964 87184 37020
rect 87184 36964 87240 37020
rect 87240 36964 87244 37020
rect 87180 36960 87244 36964
rect 87260 37020 87324 37024
rect 87260 36964 87264 37020
rect 87264 36964 87320 37020
rect 87320 36964 87324 37020
rect 87260 36960 87324 36964
rect 87340 37020 87404 37024
rect 87340 36964 87344 37020
rect 87344 36964 87400 37020
rect 87400 36964 87404 37020
rect 87340 36960 87404 36964
rect 6692 36476 6756 36480
rect 6692 36420 6696 36476
rect 6696 36420 6752 36476
rect 6752 36420 6756 36476
rect 6692 36416 6756 36420
rect 6772 36476 6836 36480
rect 6772 36420 6776 36476
rect 6776 36420 6832 36476
rect 6832 36420 6836 36476
rect 6772 36416 6836 36420
rect 6852 36476 6916 36480
rect 6852 36420 6856 36476
rect 6856 36420 6912 36476
rect 6912 36420 6916 36476
rect 6852 36416 6916 36420
rect 6932 36476 6996 36480
rect 6932 36420 6936 36476
rect 6936 36420 6992 36476
rect 6992 36420 6996 36476
rect 6932 36416 6996 36420
rect 87836 36476 87900 36480
rect 87836 36420 87840 36476
rect 87840 36420 87896 36476
rect 87896 36420 87900 36476
rect 87836 36416 87900 36420
rect 87916 36476 87980 36480
rect 87916 36420 87920 36476
rect 87920 36420 87976 36476
rect 87976 36420 87980 36476
rect 87916 36416 87980 36420
rect 87996 36476 88060 36480
rect 87996 36420 88000 36476
rect 88000 36420 88056 36476
rect 88056 36420 88060 36476
rect 87996 36416 88060 36420
rect 88076 36476 88140 36480
rect 88076 36420 88080 36476
rect 88080 36420 88136 36476
rect 88136 36420 88140 36476
rect 88076 36416 88140 36420
rect 5956 35932 6020 35936
rect 5956 35876 5960 35932
rect 5960 35876 6016 35932
rect 6016 35876 6020 35932
rect 5956 35872 6020 35876
rect 6036 35932 6100 35936
rect 6036 35876 6040 35932
rect 6040 35876 6096 35932
rect 6096 35876 6100 35932
rect 6036 35872 6100 35876
rect 6116 35932 6180 35936
rect 6116 35876 6120 35932
rect 6120 35876 6176 35932
rect 6176 35876 6180 35932
rect 6116 35872 6180 35876
rect 6196 35932 6260 35936
rect 6196 35876 6200 35932
rect 6200 35876 6256 35932
rect 6256 35876 6260 35932
rect 6196 35872 6260 35876
rect 87100 35932 87164 35936
rect 87100 35876 87104 35932
rect 87104 35876 87160 35932
rect 87160 35876 87164 35932
rect 87100 35872 87164 35876
rect 87180 35932 87244 35936
rect 87180 35876 87184 35932
rect 87184 35876 87240 35932
rect 87240 35876 87244 35932
rect 87180 35872 87244 35876
rect 87260 35932 87324 35936
rect 87260 35876 87264 35932
rect 87264 35876 87320 35932
rect 87320 35876 87324 35932
rect 87260 35872 87324 35876
rect 87340 35932 87404 35936
rect 87340 35876 87344 35932
rect 87344 35876 87400 35932
rect 87400 35876 87404 35932
rect 87340 35872 87404 35876
rect 6692 35388 6756 35392
rect 6692 35332 6696 35388
rect 6696 35332 6752 35388
rect 6752 35332 6756 35388
rect 6692 35328 6756 35332
rect 6772 35388 6836 35392
rect 6772 35332 6776 35388
rect 6776 35332 6832 35388
rect 6832 35332 6836 35388
rect 6772 35328 6836 35332
rect 6852 35388 6916 35392
rect 6852 35332 6856 35388
rect 6856 35332 6912 35388
rect 6912 35332 6916 35388
rect 6852 35328 6916 35332
rect 6932 35388 6996 35392
rect 6932 35332 6936 35388
rect 6936 35332 6992 35388
rect 6992 35332 6996 35388
rect 6932 35328 6996 35332
rect 87836 35388 87900 35392
rect 87836 35332 87840 35388
rect 87840 35332 87896 35388
rect 87896 35332 87900 35388
rect 87836 35328 87900 35332
rect 87916 35388 87980 35392
rect 87916 35332 87920 35388
rect 87920 35332 87976 35388
rect 87976 35332 87980 35388
rect 87916 35328 87980 35332
rect 87996 35388 88060 35392
rect 87996 35332 88000 35388
rect 88000 35332 88056 35388
rect 88056 35332 88060 35388
rect 87996 35328 88060 35332
rect 88076 35388 88140 35392
rect 88076 35332 88080 35388
rect 88080 35332 88136 35388
rect 88136 35332 88140 35388
rect 88076 35328 88140 35332
rect 5956 34844 6020 34848
rect 5956 34788 5960 34844
rect 5960 34788 6016 34844
rect 6016 34788 6020 34844
rect 5956 34784 6020 34788
rect 6036 34844 6100 34848
rect 6036 34788 6040 34844
rect 6040 34788 6096 34844
rect 6096 34788 6100 34844
rect 6036 34784 6100 34788
rect 6116 34844 6180 34848
rect 6116 34788 6120 34844
rect 6120 34788 6176 34844
rect 6176 34788 6180 34844
rect 6116 34784 6180 34788
rect 6196 34844 6260 34848
rect 6196 34788 6200 34844
rect 6200 34788 6256 34844
rect 6256 34788 6260 34844
rect 6196 34784 6260 34788
rect 87100 34844 87164 34848
rect 87100 34788 87104 34844
rect 87104 34788 87160 34844
rect 87160 34788 87164 34844
rect 87100 34784 87164 34788
rect 87180 34844 87244 34848
rect 87180 34788 87184 34844
rect 87184 34788 87240 34844
rect 87240 34788 87244 34844
rect 87180 34784 87244 34788
rect 87260 34844 87324 34848
rect 87260 34788 87264 34844
rect 87264 34788 87320 34844
rect 87320 34788 87324 34844
rect 87260 34784 87324 34788
rect 87340 34844 87404 34848
rect 87340 34788 87344 34844
rect 87344 34788 87400 34844
rect 87400 34788 87404 34844
rect 87340 34784 87404 34788
rect 6692 34300 6756 34304
rect 6692 34244 6696 34300
rect 6696 34244 6752 34300
rect 6752 34244 6756 34300
rect 6692 34240 6756 34244
rect 6772 34300 6836 34304
rect 6772 34244 6776 34300
rect 6776 34244 6832 34300
rect 6832 34244 6836 34300
rect 6772 34240 6836 34244
rect 6852 34300 6916 34304
rect 6852 34244 6856 34300
rect 6856 34244 6912 34300
rect 6912 34244 6916 34300
rect 6852 34240 6916 34244
rect 6932 34300 6996 34304
rect 6932 34244 6936 34300
rect 6936 34244 6992 34300
rect 6992 34244 6996 34300
rect 6932 34240 6996 34244
rect 87836 34300 87900 34304
rect 87836 34244 87840 34300
rect 87840 34244 87896 34300
rect 87896 34244 87900 34300
rect 87836 34240 87900 34244
rect 87916 34300 87980 34304
rect 87916 34244 87920 34300
rect 87920 34244 87976 34300
rect 87976 34244 87980 34300
rect 87916 34240 87980 34244
rect 87996 34300 88060 34304
rect 87996 34244 88000 34300
rect 88000 34244 88056 34300
rect 88056 34244 88060 34300
rect 87996 34240 88060 34244
rect 88076 34300 88140 34304
rect 88076 34244 88080 34300
rect 88080 34244 88136 34300
rect 88136 34244 88140 34300
rect 88076 34240 88140 34244
rect 5956 33756 6020 33760
rect 5956 33700 5960 33756
rect 5960 33700 6016 33756
rect 6016 33700 6020 33756
rect 5956 33696 6020 33700
rect 6036 33756 6100 33760
rect 6036 33700 6040 33756
rect 6040 33700 6096 33756
rect 6096 33700 6100 33756
rect 6036 33696 6100 33700
rect 6116 33756 6180 33760
rect 6116 33700 6120 33756
rect 6120 33700 6176 33756
rect 6176 33700 6180 33756
rect 6116 33696 6180 33700
rect 6196 33756 6260 33760
rect 6196 33700 6200 33756
rect 6200 33700 6256 33756
rect 6256 33700 6260 33756
rect 6196 33696 6260 33700
rect 87100 33756 87164 33760
rect 87100 33700 87104 33756
rect 87104 33700 87160 33756
rect 87160 33700 87164 33756
rect 87100 33696 87164 33700
rect 87180 33756 87244 33760
rect 87180 33700 87184 33756
rect 87184 33700 87240 33756
rect 87240 33700 87244 33756
rect 87180 33696 87244 33700
rect 87260 33756 87324 33760
rect 87260 33700 87264 33756
rect 87264 33700 87320 33756
rect 87320 33700 87324 33756
rect 87260 33696 87324 33700
rect 87340 33756 87404 33760
rect 87340 33700 87344 33756
rect 87344 33700 87400 33756
rect 87400 33700 87404 33756
rect 87340 33696 87404 33700
rect 6692 33212 6756 33216
rect 6692 33156 6696 33212
rect 6696 33156 6752 33212
rect 6752 33156 6756 33212
rect 6692 33152 6756 33156
rect 6772 33212 6836 33216
rect 6772 33156 6776 33212
rect 6776 33156 6832 33212
rect 6832 33156 6836 33212
rect 6772 33152 6836 33156
rect 6852 33212 6916 33216
rect 6852 33156 6856 33212
rect 6856 33156 6912 33212
rect 6912 33156 6916 33212
rect 6852 33152 6916 33156
rect 6932 33212 6996 33216
rect 6932 33156 6936 33212
rect 6936 33156 6992 33212
rect 6992 33156 6996 33212
rect 6932 33152 6996 33156
rect 87836 33212 87900 33216
rect 87836 33156 87840 33212
rect 87840 33156 87896 33212
rect 87896 33156 87900 33212
rect 87836 33152 87900 33156
rect 87916 33212 87980 33216
rect 87916 33156 87920 33212
rect 87920 33156 87976 33212
rect 87976 33156 87980 33212
rect 87916 33152 87980 33156
rect 87996 33212 88060 33216
rect 87996 33156 88000 33212
rect 88000 33156 88056 33212
rect 88056 33156 88060 33212
rect 87996 33152 88060 33156
rect 88076 33212 88140 33216
rect 88076 33156 88080 33212
rect 88080 33156 88136 33212
rect 88136 33156 88140 33212
rect 88076 33152 88140 33156
rect 5956 32668 6020 32672
rect 5956 32612 5960 32668
rect 5960 32612 6016 32668
rect 6016 32612 6020 32668
rect 5956 32608 6020 32612
rect 6036 32668 6100 32672
rect 6036 32612 6040 32668
rect 6040 32612 6096 32668
rect 6096 32612 6100 32668
rect 6036 32608 6100 32612
rect 6116 32668 6180 32672
rect 6116 32612 6120 32668
rect 6120 32612 6176 32668
rect 6176 32612 6180 32668
rect 6116 32608 6180 32612
rect 6196 32668 6260 32672
rect 6196 32612 6200 32668
rect 6200 32612 6256 32668
rect 6256 32612 6260 32668
rect 6196 32608 6260 32612
rect 87100 32668 87164 32672
rect 87100 32612 87104 32668
rect 87104 32612 87160 32668
rect 87160 32612 87164 32668
rect 87100 32608 87164 32612
rect 87180 32668 87244 32672
rect 87180 32612 87184 32668
rect 87184 32612 87240 32668
rect 87240 32612 87244 32668
rect 87180 32608 87244 32612
rect 87260 32668 87324 32672
rect 87260 32612 87264 32668
rect 87264 32612 87320 32668
rect 87320 32612 87324 32668
rect 87260 32608 87324 32612
rect 87340 32668 87404 32672
rect 87340 32612 87344 32668
rect 87344 32612 87400 32668
rect 87400 32612 87404 32668
rect 87340 32608 87404 32612
rect 6692 32124 6756 32128
rect 6692 32068 6696 32124
rect 6696 32068 6752 32124
rect 6752 32068 6756 32124
rect 6692 32064 6756 32068
rect 6772 32124 6836 32128
rect 6772 32068 6776 32124
rect 6776 32068 6832 32124
rect 6832 32068 6836 32124
rect 6772 32064 6836 32068
rect 6852 32124 6916 32128
rect 6852 32068 6856 32124
rect 6856 32068 6912 32124
rect 6912 32068 6916 32124
rect 6852 32064 6916 32068
rect 6932 32124 6996 32128
rect 6932 32068 6936 32124
rect 6936 32068 6992 32124
rect 6992 32068 6996 32124
rect 6932 32064 6996 32068
rect 87836 32124 87900 32128
rect 87836 32068 87840 32124
rect 87840 32068 87896 32124
rect 87896 32068 87900 32124
rect 87836 32064 87900 32068
rect 87916 32124 87980 32128
rect 87916 32068 87920 32124
rect 87920 32068 87976 32124
rect 87976 32068 87980 32124
rect 87916 32064 87980 32068
rect 87996 32124 88060 32128
rect 87996 32068 88000 32124
rect 88000 32068 88056 32124
rect 88056 32068 88060 32124
rect 87996 32064 88060 32068
rect 88076 32124 88140 32128
rect 88076 32068 88080 32124
rect 88080 32068 88136 32124
rect 88136 32068 88140 32124
rect 88076 32064 88140 32068
rect 5956 31580 6020 31584
rect 5956 31524 5960 31580
rect 5960 31524 6016 31580
rect 6016 31524 6020 31580
rect 5956 31520 6020 31524
rect 6036 31580 6100 31584
rect 6036 31524 6040 31580
rect 6040 31524 6096 31580
rect 6096 31524 6100 31580
rect 6036 31520 6100 31524
rect 6116 31580 6180 31584
rect 6116 31524 6120 31580
rect 6120 31524 6176 31580
rect 6176 31524 6180 31580
rect 6116 31520 6180 31524
rect 6196 31580 6260 31584
rect 6196 31524 6200 31580
rect 6200 31524 6256 31580
rect 6256 31524 6260 31580
rect 6196 31520 6260 31524
rect 87100 31580 87164 31584
rect 87100 31524 87104 31580
rect 87104 31524 87160 31580
rect 87160 31524 87164 31580
rect 87100 31520 87164 31524
rect 87180 31580 87244 31584
rect 87180 31524 87184 31580
rect 87184 31524 87240 31580
rect 87240 31524 87244 31580
rect 87180 31520 87244 31524
rect 87260 31580 87324 31584
rect 87260 31524 87264 31580
rect 87264 31524 87320 31580
rect 87320 31524 87324 31580
rect 87260 31520 87324 31524
rect 87340 31580 87404 31584
rect 87340 31524 87344 31580
rect 87344 31524 87400 31580
rect 87400 31524 87404 31580
rect 87340 31520 87404 31524
rect 6692 31036 6756 31040
rect 6692 30980 6696 31036
rect 6696 30980 6752 31036
rect 6752 30980 6756 31036
rect 6692 30976 6756 30980
rect 6772 31036 6836 31040
rect 6772 30980 6776 31036
rect 6776 30980 6832 31036
rect 6832 30980 6836 31036
rect 6772 30976 6836 30980
rect 6852 31036 6916 31040
rect 6852 30980 6856 31036
rect 6856 30980 6912 31036
rect 6912 30980 6916 31036
rect 6852 30976 6916 30980
rect 6932 31036 6996 31040
rect 6932 30980 6936 31036
rect 6936 30980 6992 31036
rect 6992 30980 6996 31036
rect 6932 30976 6996 30980
rect 87836 31036 87900 31040
rect 87836 30980 87840 31036
rect 87840 30980 87896 31036
rect 87896 30980 87900 31036
rect 87836 30976 87900 30980
rect 87916 31036 87980 31040
rect 87916 30980 87920 31036
rect 87920 30980 87976 31036
rect 87976 30980 87980 31036
rect 87916 30976 87980 30980
rect 87996 31036 88060 31040
rect 87996 30980 88000 31036
rect 88000 30980 88056 31036
rect 88056 30980 88060 31036
rect 87996 30976 88060 30980
rect 88076 31036 88140 31040
rect 88076 30980 88080 31036
rect 88080 30980 88136 31036
rect 88136 30980 88140 31036
rect 88076 30976 88140 30980
rect 5956 30492 6020 30496
rect 5956 30436 5960 30492
rect 5960 30436 6016 30492
rect 6016 30436 6020 30492
rect 5956 30432 6020 30436
rect 6036 30492 6100 30496
rect 6036 30436 6040 30492
rect 6040 30436 6096 30492
rect 6096 30436 6100 30492
rect 6036 30432 6100 30436
rect 6116 30492 6180 30496
rect 6116 30436 6120 30492
rect 6120 30436 6176 30492
rect 6176 30436 6180 30492
rect 6116 30432 6180 30436
rect 6196 30492 6260 30496
rect 6196 30436 6200 30492
rect 6200 30436 6256 30492
rect 6256 30436 6260 30492
rect 6196 30432 6260 30436
rect 87100 30492 87164 30496
rect 87100 30436 87104 30492
rect 87104 30436 87160 30492
rect 87160 30436 87164 30492
rect 87100 30432 87164 30436
rect 87180 30492 87244 30496
rect 87180 30436 87184 30492
rect 87184 30436 87240 30492
rect 87240 30436 87244 30492
rect 87180 30432 87244 30436
rect 87260 30492 87324 30496
rect 87260 30436 87264 30492
rect 87264 30436 87320 30492
rect 87320 30436 87324 30492
rect 87260 30432 87324 30436
rect 87340 30492 87404 30496
rect 87340 30436 87344 30492
rect 87344 30436 87400 30492
rect 87400 30436 87404 30492
rect 87340 30432 87404 30436
rect 6692 29948 6756 29952
rect 6692 29892 6696 29948
rect 6696 29892 6752 29948
rect 6752 29892 6756 29948
rect 6692 29888 6756 29892
rect 6772 29948 6836 29952
rect 6772 29892 6776 29948
rect 6776 29892 6832 29948
rect 6832 29892 6836 29948
rect 6772 29888 6836 29892
rect 6852 29948 6916 29952
rect 6852 29892 6856 29948
rect 6856 29892 6912 29948
rect 6912 29892 6916 29948
rect 6852 29888 6916 29892
rect 6932 29948 6996 29952
rect 6932 29892 6936 29948
rect 6936 29892 6992 29948
rect 6992 29892 6996 29948
rect 6932 29888 6996 29892
rect 87836 29948 87900 29952
rect 87836 29892 87840 29948
rect 87840 29892 87896 29948
rect 87896 29892 87900 29948
rect 87836 29888 87900 29892
rect 87916 29948 87980 29952
rect 87916 29892 87920 29948
rect 87920 29892 87976 29948
rect 87976 29892 87980 29948
rect 87916 29888 87980 29892
rect 87996 29948 88060 29952
rect 87996 29892 88000 29948
rect 88000 29892 88056 29948
rect 88056 29892 88060 29948
rect 87996 29888 88060 29892
rect 88076 29948 88140 29952
rect 88076 29892 88080 29948
rect 88080 29892 88136 29948
rect 88136 29892 88140 29948
rect 88076 29888 88140 29892
rect 5956 29404 6020 29408
rect 5956 29348 5960 29404
rect 5960 29348 6016 29404
rect 6016 29348 6020 29404
rect 5956 29344 6020 29348
rect 6036 29404 6100 29408
rect 6036 29348 6040 29404
rect 6040 29348 6096 29404
rect 6096 29348 6100 29404
rect 6036 29344 6100 29348
rect 6116 29404 6180 29408
rect 6116 29348 6120 29404
rect 6120 29348 6176 29404
rect 6176 29348 6180 29404
rect 6116 29344 6180 29348
rect 6196 29404 6260 29408
rect 6196 29348 6200 29404
rect 6200 29348 6256 29404
rect 6256 29348 6260 29404
rect 6196 29344 6260 29348
rect 87100 29404 87164 29408
rect 87100 29348 87104 29404
rect 87104 29348 87160 29404
rect 87160 29348 87164 29404
rect 87100 29344 87164 29348
rect 87180 29404 87244 29408
rect 87180 29348 87184 29404
rect 87184 29348 87240 29404
rect 87240 29348 87244 29404
rect 87180 29344 87244 29348
rect 87260 29404 87324 29408
rect 87260 29348 87264 29404
rect 87264 29348 87320 29404
rect 87320 29348 87324 29404
rect 87260 29344 87324 29348
rect 87340 29404 87404 29408
rect 87340 29348 87344 29404
rect 87344 29348 87400 29404
rect 87400 29348 87404 29404
rect 87340 29344 87404 29348
rect 6692 28860 6756 28864
rect 6692 28804 6696 28860
rect 6696 28804 6752 28860
rect 6752 28804 6756 28860
rect 6692 28800 6756 28804
rect 6772 28860 6836 28864
rect 6772 28804 6776 28860
rect 6776 28804 6832 28860
rect 6832 28804 6836 28860
rect 6772 28800 6836 28804
rect 6852 28860 6916 28864
rect 6852 28804 6856 28860
rect 6856 28804 6912 28860
rect 6912 28804 6916 28860
rect 6852 28800 6916 28804
rect 6932 28860 6996 28864
rect 6932 28804 6936 28860
rect 6936 28804 6992 28860
rect 6992 28804 6996 28860
rect 6932 28800 6996 28804
rect 87836 28860 87900 28864
rect 87836 28804 87840 28860
rect 87840 28804 87896 28860
rect 87896 28804 87900 28860
rect 87836 28800 87900 28804
rect 87916 28860 87980 28864
rect 87916 28804 87920 28860
rect 87920 28804 87976 28860
rect 87976 28804 87980 28860
rect 87916 28800 87980 28804
rect 87996 28860 88060 28864
rect 87996 28804 88000 28860
rect 88000 28804 88056 28860
rect 88056 28804 88060 28860
rect 87996 28800 88060 28804
rect 88076 28860 88140 28864
rect 88076 28804 88080 28860
rect 88080 28804 88136 28860
rect 88136 28804 88140 28860
rect 88076 28800 88140 28804
rect 5956 28316 6020 28320
rect 5956 28260 5960 28316
rect 5960 28260 6016 28316
rect 6016 28260 6020 28316
rect 5956 28256 6020 28260
rect 6036 28316 6100 28320
rect 6036 28260 6040 28316
rect 6040 28260 6096 28316
rect 6096 28260 6100 28316
rect 6036 28256 6100 28260
rect 6116 28316 6180 28320
rect 6116 28260 6120 28316
rect 6120 28260 6176 28316
rect 6176 28260 6180 28316
rect 6116 28256 6180 28260
rect 6196 28316 6260 28320
rect 6196 28260 6200 28316
rect 6200 28260 6256 28316
rect 6256 28260 6260 28316
rect 6196 28256 6260 28260
rect 87100 28316 87164 28320
rect 87100 28260 87104 28316
rect 87104 28260 87160 28316
rect 87160 28260 87164 28316
rect 87100 28256 87164 28260
rect 87180 28316 87244 28320
rect 87180 28260 87184 28316
rect 87184 28260 87240 28316
rect 87240 28260 87244 28316
rect 87180 28256 87244 28260
rect 87260 28316 87324 28320
rect 87260 28260 87264 28316
rect 87264 28260 87320 28316
rect 87320 28260 87324 28316
rect 87260 28256 87324 28260
rect 87340 28316 87404 28320
rect 87340 28260 87344 28316
rect 87344 28260 87400 28316
rect 87400 28260 87404 28316
rect 87340 28256 87404 28260
rect 6692 27772 6756 27776
rect 6692 27716 6696 27772
rect 6696 27716 6752 27772
rect 6752 27716 6756 27772
rect 6692 27712 6756 27716
rect 6772 27772 6836 27776
rect 6772 27716 6776 27772
rect 6776 27716 6832 27772
rect 6832 27716 6836 27772
rect 6772 27712 6836 27716
rect 6852 27772 6916 27776
rect 6852 27716 6856 27772
rect 6856 27716 6912 27772
rect 6912 27716 6916 27772
rect 6852 27712 6916 27716
rect 6932 27772 6996 27776
rect 6932 27716 6936 27772
rect 6936 27716 6992 27772
rect 6992 27716 6996 27772
rect 6932 27712 6996 27716
rect 87836 27772 87900 27776
rect 87836 27716 87840 27772
rect 87840 27716 87896 27772
rect 87896 27716 87900 27772
rect 87836 27712 87900 27716
rect 87916 27772 87980 27776
rect 87916 27716 87920 27772
rect 87920 27716 87976 27772
rect 87976 27716 87980 27772
rect 87916 27712 87980 27716
rect 87996 27772 88060 27776
rect 87996 27716 88000 27772
rect 88000 27716 88056 27772
rect 88056 27716 88060 27772
rect 87996 27712 88060 27716
rect 88076 27772 88140 27776
rect 88076 27716 88080 27772
rect 88080 27716 88136 27772
rect 88136 27716 88140 27772
rect 88076 27712 88140 27716
rect 5956 27228 6020 27232
rect 5956 27172 5960 27228
rect 5960 27172 6016 27228
rect 6016 27172 6020 27228
rect 5956 27168 6020 27172
rect 6036 27228 6100 27232
rect 6036 27172 6040 27228
rect 6040 27172 6096 27228
rect 6096 27172 6100 27228
rect 6036 27168 6100 27172
rect 6116 27228 6180 27232
rect 6116 27172 6120 27228
rect 6120 27172 6176 27228
rect 6176 27172 6180 27228
rect 6116 27168 6180 27172
rect 6196 27228 6260 27232
rect 6196 27172 6200 27228
rect 6200 27172 6256 27228
rect 6256 27172 6260 27228
rect 6196 27168 6260 27172
rect 87100 27228 87164 27232
rect 87100 27172 87104 27228
rect 87104 27172 87160 27228
rect 87160 27172 87164 27228
rect 87100 27168 87164 27172
rect 87180 27228 87244 27232
rect 87180 27172 87184 27228
rect 87184 27172 87240 27228
rect 87240 27172 87244 27228
rect 87180 27168 87244 27172
rect 87260 27228 87324 27232
rect 87260 27172 87264 27228
rect 87264 27172 87320 27228
rect 87320 27172 87324 27228
rect 87260 27168 87324 27172
rect 87340 27228 87404 27232
rect 87340 27172 87344 27228
rect 87344 27172 87400 27228
rect 87400 27172 87404 27228
rect 87340 27168 87404 27172
rect 6692 26684 6756 26688
rect 6692 26628 6696 26684
rect 6696 26628 6752 26684
rect 6752 26628 6756 26684
rect 6692 26624 6756 26628
rect 6772 26684 6836 26688
rect 6772 26628 6776 26684
rect 6776 26628 6832 26684
rect 6832 26628 6836 26684
rect 6772 26624 6836 26628
rect 6852 26684 6916 26688
rect 6852 26628 6856 26684
rect 6856 26628 6912 26684
rect 6912 26628 6916 26684
rect 6852 26624 6916 26628
rect 6932 26684 6996 26688
rect 6932 26628 6936 26684
rect 6936 26628 6992 26684
rect 6992 26628 6996 26684
rect 6932 26624 6996 26628
rect 87836 26684 87900 26688
rect 87836 26628 87840 26684
rect 87840 26628 87896 26684
rect 87896 26628 87900 26684
rect 87836 26624 87900 26628
rect 87916 26684 87980 26688
rect 87916 26628 87920 26684
rect 87920 26628 87976 26684
rect 87976 26628 87980 26684
rect 87916 26624 87980 26628
rect 87996 26684 88060 26688
rect 87996 26628 88000 26684
rect 88000 26628 88056 26684
rect 88056 26628 88060 26684
rect 87996 26624 88060 26628
rect 88076 26684 88140 26688
rect 88076 26628 88080 26684
rect 88080 26628 88136 26684
rect 88136 26628 88140 26684
rect 88076 26624 88140 26628
rect 5956 26140 6020 26144
rect 5956 26084 5960 26140
rect 5960 26084 6016 26140
rect 6016 26084 6020 26140
rect 5956 26080 6020 26084
rect 6036 26140 6100 26144
rect 6036 26084 6040 26140
rect 6040 26084 6096 26140
rect 6096 26084 6100 26140
rect 6036 26080 6100 26084
rect 6116 26140 6180 26144
rect 6116 26084 6120 26140
rect 6120 26084 6176 26140
rect 6176 26084 6180 26140
rect 6116 26080 6180 26084
rect 6196 26140 6260 26144
rect 6196 26084 6200 26140
rect 6200 26084 6256 26140
rect 6256 26084 6260 26140
rect 6196 26080 6260 26084
rect 87100 26140 87164 26144
rect 87100 26084 87104 26140
rect 87104 26084 87160 26140
rect 87160 26084 87164 26140
rect 87100 26080 87164 26084
rect 87180 26140 87244 26144
rect 87180 26084 87184 26140
rect 87184 26084 87240 26140
rect 87240 26084 87244 26140
rect 87180 26080 87244 26084
rect 87260 26140 87324 26144
rect 87260 26084 87264 26140
rect 87264 26084 87320 26140
rect 87320 26084 87324 26140
rect 87260 26080 87324 26084
rect 87340 26140 87404 26144
rect 87340 26084 87344 26140
rect 87344 26084 87400 26140
rect 87400 26084 87404 26140
rect 87340 26080 87404 26084
rect 6692 25596 6756 25600
rect 6692 25540 6696 25596
rect 6696 25540 6752 25596
rect 6752 25540 6756 25596
rect 6692 25536 6756 25540
rect 6772 25596 6836 25600
rect 6772 25540 6776 25596
rect 6776 25540 6832 25596
rect 6832 25540 6836 25596
rect 6772 25536 6836 25540
rect 6852 25596 6916 25600
rect 6852 25540 6856 25596
rect 6856 25540 6912 25596
rect 6912 25540 6916 25596
rect 6852 25536 6916 25540
rect 6932 25596 6996 25600
rect 6932 25540 6936 25596
rect 6936 25540 6992 25596
rect 6992 25540 6996 25596
rect 6932 25536 6996 25540
rect 87836 25596 87900 25600
rect 87836 25540 87840 25596
rect 87840 25540 87896 25596
rect 87896 25540 87900 25596
rect 87836 25536 87900 25540
rect 87916 25596 87980 25600
rect 87916 25540 87920 25596
rect 87920 25540 87976 25596
rect 87976 25540 87980 25596
rect 87916 25536 87980 25540
rect 87996 25596 88060 25600
rect 87996 25540 88000 25596
rect 88000 25540 88056 25596
rect 88056 25540 88060 25596
rect 87996 25536 88060 25540
rect 88076 25596 88140 25600
rect 88076 25540 88080 25596
rect 88080 25540 88136 25596
rect 88136 25540 88140 25596
rect 88076 25536 88140 25540
rect 5956 25052 6020 25056
rect 5956 24996 5960 25052
rect 5960 24996 6016 25052
rect 6016 24996 6020 25052
rect 5956 24992 6020 24996
rect 6036 25052 6100 25056
rect 6036 24996 6040 25052
rect 6040 24996 6096 25052
rect 6096 24996 6100 25052
rect 6036 24992 6100 24996
rect 6116 25052 6180 25056
rect 6116 24996 6120 25052
rect 6120 24996 6176 25052
rect 6176 24996 6180 25052
rect 6116 24992 6180 24996
rect 6196 25052 6260 25056
rect 6196 24996 6200 25052
rect 6200 24996 6256 25052
rect 6256 24996 6260 25052
rect 6196 24992 6260 24996
rect 87100 25052 87164 25056
rect 87100 24996 87104 25052
rect 87104 24996 87160 25052
rect 87160 24996 87164 25052
rect 87100 24992 87164 24996
rect 87180 25052 87244 25056
rect 87180 24996 87184 25052
rect 87184 24996 87240 25052
rect 87240 24996 87244 25052
rect 87180 24992 87244 24996
rect 87260 25052 87324 25056
rect 87260 24996 87264 25052
rect 87264 24996 87320 25052
rect 87320 24996 87324 25052
rect 87260 24992 87324 24996
rect 87340 25052 87404 25056
rect 87340 24996 87344 25052
rect 87344 24996 87400 25052
rect 87400 24996 87404 25052
rect 87340 24992 87404 24996
rect 6692 24508 6756 24512
rect 6692 24452 6696 24508
rect 6696 24452 6752 24508
rect 6752 24452 6756 24508
rect 6692 24448 6756 24452
rect 6772 24508 6836 24512
rect 6772 24452 6776 24508
rect 6776 24452 6832 24508
rect 6832 24452 6836 24508
rect 6772 24448 6836 24452
rect 6852 24508 6916 24512
rect 6852 24452 6856 24508
rect 6856 24452 6912 24508
rect 6912 24452 6916 24508
rect 6852 24448 6916 24452
rect 6932 24508 6996 24512
rect 6932 24452 6936 24508
rect 6936 24452 6992 24508
rect 6992 24452 6996 24508
rect 6932 24448 6996 24452
rect 87836 24508 87900 24512
rect 87836 24452 87840 24508
rect 87840 24452 87896 24508
rect 87896 24452 87900 24508
rect 87836 24448 87900 24452
rect 87916 24508 87980 24512
rect 87916 24452 87920 24508
rect 87920 24452 87976 24508
rect 87976 24452 87980 24508
rect 87916 24448 87980 24452
rect 87996 24508 88060 24512
rect 87996 24452 88000 24508
rect 88000 24452 88056 24508
rect 88056 24452 88060 24508
rect 87996 24448 88060 24452
rect 88076 24508 88140 24512
rect 88076 24452 88080 24508
rect 88080 24452 88136 24508
rect 88136 24452 88140 24508
rect 88076 24448 88140 24452
rect 5956 23964 6020 23968
rect 5956 23908 5960 23964
rect 5960 23908 6016 23964
rect 6016 23908 6020 23964
rect 5956 23904 6020 23908
rect 6036 23964 6100 23968
rect 6036 23908 6040 23964
rect 6040 23908 6096 23964
rect 6096 23908 6100 23964
rect 6036 23904 6100 23908
rect 6116 23964 6180 23968
rect 6116 23908 6120 23964
rect 6120 23908 6176 23964
rect 6176 23908 6180 23964
rect 6116 23904 6180 23908
rect 6196 23964 6260 23968
rect 6196 23908 6200 23964
rect 6200 23908 6256 23964
rect 6256 23908 6260 23964
rect 6196 23904 6260 23908
rect 87100 23964 87164 23968
rect 87100 23908 87104 23964
rect 87104 23908 87160 23964
rect 87160 23908 87164 23964
rect 87100 23904 87164 23908
rect 87180 23964 87244 23968
rect 87180 23908 87184 23964
rect 87184 23908 87240 23964
rect 87240 23908 87244 23964
rect 87180 23904 87244 23908
rect 87260 23964 87324 23968
rect 87260 23908 87264 23964
rect 87264 23908 87320 23964
rect 87320 23908 87324 23964
rect 87260 23904 87324 23908
rect 87340 23964 87404 23968
rect 87340 23908 87344 23964
rect 87344 23908 87400 23964
rect 87400 23908 87404 23964
rect 87340 23904 87404 23908
rect 6692 23420 6756 23424
rect 6692 23364 6696 23420
rect 6696 23364 6752 23420
rect 6752 23364 6756 23420
rect 6692 23360 6756 23364
rect 6772 23420 6836 23424
rect 6772 23364 6776 23420
rect 6776 23364 6832 23420
rect 6832 23364 6836 23420
rect 6772 23360 6836 23364
rect 6852 23420 6916 23424
rect 6852 23364 6856 23420
rect 6856 23364 6912 23420
rect 6912 23364 6916 23420
rect 6852 23360 6916 23364
rect 6932 23420 6996 23424
rect 6932 23364 6936 23420
rect 6936 23364 6992 23420
rect 6992 23364 6996 23420
rect 6932 23360 6996 23364
rect 87836 23420 87900 23424
rect 87836 23364 87840 23420
rect 87840 23364 87896 23420
rect 87896 23364 87900 23420
rect 87836 23360 87900 23364
rect 87916 23420 87980 23424
rect 87916 23364 87920 23420
rect 87920 23364 87976 23420
rect 87976 23364 87980 23420
rect 87916 23360 87980 23364
rect 87996 23420 88060 23424
rect 87996 23364 88000 23420
rect 88000 23364 88056 23420
rect 88056 23364 88060 23420
rect 87996 23360 88060 23364
rect 88076 23420 88140 23424
rect 88076 23364 88080 23420
rect 88080 23364 88136 23420
rect 88136 23364 88140 23420
rect 88076 23360 88140 23364
rect 5956 22876 6020 22880
rect 5956 22820 5960 22876
rect 5960 22820 6016 22876
rect 6016 22820 6020 22876
rect 5956 22816 6020 22820
rect 6036 22876 6100 22880
rect 6036 22820 6040 22876
rect 6040 22820 6096 22876
rect 6096 22820 6100 22876
rect 6036 22816 6100 22820
rect 6116 22876 6180 22880
rect 6116 22820 6120 22876
rect 6120 22820 6176 22876
rect 6176 22820 6180 22876
rect 6116 22816 6180 22820
rect 6196 22876 6260 22880
rect 6196 22820 6200 22876
rect 6200 22820 6256 22876
rect 6256 22820 6260 22876
rect 6196 22816 6260 22820
rect 87100 22876 87164 22880
rect 87100 22820 87104 22876
rect 87104 22820 87160 22876
rect 87160 22820 87164 22876
rect 87100 22816 87164 22820
rect 87180 22876 87244 22880
rect 87180 22820 87184 22876
rect 87184 22820 87240 22876
rect 87240 22820 87244 22876
rect 87180 22816 87244 22820
rect 87260 22876 87324 22880
rect 87260 22820 87264 22876
rect 87264 22820 87320 22876
rect 87320 22820 87324 22876
rect 87260 22816 87324 22820
rect 87340 22876 87404 22880
rect 87340 22820 87344 22876
rect 87344 22820 87400 22876
rect 87400 22820 87404 22876
rect 87340 22816 87404 22820
rect 6692 22332 6756 22336
rect 6692 22276 6696 22332
rect 6696 22276 6752 22332
rect 6752 22276 6756 22332
rect 6692 22272 6756 22276
rect 6772 22332 6836 22336
rect 6772 22276 6776 22332
rect 6776 22276 6832 22332
rect 6832 22276 6836 22332
rect 6772 22272 6836 22276
rect 6852 22332 6916 22336
rect 6852 22276 6856 22332
rect 6856 22276 6912 22332
rect 6912 22276 6916 22332
rect 6852 22272 6916 22276
rect 6932 22332 6996 22336
rect 6932 22276 6936 22332
rect 6936 22276 6992 22332
rect 6992 22276 6996 22332
rect 6932 22272 6996 22276
rect 87836 22332 87900 22336
rect 87836 22276 87840 22332
rect 87840 22276 87896 22332
rect 87896 22276 87900 22332
rect 87836 22272 87900 22276
rect 87916 22332 87980 22336
rect 87916 22276 87920 22332
rect 87920 22276 87976 22332
rect 87976 22276 87980 22332
rect 87916 22272 87980 22276
rect 87996 22332 88060 22336
rect 87996 22276 88000 22332
rect 88000 22276 88056 22332
rect 88056 22276 88060 22332
rect 87996 22272 88060 22276
rect 88076 22332 88140 22336
rect 88076 22276 88080 22332
rect 88080 22276 88136 22332
rect 88136 22276 88140 22332
rect 88076 22272 88140 22276
rect 5956 21788 6020 21792
rect 5956 21732 5960 21788
rect 5960 21732 6016 21788
rect 6016 21732 6020 21788
rect 5956 21728 6020 21732
rect 6036 21788 6100 21792
rect 6036 21732 6040 21788
rect 6040 21732 6096 21788
rect 6096 21732 6100 21788
rect 6036 21728 6100 21732
rect 6116 21788 6180 21792
rect 6116 21732 6120 21788
rect 6120 21732 6176 21788
rect 6176 21732 6180 21788
rect 6116 21728 6180 21732
rect 6196 21788 6260 21792
rect 6196 21732 6200 21788
rect 6200 21732 6256 21788
rect 6256 21732 6260 21788
rect 6196 21728 6260 21732
rect 87100 21788 87164 21792
rect 87100 21732 87104 21788
rect 87104 21732 87160 21788
rect 87160 21732 87164 21788
rect 87100 21728 87164 21732
rect 87180 21788 87244 21792
rect 87180 21732 87184 21788
rect 87184 21732 87240 21788
rect 87240 21732 87244 21788
rect 87180 21728 87244 21732
rect 87260 21788 87324 21792
rect 87260 21732 87264 21788
rect 87264 21732 87320 21788
rect 87320 21732 87324 21788
rect 87260 21728 87324 21732
rect 87340 21788 87404 21792
rect 87340 21732 87344 21788
rect 87344 21732 87400 21788
rect 87400 21732 87404 21788
rect 87340 21728 87404 21732
rect 6692 21244 6756 21248
rect 6692 21188 6696 21244
rect 6696 21188 6752 21244
rect 6752 21188 6756 21244
rect 6692 21184 6756 21188
rect 6772 21244 6836 21248
rect 6772 21188 6776 21244
rect 6776 21188 6832 21244
rect 6832 21188 6836 21244
rect 6772 21184 6836 21188
rect 6852 21244 6916 21248
rect 6852 21188 6856 21244
rect 6856 21188 6912 21244
rect 6912 21188 6916 21244
rect 6852 21184 6916 21188
rect 6932 21244 6996 21248
rect 6932 21188 6936 21244
rect 6936 21188 6992 21244
rect 6992 21188 6996 21244
rect 6932 21184 6996 21188
rect 87836 21244 87900 21248
rect 87836 21188 87840 21244
rect 87840 21188 87896 21244
rect 87896 21188 87900 21244
rect 87836 21184 87900 21188
rect 87916 21244 87980 21248
rect 87916 21188 87920 21244
rect 87920 21188 87976 21244
rect 87976 21188 87980 21244
rect 87916 21184 87980 21188
rect 87996 21244 88060 21248
rect 87996 21188 88000 21244
rect 88000 21188 88056 21244
rect 88056 21188 88060 21244
rect 87996 21184 88060 21188
rect 88076 21244 88140 21248
rect 88076 21188 88080 21244
rect 88080 21188 88136 21244
rect 88136 21188 88140 21244
rect 88076 21184 88140 21188
rect 5956 20700 6020 20704
rect 5956 20644 5960 20700
rect 5960 20644 6016 20700
rect 6016 20644 6020 20700
rect 5956 20640 6020 20644
rect 6036 20700 6100 20704
rect 6036 20644 6040 20700
rect 6040 20644 6096 20700
rect 6096 20644 6100 20700
rect 6036 20640 6100 20644
rect 6116 20700 6180 20704
rect 6116 20644 6120 20700
rect 6120 20644 6176 20700
rect 6176 20644 6180 20700
rect 6116 20640 6180 20644
rect 6196 20700 6260 20704
rect 6196 20644 6200 20700
rect 6200 20644 6256 20700
rect 6256 20644 6260 20700
rect 6196 20640 6260 20644
rect 87100 20700 87164 20704
rect 87100 20644 87104 20700
rect 87104 20644 87160 20700
rect 87160 20644 87164 20700
rect 87100 20640 87164 20644
rect 87180 20700 87244 20704
rect 87180 20644 87184 20700
rect 87184 20644 87240 20700
rect 87240 20644 87244 20700
rect 87180 20640 87244 20644
rect 87260 20700 87324 20704
rect 87260 20644 87264 20700
rect 87264 20644 87320 20700
rect 87320 20644 87324 20700
rect 87260 20640 87324 20644
rect 87340 20700 87404 20704
rect 87340 20644 87344 20700
rect 87344 20644 87400 20700
rect 87400 20644 87404 20700
rect 87340 20640 87404 20644
rect 6692 20156 6756 20160
rect 6692 20100 6696 20156
rect 6696 20100 6752 20156
rect 6752 20100 6756 20156
rect 6692 20096 6756 20100
rect 6772 20156 6836 20160
rect 6772 20100 6776 20156
rect 6776 20100 6832 20156
rect 6832 20100 6836 20156
rect 6772 20096 6836 20100
rect 6852 20156 6916 20160
rect 6852 20100 6856 20156
rect 6856 20100 6912 20156
rect 6912 20100 6916 20156
rect 6852 20096 6916 20100
rect 6932 20156 6996 20160
rect 6932 20100 6936 20156
rect 6936 20100 6992 20156
rect 6992 20100 6996 20156
rect 6932 20096 6996 20100
rect 87836 20156 87900 20160
rect 87836 20100 87840 20156
rect 87840 20100 87896 20156
rect 87896 20100 87900 20156
rect 87836 20096 87900 20100
rect 87916 20156 87980 20160
rect 87916 20100 87920 20156
rect 87920 20100 87976 20156
rect 87976 20100 87980 20156
rect 87916 20096 87980 20100
rect 87996 20156 88060 20160
rect 87996 20100 88000 20156
rect 88000 20100 88056 20156
rect 88056 20100 88060 20156
rect 87996 20096 88060 20100
rect 88076 20156 88140 20160
rect 88076 20100 88080 20156
rect 88080 20100 88136 20156
rect 88136 20100 88140 20156
rect 88076 20096 88140 20100
rect 5956 19612 6020 19616
rect 5956 19556 5960 19612
rect 5960 19556 6016 19612
rect 6016 19556 6020 19612
rect 5956 19552 6020 19556
rect 6036 19612 6100 19616
rect 6036 19556 6040 19612
rect 6040 19556 6096 19612
rect 6096 19556 6100 19612
rect 6036 19552 6100 19556
rect 6116 19612 6180 19616
rect 6116 19556 6120 19612
rect 6120 19556 6176 19612
rect 6176 19556 6180 19612
rect 6116 19552 6180 19556
rect 6196 19612 6260 19616
rect 6196 19556 6200 19612
rect 6200 19556 6256 19612
rect 6256 19556 6260 19612
rect 6196 19552 6260 19556
rect 87100 19612 87164 19616
rect 87100 19556 87104 19612
rect 87104 19556 87160 19612
rect 87160 19556 87164 19612
rect 87100 19552 87164 19556
rect 87180 19612 87244 19616
rect 87180 19556 87184 19612
rect 87184 19556 87240 19612
rect 87240 19556 87244 19612
rect 87180 19552 87244 19556
rect 87260 19612 87324 19616
rect 87260 19556 87264 19612
rect 87264 19556 87320 19612
rect 87320 19556 87324 19612
rect 87260 19552 87324 19556
rect 87340 19612 87404 19616
rect 87340 19556 87344 19612
rect 87344 19556 87400 19612
rect 87400 19556 87404 19612
rect 87340 19552 87404 19556
rect 6692 19068 6756 19072
rect 6692 19012 6696 19068
rect 6696 19012 6752 19068
rect 6752 19012 6756 19068
rect 6692 19008 6756 19012
rect 6772 19068 6836 19072
rect 6772 19012 6776 19068
rect 6776 19012 6832 19068
rect 6832 19012 6836 19068
rect 6772 19008 6836 19012
rect 6852 19068 6916 19072
rect 6852 19012 6856 19068
rect 6856 19012 6912 19068
rect 6912 19012 6916 19068
rect 6852 19008 6916 19012
rect 6932 19068 6996 19072
rect 6932 19012 6936 19068
rect 6936 19012 6992 19068
rect 6992 19012 6996 19068
rect 6932 19008 6996 19012
rect 87836 19068 87900 19072
rect 87836 19012 87840 19068
rect 87840 19012 87896 19068
rect 87896 19012 87900 19068
rect 87836 19008 87900 19012
rect 87916 19068 87980 19072
rect 87916 19012 87920 19068
rect 87920 19012 87976 19068
rect 87976 19012 87980 19068
rect 87916 19008 87980 19012
rect 87996 19068 88060 19072
rect 87996 19012 88000 19068
rect 88000 19012 88056 19068
rect 88056 19012 88060 19068
rect 87996 19008 88060 19012
rect 88076 19068 88140 19072
rect 88076 19012 88080 19068
rect 88080 19012 88136 19068
rect 88136 19012 88140 19068
rect 88076 19008 88140 19012
rect 5956 18524 6020 18528
rect 5956 18468 5960 18524
rect 5960 18468 6016 18524
rect 6016 18468 6020 18524
rect 5956 18464 6020 18468
rect 6036 18524 6100 18528
rect 6036 18468 6040 18524
rect 6040 18468 6096 18524
rect 6096 18468 6100 18524
rect 6036 18464 6100 18468
rect 6116 18524 6180 18528
rect 6116 18468 6120 18524
rect 6120 18468 6176 18524
rect 6176 18468 6180 18524
rect 6116 18464 6180 18468
rect 6196 18524 6260 18528
rect 6196 18468 6200 18524
rect 6200 18468 6256 18524
rect 6256 18468 6260 18524
rect 6196 18464 6260 18468
rect 87100 18524 87164 18528
rect 87100 18468 87104 18524
rect 87104 18468 87160 18524
rect 87160 18468 87164 18524
rect 87100 18464 87164 18468
rect 87180 18524 87244 18528
rect 87180 18468 87184 18524
rect 87184 18468 87240 18524
rect 87240 18468 87244 18524
rect 87180 18464 87244 18468
rect 87260 18524 87324 18528
rect 87260 18468 87264 18524
rect 87264 18468 87320 18524
rect 87320 18468 87324 18524
rect 87260 18464 87324 18468
rect 87340 18524 87404 18528
rect 87340 18468 87344 18524
rect 87344 18468 87400 18524
rect 87400 18468 87404 18524
rect 87340 18464 87404 18468
rect 6692 17980 6756 17984
rect 6692 17924 6696 17980
rect 6696 17924 6752 17980
rect 6752 17924 6756 17980
rect 6692 17920 6756 17924
rect 6772 17980 6836 17984
rect 6772 17924 6776 17980
rect 6776 17924 6832 17980
rect 6832 17924 6836 17980
rect 6772 17920 6836 17924
rect 6852 17980 6916 17984
rect 6852 17924 6856 17980
rect 6856 17924 6912 17980
rect 6912 17924 6916 17980
rect 6852 17920 6916 17924
rect 6932 17980 6996 17984
rect 6932 17924 6936 17980
rect 6936 17924 6992 17980
rect 6992 17924 6996 17980
rect 6932 17920 6996 17924
rect 87836 17980 87900 17984
rect 87836 17924 87840 17980
rect 87840 17924 87896 17980
rect 87896 17924 87900 17980
rect 87836 17920 87900 17924
rect 87916 17980 87980 17984
rect 87916 17924 87920 17980
rect 87920 17924 87976 17980
rect 87976 17924 87980 17980
rect 87916 17920 87980 17924
rect 87996 17980 88060 17984
rect 87996 17924 88000 17980
rect 88000 17924 88056 17980
rect 88056 17924 88060 17980
rect 87996 17920 88060 17924
rect 88076 17980 88140 17984
rect 88076 17924 88080 17980
rect 88080 17924 88136 17980
rect 88136 17924 88140 17980
rect 88076 17920 88140 17924
rect 5956 17436 6020 17440
rect 5956 17380 5960 17436
rect 5960 17380 6016 17436
rect 6016 17380 6020 17436
rect 5956 17376 6020 17380
rect 6036 17436 6100 17440
rect 6036 17380 6040 17436
rect 6040 17380 6096 17436
rect 6096 17380 6100 17436
rect 6036 17376 6100 17380
rect 6116 17436 6180 17440
rect 6116 17380 6120 17436
rect 6120 17380 6176 17436
rect 6176 17380 6180 17436
rect 6116 17376 6180 17380
rect 6196 17436 6260 17440
rect 6196 17380 6200 17436
rect 6200 17380 6256 17436
rect 6256 17380 6260 17436
rect 6196 17376 6260 17380
rect 87100 17436 87164 17440
rect 87100 17380 87104 17436
rect 87104 17380 87160 17436
rect 87160 17380 87164 17436
rect 87100 17376 87164 17380
rect 87180 17436 87244 17440
rect 87180 17380 87184 17436
rect 87184 17380 87240 17436
rect 87240 17380 87244 17436
rect 87180 17376 87244 17380
rect 87260 17436 87324 17440
rect 87260 17380 87264 17436
rect 87264 17380 87320 17436
rect 87320 17380 87324 17436
rect 87260 17376 87324 17380
rect 87340 17436 87404 17440
rect 87340 17380 87344 17436
rect 87344 17380 87400 17436
rect 87400 17380 87404 17436
rect 87340 17376 87404 17380
rect 6692 16892 6756 16896
rect 6692 16836 6696 16892
rect 6696 16836 6752 16892
rect 6752 16836 6756 16892
rect 6692 16832 6756 16836
rect 6772 16892 6836 16896
rect 6772 16836 6776 16892
rect 6776 16836 6832 16892
rect 6832 16836 6836 16892
rect 6772 16832 6836 16836
rect 6852 16892 6916 16896
rect 6852 16836 6856 16892
rect 6856 16836 6912 16892
rect 6912 16836 6916 16892
rect 6852 16832 6916 16836
rect 6932 16892 6996 16896
rect 6932 16836 6936 16892
rect 6936 16836 6992 16892
rect 6992 16836 6996 16892
rect 6932 16832 6996 16836
rect 87836 16892 87900 16896
rect 87836 16836 87840 16892
rect 87840 16836 87896 16892
rect 87896 16836 87900 16892
rect 87836 16832 87900 16836
rect 87916 16892 87980 16896
rect 87916 16836 87920 16892
rect 87920 16836 87976 16892
rect 87976 16836 87980 16892
rect 87916 16832 87980 16836
rect 87996 16892 88060 16896
rect 87996 16836 88000 16892
rect 88000 16836 88056 16892
rect 88056 16836 88060 16892
rect 87996 16832 88060 16836
rect 88076 16892 88140 16896
rect 88076 16836 88080 16892
rect 88080 16836 88136 16892
rect 88136 16836 88140 16892
rect 88076 16832 88140 16836
rect 5956 16348 6020 16352
rect 5956 16292 5960 16348
rect 5960 16292 6016 16348
rect 6016 16292 6020 16348
rect 5956 16288 6020 16292
rect 6036 16348 6100 16352
rect 6036 16292 6040 16348
rect 6040 16292 6096 16348
rect 6096 16292 6100 16348
rect 6036 16288 6100 16292
rect 6116 16348 6180 16352
rect 6116 16292 6120 16348
rect 6120 16292 6176 16348
rect 6176 16292 6180 16348
rect 6116 16288 6180 16292
rect 6196 16348 6260 16352
rect 6196 16292 6200 16348
rect 6200 16292 6256 16348
rect 6256 16292 6260 16348
rect 6196 16288 6260 16292
rect 87100 16348 87164 16352
rect 87100 16292 87104 16348
rect 87104 16292 87160 16348
rect 87160 16292 87164 16348
rect 87100 16288 87164 16292
rect 87180 16348 87244 16352
rect 87180 16292 87184 16348
rect 87184 16292 87240 16348
rect 87240 16292 87244 16348
rect 87180 16288 87244 16292
rect 87260 16348 87324 16352
rect 87260 16292 87264 16348
rect 87264 16292 87320 16348
rect 87320 16292 87324 16348
rect 87260 16288 87324 16292
rect 87340 16348 87404 16352
rect 87340 16292 87344 16348
rect 87344 16292 87400 16348
rect 87400 16292 87404 16348
rect 87340 16288 87404 16292
rect 6692 15804 6756 15808
rect 6692 15748 6696 15804
rect 6696 15748 6752 15804
rect 6752 15748 6756 15804
rect 6692 15744 6756 15748
rect 6772 15804 6836 15808
rect 6772 15748 6776 15804
rect 6776 15748 6832 15804
rect 6832 15748 6836 15804
rect 6772 15744 6836 15748
rect 6852 15804 6916 15808
rect 6852 15748 6856 15804
rect 6856 15748 6912 15804
rect 6912 15748 6916 15804
rect 6852 15744 6916 15748
rect 6932 15804 6996 15808
rect 6932 15748 6936 15804
rect 6936 15748 6992 15804
rect 6992 15748 6996 15804
rect 6932 15744 6996 15748
rect 87836 15804 87900 15808
rect 87836 15748 87840 15804
rect 87840 15748 87896 15804
rect 87896 15748 87900 15804
rect 87836 15744 87900 15748
rect 87916 15804 87980 15808
rect 87916 15748 87920 15804
rect 87920 15748 87976 15804
rect 87976 15748 87980 15804
rect 87916 15744 87980 15748
rect 87996 15804 88060 15808
rect 87996 15748 88000 15804
rect 88000 15748 88056 15804
rect 88056 15748 88060 15804
rect 87996 15744 88060 15748
rect 88076 15804 88140 15808
rect 88076 15748 88080 15804
rect 88080 15748 88136 15804
rect 88136 15748 88140 15804
rect 88076 15744 88140 15748
rect 5956 15260 6020 15264
rect 5956 15204 5960 15260
rect 5960 15204 6016 15260
rect 6016 15204 6020 15260
rect 5956 15200 6020 15204
rect 6036 15260 6100 15264
rect 6036 15204 6040 15260
rect 6040 15204 6096 15260
rect 6096 15204 6100 15260
rect 6036 15200 6100 15204
rect 6116 15260 6180 15264
rect 6116 15204 6120 15260
rect 6120 15204 6176 15260
rect 6176 15204 6180 15260
rect 6116 15200 6180 15204
rect 6196 15260 6260 15264
rect 6196 15204 6200 15260
rect 6200 15204 6256 15260
rect 6256 15204 6260 15260
rect 6196 15200 6260 15204
rect 87100 15260 87164 15264
rect 87100 15204 87104 15260
rect 87104 15204 87160 15260
rect 87160 15204 87164 15260
rect 87100 15200 87164 15204
rect 87180 15260 87244 15264
rect 87180 15204 87184 15260
rect 87184 15204 87240 15260
rect 87240 15204 87244 15260
rect 87180 15200 87244 15204
rect 87260 15260 87324 15264
rect 87260 15204 87264 15260
rect 87264 15204 87320 15260
rect 87320 15204 87324 15260
rect 87260 15200 87324 15204
rect 87340 15260 87404 15264
rect 87340 15204 87344 15260
rect 87344 15204 87400 15260
rect 87400 15204 87404 15260
rect 87340 15200 87404 15204
rect 6692 14716 6756 14720
rect 6692 14660 6696 14716
rect 6696 14660 6752 14716
rect 6752 14660 6756 14716
rect 6692 14656 6756 14660
rect 6772 14716 6836 14720
rect 6772 14660 6776 14716
rect 6776 14660 6832 14716
rect 6832 14660 6836 14716
rect 6772 14656 6836 14660
rect 6852 14716 6916 14720
rect 6852 14660 6856 14716
rect 6856 14660 6912 14716
rect 6912 14660 6916 14716
rect 6852 14656 6916 14660
rect 6932 14716 6996 14720
rect 6932 14660 6936 14716
rect 6936 14660 6992 14716
rect 6992 14660 6996 14716
rect 6932 14656 6996 14660
rect 87836 14716 87900 14720
rect 87836 14660 87840 14716
rect 87840 14660 87896 14716
rect 87896 14660 87900 14716
rect 87836 14656 87900 14660
rect 87916 14716 87980 14720
rect 87916 14660 87920 14716
rect 87920 14660 87976 14716
rect 87976 14660 87980 14716
rect 87916 14656 87980 14660
rect 87996 14716 88060 14720
rect 87996 14660 88000 14716
rect 88000 14660 88056 14716
rect 88056 14660 88060 14716
rect 87996 14656 88060 14660
rect 88076 14716 88140 14720
rect 88076 14660 88080 14716
rect 88080 14660 88136 14716
rect 88136 14660 88140 14716
rect 88076 14656 88140 14660
rect 5956 14172 6020 14176
rect 5956 14116 5960 14172
rect 5960 14116 6016 14172
rect 6016 14116 6020 14172
rect 5956 14112 6020 14116
rect 6036 14172 6100 14176
rect 6036 14116 6040 14172
rect 6040 14116 6096 14172
rect 6096 14116 6100 14172
rect 6036 14112 6100 14116
rect 6116 14172 6180 14176
rect 6116 14116 6120 14172
rect 6120 14116 6176 14172
rect 6176 14116 6180 14172
rect 6116 14112 6180 14116
rect 6196 14172 6260 14176
rect 6196 14116 6200 14172
rect 6200 14116 6256 14172
rect 6256 14116 6260 14172
rect 6196 14112 6260 14116
rect 87100 14172 87164 14176
rect 87100 14116 87104 14172
rect 87104 14116 87160 14172
rect 87160 14116 87164 14172
rect 87100 14112 87164 14116
rect 87180 14172 87244 14176
rect 87180 14116 87184 14172
rect 87184 14116 87240 14172
rect 87240 14116 87244 14172
rect 87180 14112 87244 14116
rect 87260 14172 87324 14176
rect 87260 14116 87264 14172
rect 87264 14116 87320 14172
rect 87320 14116 87324 14172
rect 87260 14112 87324 14116
rect 87340 14172 87404 14176
rect 87340 14116 87344 14172
rect 87344 14116 87400 14172
rect 87400 14116 87404 14172
rect 87340 14112 87404 14116
rect 6692 13628 6756 13632
rect 6692 13572 6696 13628
rect 6696 13572 6752 13628
rect 6752 13572 6756 13628
rect 6692 13568 6756 13572
rect 6772 13628 6836 13632
rect 6772 13572 6776 13628
rect 6776 13572 6832 13628
rect 6832 13572 6836 13628
rect 6772 13568 6836 13572
rect 6852 13628 6916 13632
rect 6852 13572 6856 13628
rect 6856 13572 6912 13628
rect 6912 13572 6916 13628
rect 6852 13568 6916 13572
rect 6932 13628 6996 13632
rect 6932 13572 6936 13628
rect 6936 13572 6992 13628
rect 6992 13572 6996 13628
rect 6932 13568 6996 13572
rect 87836 13628 87900 13632
rect 87836 13572 87840 13628
rect 87840 13572 87896 13628
rect 87896 13572 87900 13628
rect 87836 13568 87900 13572
rect 87916 13628 87980 13632
rect 87916 13572 87920 13628
rect 87920 13572 87976 13628
rect 87976 13572 87980 13628
rect 87916 13568 87980 13572
rect 87996 13628 88060 13632
rect 87996 13572 88000 13628
rect 88000 13572 88056 13628
rect 88056 13572 88060 13628
rect 87996 13568 88060 13572
rect 88076 13628 88140 13632
rect 88076 13572 88080 13628
rect 88080 13572 88136 13628
rect 88136 13572 88140 13628
rect 88076 13568 88140 13572
rect 5956 13084 6020 13088
rect 5956 13028 5960 13084
rect 5960 13028 6016 13084
rect 6016 13028 6020 13084
rect 5956 13024 6020 13028
rect 6036 13084 6100 13088
rect 6036 13028 6040 13084
rect 6040 13028 6096 13084
rect 6096 13028 6100 13084
rect 6036 13024 6100 13028
rect 6116 13084 6180 13088
rect 6116 13028 6120 13084
rect 6120 13028 6176 13084
rect 6176 13028 6180 13084
rect 6116 13024 6180 13028
rect 6196 13084 6260 13088
rect 6196 13028 6200 13084
rect 6200 13028 6256 13084
rect 6256 13028 6260 13084
rect 6196 13024 6260 13028
rect 87100 13084 87164 13088
rect 87100 13028 87104 13084
rect 87104 13028 87160 13084
rect 87160 13028 87164 13084
rect 87100 13024 87164 13028
rect 87180 13084 87244 13088
rect 87180 13028 87184 13084
rect 87184 13028 87240 13084
rect 87240 13028 87244 13084
rect 87180 13024 87244 13028
rect 87260 13084 87324 13088
rect 87260 13028 87264 13084
rect 87264 13028 87320 13084
rect 87320 13028 87324 13084
rect 87260 13024 87324 13028
rect 87340 13084 87404 13088
rect 87340 13028 87344 13084
rect 87344 13028 87400 13084
rect 87400 13028 87404 13084
rect 87340 13024 87404 13028
rect 6692 12540 6756 12544
rect 6692 12484 6696 12540
rect 6696 12484 6752 12540
rect 6752 12484 6756 12540
rect 6692 12480 6756 12484
rect 6772 12540 6836 12544
rect 6772 12484 6776 12540
rect 6776 12484 6832 12540
rect 6832 12484 6836 12540
rect 6772 12480 6836 12484
rect 6852 12540 6916 12544
rect 6852 12484 6856 12540
rect 6856 12484 6912 12540
rect 6912 12484 6916 12540
rect 6852 12480 6916 12484
rect 6932 12540 6996 12544
rect 6932 12484 6936 12540
rect 6936 12484 6992 12540
rect 6992 12484 6996 12540
rect 6932 12480 6996 12484
rect 87836 12540 87900 12544
rect 87836 12484 87840 12540
rect 87840 12484 87896 12540
rect 87896 12484 87900 12540
rect 87836 12480 87900 12484
rect 87916 12540 87980 12544
rect 87916 12484 87920 12540
rect 87920 12484 87976 12540
rect 87976 12484 87980 12540
rect 87916 12480 87980 12484
rect 87996 12540 88060 12544
rect 87996 12484 88000 12540
rect 88000 12484 88056 12540
rect 88056 12484 88060 12540
rect 87996 12480 88060 12484
rect 88076 12540 88140 12544
rect 88076 12484 88080 12540
rect 88080 12484 88136 12540
rect 88136 12484 88140 12540
rect 88076 12480 88140 12484
rect 5956 11996 6020 12000
rect 5956 11940 5960 11996
rect 5960 11940 6016 11996
rect 6016 11940 6020 11996
rect 5956 11936 6020 11940
rect 6036 11996 6100 12000
rect 6036 11940 6040 11996
rect 6040 11940 6096 11996
rect 6096 11940 6100 11996
rect 6036 11936 6100 11940
rect 6116 11996 6180 12000
rect 6116 11940 6120 11996
rect 6120 11940 6176 11996
rect 6176 11940 6180 11996
rect 6116 11936 6180 11940
rect 6196 11996 6260 12000
rect 6196 11940 6200 11996
rect 6200 11940 6256 11996
rect 6256 11940 6260 11996
rect 6196 11936 6260 11940
rect 87100 11996 87164 12000
rect 87100 11940 87104 11996
rect 87104 11940 87160 11996
rect 87160 11940 87164 11996
rect 87100 11936 87164 11940
rect 87180 11996 87244 12000
rect 87180 11940 87184 11996
rect 87184 11940 87240 11996
rect 87240 11940 87244 11996
rect 87180 11936 87244 11940
rect 87260 11996 87324 12000
rect 87260 11940 87264 11996
rect 87264 11940 87320 11996
rect 87320 11940 87324 11996
rect 87260 11936 87324 11940
rect 87340 11996 87404 12000
rect 87340 11940 87344 11996
rect 87344 11940 87400 11996
rect 87400 11940 87404 11996
rect 87340 11936 87404 11940
rect 6692 11452 6756 11456
rect 6692 11396 6696 11452
rect 6696 11396 6752 11452
rect 6752 11396 6756 11452
rect 6692 11392 6756 11396
rect 6772 11452 6836 11456
rect 6772 11396 6776 11452
rect 6776 11396 6832 11452
rect 6832 11396 6836 11452
rect 6772 11392 6836 11396
rect 6852 11452 6916 11456
rect 6852 11396 6856 11452
rect 6856 11396 6912 11452
rect 6912 11396 6916 11452
rect 6852 11392 6916 11396
rect 6932 11452 6996 11456
rect 6932 11396 6936 11452
rect 6936 11396 6992 11452
rect 6992 11396 6996 11452
rect 6932 11392 6996 11396
rect 87836 11452 87900 11456
rect 87836 11396 87840 11452
rect 87840 11396 87896 11452
rect 87896 11396 87900 11452
rect 87836 11392 87900 11396
rect 87916 11452 87980 11456
rect 87916 11396 87920 11452
rect 87920 11396 87976 11452
rect 87976 11396 87980 11452
rect 87916 11392 87980 11396
rect 87996 11452 88060 11456
rect 87996 11396 88000 11452
rect 88000 11396 88056 11452
rect 88056 11396 88060 11452
rect 87996 11392 88060 11396
rect 88076 11452 88140 11456
rect 88076 11396 88080 11452
rect 88080 11396 88136 11452
rect 88136 11396 88140 11452
rect 88076 11392 88140 11396
rect 5956 10908 6020 10912
rect 5956 10852 5960 10908
rect 5960 10852 6016 10908
rect 6016 10852 6020 10908
rect 5956 10848 6020 10852
rect 6036 10908 6100 10912
rect 6036 10852 6040 10908
rect 6040 10852 6096 10908
rect 6096 10852 6100 10908
rect 6036 10848 6100 10852
rect 6116 10908 6180 10912
rect 6116 10852 6120 10908
rect 6120 10852 6176 10908
rect 6176 10852 6180 10908
rect 6116 10848 6180 10852
rect 6196 10908 6260 10912
rect 6196 10852 6200 10908
rect 6200 10852 6256 10908
rect 6256 10852 6260 10908
rect 6196 10848 6260 10852
rect 87100 10908 87164 10912
rect 87100 10852 87104 10908
rect 87104 10852 87160 10908
rect 87160 10852 87164 10908
rect 87100 10848 87164 10852
rect 87180 10908 87244 10912
rect 87180 10852 87184 10908
rect 87184 10852 87240 10908
rect 87240 10852 87244 10908
rect 87180 10848 87244 10852
rect 87260 10908 87324 10912
rect 87260 10852 87264 10908
rect 87264 10852 87320 10908
rect 87320 10852 87324 10908
rect 87260 10848 87324 10852
rect 87340 10908 87404 10912
rect 87340 10852 87344 10908
rect 87344 10852 87400 10908
rect 87400 10852 87404 10908
rect 87340 10848 87404 10852
rect 6692 10364 6756 10368
rect 6692 10308 6696 10364
rect 6696 10308 6752 10364
rect 6752 10308 6756 10364
rect 6692 10304 6756 10308
rect 6772 10364 6836 10368
rect 6772 10308 6776 10364
rect 6776 10308 6832 10364
rect 6832 10308 6836 10364
rect 6772 10304 6836 10308
rect 6852 10364 6916 10368
rect 6852 10308 6856 10364
rect 6856 10308 6912 10364
rect 6912 10308 6916 10364
rect 6852 10304 6916 10308
rect 6932 10364 6996 10368
rect 6932 10308 6936 10364
rect 6936 10308 6992 10364
rect 6992 10308 6996 10364
rect 6932 10304 6996 10308
rect 87836 10364 87900 10368
rect 87836 10308 87840 10364
rect 87840 10308 87896 10364
rect 87896 10308 87900 10364
rect 87836 10304 87900 10308
rect 87916 10364 87980 10368
rect 87916 10308 87920 10364
rect 87920 10308 87976 10364
rect 87976 10308 87980 10364
rect 87916 10304 87980 10308
rect 87996 10364 88060 10368
rect 87996 10308 88000 10364
rect 88000 10308 88056 10364
rect 88056 10308 88060 10364
rect 87996 10304 88060 10308
rect 88076 10364 88140 10368
rect 88076 10308 88080 10364
rect 88080 10308 88136 10364
rect 88136 10308 88140 10364
rect 88076 10304 88140 10308
rect 5956 9820 6020 9824
rect 5956 9764 5960 9820
rect 5960 9764 6016 9820
rect 6016 9764 6020 9820
rect 5956 9760 6020 9764
rect 6036 9820 6100 9824
rect 6036 9764 6040 9820
rect 6040 9764 6096 9820
rect 6096 9764 6100 9820
rect 6036 9760 6100 9764
rect 6116 9820 6180 9824
rect 6116 9764 6120 9820
rect 6120 9764 6176 9820
rect 6176 9764 6180 9820
rect 6116 9760 6180 9764
rect 6196 9820 6260 9824
rect 6196 9764 6200 9820
rect 6200 9764 6256 9820
rect 6256 9764 6260 9820
rect 6196 9760 6260 9764
rect 87100 9820 87164 9824
rect 87100 9764 87104 9820
rect 87104 9764 87160 9820
rect 87160 9764 87164 9820
rect 87100 9760 87164 9764
rect 87180 9820 87244 9824
rect 87180 9764 87184 9820
rect 87184 9764 87240 9820
rect 87240 9764 87244 9820
rect 87180 9760 87244 9764
rect 87260 9820 87324 9824
rect 87260 9764 87264 9820
rect 87264 9764 87320 9820
rect 87320 9764 87324 9820
rect 87260 9760 87324 9764
rect 87340 9820 87404 9824
rect 87340 9764 87344 9820
rect 87344 9764 87400 9820
rect 87400 9764 87404 9820
rect 87340 9760 87404 9764
rect 6692 9276 6756 9280
rect 6692 9220 6696 9276
rect 6696 9220 6752 9276
rect 6752 9220 6756 9276
rect 6692 9216 6756 9220
rect 6772 9276 6836 9280
rect 6772 9220 6776 9276
rect 6776 9220 6832 9276
rect 6832 9220 6836 9276
rect 6772 9216 6836 9220
rect 6852 9276 6916 9280
rect 6852 9220 6856 9276
rect 6856 9220 6912 9276
rect 6912 9220 6916 9276
rect 6852 9216 6916 9220
rect 6932 9276 6996 9280
rect 6932 9220 6936 9276
rect 6936 9220 6992 9276
rect 6992 9220 6996 9276
rect 6932 9216 6996 9220
rect 87836 9276 87900 9280
rect 87836 9220 87840 9276
rect 87840 9220 87896 9276
rect 87896 9220 87900 9276
rect 87836 9216 87900 9220
rect 87916 9276 87980 9280
rect 87916 9220 87920 9276
rect 87920 9220 87976 9276
rect 87976 9220 87980 9276
rect 87916 9216 87980 9220
rect 87996 9276 88060 9280
rect 87996 9220 88000 9276
rect 88000 9220 88056 9276
rect 88056 9220 88060 9276
rect 87996 9216 88060 9220
rect 88076 9276 88140 9280
rect 88076 9220 88080 9276
rect 88080 9220 88136 9276
rect 88136 9220 88140 9276
rect 88076 9216 88140 9220
rect 5956 8732 6020 8736
rect 5956 8676 5960 8732
rect 5960 8676 6016 8732
rect 6016 8676 6020 8732
rect 5956 8672 6020 8676
rect 6036 8732 6100 8736
rect 6036 8676 6040 8732
rect 6040 8676 6096 8732
rect 6096 8676 6100 8732
rect 6036 8672 6100 8676
rect 6116 8732 6180 8736
rect 6116 8676 6120 8732
rect 6120 8676 6176 8732
rect 6176 8676 6180 8732
rect 6116 8672 6180 8676
rect 6196 8732 6260 8736
rect 6196 8676 6200 8732
rect 6200 8676 6256 8732
rect 6256 8676 6260 8732
rect 6196 8672 6260 8676
rect 87100 8732 87164 8736
rect 87100 8676 87104 8732
rect 87104 8676 87160 8732
rect 87160 8676 87164 8732
rect 87100 8672 87164 8676
rect 87180 8732 87244 8736
rect 87180 8676 87184 8732
rect 87184 8676 87240 8732
rect 87240 8676 87244 8732
rect 87180 8672 87244 8676
rect 87260 8732 87324 8736
rect 87260 8676 87264 8732
rect 87264 8676 87320 8732
rect 87320 8676 87324 8732
rect 87260 8672 87324 8676
rect 87340 8732 87404 8736
rect 87340 8676 87344 8732
rect 87344 8676 87400 8732
rect 87400 8676 87404 8732
rect 87340 8672 87404 8676
rect 6692 8188 6756 8192
rect 6692 8132 6696 8188
rect 6696 8132 6752 8188
rect 6752 8132 6756 8188
rect 6692 8128 6756 8132
rect 6772 8188 6836 8192
rect 6772 8132 6776 8188
rect 6776 8132 6832 8188
rect 6832 8132 6836 8188
rect 6772 8128 6836 8132
rect 6852 8188 6916 8192
rect 6852 8132 6856 8188
rect 6856 8132 6912 8188
rect 6912 8132 6916 8188
rect 6852 8128 6916 8132
rect 6932 8188 6996 8192
rect 6932 8132 6936 8188
rect 6936 8132 6992 8188
rect 6992 8132 6996 8188
rect 6932 8128 6996 8132
rect 87836 8188 87900 8192
rect 87836 8132 87840 8188
rect 87840 8132 87896 8188
rect 87896 8132 87900 8188
rect 87836 8128 87900 8132
rect 87916 8188 87980 8192
rect 87916 8132 87920 8188
rect 87920 8132 87976 8188
rect 87976 8132 87980 8188
rect 87916 8128 87980 8132
rect 87996 8188 88060 8192
rect 87996 8132 88000 8188
rect 88000 8132 88056 8188
rect 88056 8132 88060 8188
rect 87996 8128 88060 8132
rect 88076 8188 88140 8192
rect 88076 8132 88080 8188
rect 88080 8132 88136 8188
rect 88136 8132 88140 8188
rect 88076 8128 88140 8132
rect 5956 7644 6020 7648
rect 5956 7588 5960 7644
rect 5960 7588 6016 7644
rect 6016 7588 6020 7644
rect 5956 7584 6020 7588
rect 6036 7644 6100 7648
rect 6036 7588 6040 7644
rect 6040 7588 6096 7644
rect 6096 7588 6100 7644
rect 6036 7584 6100 7588
rect 6116 7644 6180 7648
rect 6116 7588 6120 7644
rect 6120 7588 6176 7644
rect 6176 7588 6180 7644
rect 6116 7584 6180 7588
rect 6196 7644 6260 7648
rect 6196 7588 6200 7644
rect 6200 7588 6256 7644
rect 6256 7588 6260 7644
rect 6196 7584 6260 7588
rect 18724 7644 18788 7648
rect 18724 7588 18728 7644
rect 18728 7588 18784 7644
rect 18784 7588 18788 7644
rect 18724 7584 18788 7588
rect 18804 7644 18868 7648
rect 18804 7588 18808 7644
rect 18808 7588 18864 7644
rect 18864 7588 18868 7644
rect 18804 7584 18868 7588
rect 18884 7644 18948 7648
rect 18884 7588 18888 7644
rect 18888 7588 18944 7644
rect 18944 7588 18948 7644
rect 18884 7584 18948 7588
rect 18964 7644 19028 7648
rect 18964 7588 18968 7644
rect 18968 7588 19024 7644
rect 19024 7588 19028 7644
rect 18964 7584 19028 7588
rect 37724 7644 37788 7648
rect 37724 7588 37728 7644
rect 37728 7588 37784 7644
rect 37784 7588 37788 7644
rect 37724 7584 37788 7588
rect 37804 7644 37868 7648
rect 37804 7588 37808 7644
rect 37808 7588 37864 7644
rect 37864 7588 37868 7644
rect 37804 7584 37868 7588
rect 37884 7644 37948 7648
rect 37884 7588 37888 7644
rect 37888 7588 37944 7644
rect 37944 7588 37948 7644
rect 37884 7584 37948 7588
rect 37964 7644 38028 7648
rect 37964 7588 37968 7644
rect 37968 7588 38024 7644
rect 38024 7588 38028 7644
rect 37964 7584 38028 7588
rect 56724 7644 56788 7648
rect 56724 7588 56728 7644
rect 56728 7588 56784 7644
rect 56784 7588 56788 7644
rect 56724 7584 56788 7588
rect 56804 7644 56868 7648
rect 56804 7588 56808 7644
rect 56808 7588 56864 7644
rect 56864 7588 56868 7644
rect 56804 7584 56868 7588
rect 56884 7644 56948 7648
rect 56884 7588 56888 7644
rect 56888 7588 56944 7644
rect 56944 7588 56948 7644
rect 56884 7584 56948 7588
rect 56964 7644 57028 7648
rect 56964 7588 56968 7644
rect 56968 7588 57024 7644
rect 57024 7588 57028 7644
rect 56964 7584 57028 7588
rect 75724 7644 75788 7648
rect 75724 7588 75728 7644
rect 75728 7588 75784 7644
rect 75784 7588 75788 7644
rect 75724 7584 75788 7588
rect 75804 7644 75868 7648
rect 75804 7588 75808 7644
rect 75808 7588 75864 7644
rect 75864 7588 75868 7644
rect 75804 7584 75868 7588
rect 75884 7644 75948 7648
rect 75884 7588 75888 7644
rect 75888 7588 75944 7644
rect 75944 7588 75948 7644
rect 75884 7584 75948 7588
rect 75964 7644 76028 7648
rect 75964 7588 75968 7644
rect 75968 7588 76024 7644
rect 76024 7588 76028 7644
rect 75964 7584 76028 7588
rect 87100 7644 87164 7648
rect 87100 7588 87104 7644
rect 87104 7588 87160 7644
rect 87160 7588 87164 7644
rect 87100 7584 87164 7588
rect 87180 7644 87244 7648
rect 87180 7588 87184 7644
rect 87184 7588 87240 7644
rect 87240 7588 87244 7644
rect 87180 7584 87244 7588
rect 87260 7644 87324 7648
rect 87260 7588 87264 7644
rect 87264 7588 87320 7644
rect 87320 7588 87324 7644
rect 87260 7584 87324 7588
rect 87340 7644 87404 7648
rect 87340 7588 87344 7644
rect 87344 7588 87400 7644
rect 87400 7588 87404 7644
rect 87340 7584 87404 7588
rect 6692 7100 6756 7104
rect 6692 7044 6696 7100
rect 6696 7044 6752 7100
rect 6752 7044 6756 7100
rect 6692 7040 6756 7044
rect 6772 7100 6836 7104
rect 6772 7044 6776 7100
rect 6776 7044 6832 7100
rect 6832 7044 6836 7100
rect 6772 7040 6836 7044
rect 6852 7100 6916 7104
rect 6852 7044 6856 7100
rect 6856 7044 6912 7100
rect 6912 7044 6916 7100
rect 6852 7040 6916 7044
rect 6932 7100 6996 7104
rect 6932 7044 6936 7100
rect 6936 7044 6992 7100
rect 6992 7044 6996 7100
rect 6932 7040 6996 7044
rect 19384 7100 19448 7104
rect 19384 7044 19388 7100
rect 19388 7044 19444 7100
rect 19444 7044 19448 7100
rect 19384 7040 19448 7044
rect 19464 7100 19528 7104
rect 19464 7044 19468 7100
rect 19468 7044 19524 7100
rect 19524 7044 19528 7100
rect 19464 7040 19528 7044
rect 19544 7100 19608 7104
rect 19544 7044 19548 7100
rect 19548 7044 19604 7100
rect 19604 7044 19608 7100
rect 19544 7040 19608 7044
rect 19624 7100 19688 7104
rect 19624 7044 19628 7100
rect 19628 7044 19684 7100
rect 19684 7044 19688 7100
rect 19624 7040 19688 7044
rect 38384 7100 38448 7104
rect 38384 7044 38388 7100
rect 38388 7044 38444 7100
rect 38444 7044 38448 7100
rect 38384 7040 38448 7044
rect 38464 7100 38528 7104
rect 38464 7044 38468 7100
rect 38468 7044 38524 7100
rect 38524 7044 38528 7100
rect 38464 7040 38528 7044
rect 38544 7100 38608 7104
rect 38544 7044 38548 7100
rect 38548 7044 38604 7100
rect 38604 7044 38608 7100
rect 38544 7040 38608 7044
rect 38624 7100 38688 7104
rect 38624 7044 38628 7100
rect 38628 7044 38684 7100
rect 38684 7044 38688 7100
rect 38624 7040 38688 7044
rect 57384 7100 57448 7104
rect 57384 7044 57388 7100
rect 57388 7044 57444 7100
rect 57444 7044 57448 7100
rect 57384 7040 57448 7044
rect 57464 7100 57528 7104
rect 57464 7044 57468 7100
rect 57468 7044 57524 7100
rect 57524 7044 57528 7100
rect 57464 7040 57528 7044
rect 57544 7100 57608 7104
rect 57544 7044 57548 7100
rect 57548 7044 57604 7100
rect 57604 7044 57608 7100
rect 57544 7040 57608 7044
rect 57624 7100 57688 7104
rect 57624 7044 57628 7100
rect 57628 7044 57684 7100
rect 57684 7044 57688 7100
rect 57624 7040 57688 7044
rect 76384 7100 76448 7104
rect 76384 7044 76388 7100
rect 76388 7044 76444 7100
rect 76444 7044 76448 7100
rect 76384 7040 76448 7044
rect 76464 7100 76528 7104
rect 76464 7044 76468 7100
rect 76468 7044 76524 7100
rect 76524 7044 76528 7100
rect 76464 7040 76528 7044
rect 76544 7100 76608 7104
rect 76544 7044 76548 7100
rect 76548 7044 76604 7100
rect 76604 7044 76608 7100
rect 76544 7040 76608 7044
rect 76624 7100 76688 7104
rect 76624 7044 76628 7100
rect 76628 7044 76684 7100
rect 76684 7044 76688 7100
rect 76624 7040 76688 7044
rect 87836 7100 87900 7104
rect 87836 7044 87840 7100
rect 87840 7044 87896 7100
rect 87896 7044 87900 7100
rect 87836 7040 87900 7044
rect 87916 7100 87980 7104
rect 87916 7044 87920 7100
rect 87920 7044 87976 7100
rect 87976 7044 87980 7100
rect 87916 7040 87980 7044
rect 87996 7100 88060 7104
rect 87996 7044 88000 7100
rect 88000 7044 88056 7100
rect 88056 7044 88060 7100
rect 87996 7040 88060 7044
rect 88076 7100 88140 7104
rect 88076 7044 88080 7100
rect 88080 7044 88136 7100
rect 88136 7044 88140 7100
rect 88076 7040 88140 7044
rect 18724 6556 18788 6560
rect 18724 6500 18728 6556
rect 18728 6500 18784 6556
rect 18784 6500 18788 6556
rect 18724 6496 18788 6500
rect 18804 6556 18868 6560
rect 18804 6500 18808 6556
rect 18808 6500 18864 6556
rect 18864 6500 18868 6556
rect 18804 6496 18868 6500
rect 18884 6556 18948 6560
rect 18884 6500 18888 6556
rect 18888 6500 18944 6556
rect 18944 6500 18948 6556
rect 18884 6496 18948 6500
rect 18964 6556 19028 6560
rect 18964 6500 18968 6556
rect 18968 6500 19024 6556
rect 19024 6500 19028 6556
rect 18964 6496 19028 6500
rect 37724 6556 37788 6560
rect 37724 6500 37728 6556
rect 37728 6500 37784 6556
rect 37784 6500 37788 6556
rect 37724 6496 37788 6500
rect 37804 6556 37868 6560
rect 37804 6500 37808 6556
rect 37808 6500 37864 6556
rect 37864 6500 37868 6556
rect 37804 6496 37868 6500
rect 37884 6556 37948 6560
rect 37884 6500 37888 6556
rect 37888 6500 37944 6556
rect 37944 6500 37948 6556
rect 37884 6496 37948 6500
rect 37964 6556 38028 6560
rect 37964 6500 37968 6556
rect 37968 6500 38024 6556
rect 38024 6500 38028 6556
rect 37964 6496 38028 6500
rect 56724 6556 56788 6560
rect 56724 6500 56728 6556
rect 56728 6500 56784 6556
rect 56784 6500 56788 6556
rect 56724 6496 56788 6500
rect 56804 6556 56868 6560
rect 56804 6500 56808 6556
rect 56808 6500 56864 6556
rect 56864 6500 56868 6556
rect 56804 6496 56868 6500
rect 56884 6556 56948 6560
rect 56884 6500 56888 6556
rect 56888 6500 56944 6556
rect 56944 6500 56948 6556
rect 56884 6496 56948 6500
rect 56964 6556 57028 6560
rect 56964 6500 56968 6556
rect 56968 6500 57024 6556
rect 57024 6500 57028 6556
rect 56964 6496 57028 6500
rect 75724 6556 75788 6560
rect 75724 6500 75728 6556
rect 75728 6500 75784 6556
rect 75784 6500 75788 6556
rect 75724 6496 75788 6500
rect 75804 6556 75868 6560
rect 75804 6500 75808 6556
rect 75808 6500 75864 6556
rect 75864 6500 75868 6556
rect 75804 6496 75868 6500
rect 75884 6556 75948 6560
rect 75884 6500 75888 6556
rect 75888 6500 75944 6556
rect 75944 6500 75948 6556
rect 75884 6496 75948 6500
rect 75964 6556 76028 6560
rect 75964 6500 75968 6556
rect 75968 6500 76024 6556
rect 76024 6500 76028 6556
rect 75964 6496 76028 6500
rect 19384 6012 19448 6016
rect 19384 5956 19388 6012
rect 19388 5956 19444 6012
rect 19444 5956 19448 6012
rect 19384 5952 19448 5956
rect 19464 6012 19528 6016
rect 19464 5956 19468 6012
rect 19468 5956 19524 6012
rect 19524 5956 19528 6012
rect 19464 5952 19528 5956
rect 19544 6012 19608 6016
rect 19544 5956 19548 6012
rect 19548 5956 19604 6012
rect 19604 5956 19608 6012
rect 19544 5952 19608 5956
rect 19624 6012 19688 6016
rect 19624 5956 19628 6012
rect 19628 5956 19684 6012
rect 19684 5956 19688 6012
rect 19624 5952 19688 5956
rect 38384 6012 38448 6016
rect 38384 5956 38388 6012
rect 38388 5956 38444 6012
rect 38444 5956 38448 6012
rect 38384 5952 38448 5956
rect 38464 6012 38528 6016
rect 38464 5956 38468 6012
rect 38468 5956 38524 6012
rect 38524 5956 38528 6012
rect 38464 5952 38528 5956
rect 38544 6012 38608 6016
rect 38544 5956 38548 6012
rect 38548 5956 38604 6012
rect 38604 5956 38608 6012
rect 38544 5952 38608 5956
rect 38624 6012 38688 6016
rect 38624 5956 38628 6012
rect 38628 5956 38684 6012
rect 38684 5956 38688 6012
rect 38624 5952 38688 5956
rect 57384 6012 57448 6016
rect 57384 5956 57388 6012
rect 57388 5956 57444 6012
rect 57444 5956 57448 6012
rect 57384 5952 57448 5956
rect 57464 6012 57528 6016
rect 57464 5956 57468 6012
rect 57468 5956 57524 6012
rect 57524 5956 57528 6012
rect 57464 5952 57528 5956
rect 57544 6012 57608 6016
rect 57544 5956 57548 6012
rect 57548 5956 57604 6012
rect 57604 5956 57608 6012
rect 57544 5952 57608 5956
rect 57624 6012 57688 6016
rect 57624 5956 57628 6012
rect 57628 5956 57684 6012
rect 57684 5956 57688 6012
rect 57624 5952 57688 5956
rect 76384 6012 76448 6016
rect 76384 5956 76388 6012
rect 76388 5956 76444 6012
rect 76444 5956 76448 6012
rect 76384 5952 76448 5956
rect 76464 6012 76528 6016
rect 76464 5956 76468 6012
rect 76468 5956 76524 6012
rect 76524 5956 76528 6012
rect 76464 5952 76528 5956
rect 76544 6012 76608 6016
rect 76544 5956 76548 6012
rect 76548 5956 76604 6012
rect 76604 5956 76608 6012
rect 76544 5952 76608 5956
rect 76624 6012 76688 6016
rect 76624 5956 76628 6012
rect 76628 5956 76684 6012
rect 76684 5956 76688 6012
rect 76624 5952 76688 5956
rect 18724 5468 18788 5472
rect 18724 5412 18728 5468
rect 18728 5412 18784 5468
rect 18784 5412 18788 5468
rect 18724 5408 18788 5412
rect 18804 5468 18868 5472
rect 18804 5412 18808 5468
rect 18808 5412 18864 5468
rect 18864 5412 18868 5468
rect 18804 5408 18868 5412
rect 18884 5468 18948 5472
rect 18884 5412 18888 5468
rect 18888 5412 18944 5468
rect 18944 5412 18948 5468
rect 18884 5408 18948 5412
rect 18964 5468 19028 5472
rect 18964 5412 18968 5468
rect 18968 5412 19024 5468
rect 19024 5412 19028 5468
rect 18964 5408 19028 5412
rect 37724 5468 37788 5472
rect 37724 5412 37728 5468
rect 37728 5412 37784 5468
rect 37784 5412 37788 5468
rect 37724 5408 37788 5412
rect 37804 5468 37868 5472
rect 37804 5412 37808 5468
rect 37808 5412 37864 5468
rect 37864 5412 37868 5468
rect 37804 5408 37868 5412
rect 37884 5468 37948 5472
rect 37884 5412 37888 5468
rect 37888 5412 37944 5468
rect 37944 5412 37948 5468
rect 37884 5408 37948 5412
rect 37964 5468 38028 5472
rect 37964 5412 37968 5468
rect 37968 5412 38024 5468
rect 38024 5412 38028 5468
rect 37964 5408 38028 5412
rect 56724 5468 56788 5472
rect 56724 5412 56728 5468
rect 56728 5412 56784 5468
rect 56784 5412 56788 5468
rect 56724 5408 56788 5412
rect 56804 5468 56868 5472
rect 56804 5412 56808 5468
rect 56808 5412 56864 5468
rect 56864 5412 56868 5468
rect 56804 5408 56868 5412
rect 56884 5468 56948 5472
rect 56884 5412 56888 5468
rect 56888 5412 56944 5468
rect 56944 5412 56948 5468
rect 56884 5408 56948 5412
rect 56964 5468 57028 5472
rect 56964 5412 56968 5468
rect 56968 5412 57024 5468
rect 57024 5412 57028 5468
rect 56964 5408 57028 5412
rect 75724 5468 75788 5472
rect 75724 5412 75728 5468
rect 75728 5412 75784 5468
rect 75784 5412 75788 5468
rect 75724 5408 75788 5412
rect 75804 5468 75868 5472
rect 75804 5412 75808 5468
rect 75808 5412 75864 5468
rect 75864 5412 75868 5468
rect 75804 5408 75868 5412
rect 75884 5468 75948 5472
rect 75884 5412 75888 5468
rect 75888 5412 75944 5468
rect 75944 5412 75948 5468
rect 75884 5408 75948 5412
rect 75964 5468 76028 5472
rect 75964 5412 75968 5468
rect 75968 5412 76024 5468
rect 76024 5412 76028 5468
rect 75964 5408 76028 5412
rect 19384 4924 19448 4928
rect 19384 4868 19388 4924
rect 19388 4868 19444 4924
rect 19444 4868 19448 4924
rect 19384 4864 19448 4868
rect 19464 4924 19528 4928
rect 19464 4868 19468 4924
rect 19468 4868 19524 4924
rect 19524 4868 19528 4924
rect 19464 4864 19528 4868
rect 19544 4924 19608 4928
rect 19544 4868 19548 4924
rect 19548 4868 19604 4924
rect 19604 4868 19608 4924
rect 19544 4864 19608 4868
rect 19624 4924 19688 4928
rect 19624 4868 19628 4924
rect 19628 4868 19684 4924
rect 19684 4868 19688 4924
rect 19624 4864 19688 4868
rect 38384 4924 38448 4928
rect 38384 4868 38388 4924
rect 38388 4868 38444 4924
rect 38444 4868 38448 4924
rect 38384 4864 38448 4868
rect 38464 4924 38528 4928
rect 38464 4868 38468 4924
rect 38468 4868 38524 4924
rect 38524 4868 38528 4924
rect 38464 4864 38528 4868
rect 38544 4924 38608 4928
rect 38544 4868 38548 4924
rect 38548 4868 38604 4924
rect 38604 4868 38608 4924
rect 38544 4864 38608 4868
rect 38624 4924 38688 4928
rect 38624 4868 38628 4924
rect 38628 4868 38684 4924
rect 38684 4868 38688 4924
rect 38624 4864 38688 4868
rect 57384 4924 57448 4928
rect 57384 4868 57388 4924
rect 57388 4868 57444 4924
rect 57444 4868 57448 4924
rect 57384 4864 57448 4868
rect 57464 4924 57528 4928
rect 57464 4868 57468 4924
rect 57468 4868 57524 4924
rect 57524 4868 57528 4924
rect 57464 4864 57528 4868
rect 57544 4924 57608 4928
rect 57544 4868 57548 4924
rect 57548 4868 57604 4924
rect 57604 4868 57608 4924
rect 57544 4864 57608 4868
rect 57624 4924 57688 4928
rect 57624 4868 57628 4924
rect 57628 4868 57684 4924
rect 57684 4868 57688 4924
rect 57624 4864 57688 4868
rect 76384 4924 76448 4928
rect 76384 4868 76388 4924
rect 76388 4868 76444 4924
rect 76444 4868 76448 4924
rect 76384 4864 76448 4868
rect 76464 4924 76528 4928
rect 76464 4868 76468 4924
rect 76468 4868 76524 4924
rect 76524 4868 76528 4924
rect 76464 4864 76528 4868
rect 76544 4924 76608 4928
rect 76544 4868 76548 4924
rect 76548 4868 76604 4924
rect 76604 4868 76608 4924
rect 76544 4864 76608 4868
rect 76624 4924 76688 4928
rect 76624 4868 76628 4924
rect 76628 4868 76684 4924
rect 76684 4868 76688 4924
rect 76624 4864 76688 4868
<< metal4 >>
rect 2696 91354 3016 91396
rect 2696 91118 2738 91354
rect 2974 91118 3016 91354
rect 2696 76674 3016 91118
rect 2696 76438 2738 76674
rect 2974 76438 3016 76674
rect 2696 57674 3016 76438
rect 2696 57438 2738 57674
rect 2974 57438 3016 57674
rect 2696 38674 3016 57438
rect 2696 38438 2738 38674
rect 2974 38438 3016 38674
rect 2696 19674 3016 38438
rect 2696 19438 2738 19674
rect 2974 19438 3016 19674
rect 2696 2994 3016 19438
rect 3356 90694 3676 90736
rect 3356 90458 3398 90694
rect 3634 90458 3676 90694
rect 3356 76014 3676 90458
rect 18716 90694 19036 91396
rect 18716 90458 18758 90694
rect 18994 90458 19036 90694
rect 18716 89248 19036 90458
rect 18716 89184 18724 89248
rect 18788 89184 18804 89248
rect 18868 89184 18884 89248
rect 18948 89184 18964 89248
rect 19028 89184 19036 89248
rect 18716 88160 19036 89184
rect 18716 88096 18724 88160
rect 18788 88096 18804 88160
rect 18868 88096 18884 88160
rect 18948 88096 18964 88160
rect 19028 88096 19036 88160
rect 3356 75778 3398 76014
rect 3634 75778 3676 76014
rect 3356 57014 3676 75778
rect 3356 56778 3398 57014
rect 3634 56778 3676 57014
rect 3356 38014 3676 56778
rect 3356 37778 3398 38014
rect 3634 37778 3676 38014
rect 3356 19014 3676 37778
rect 3356 18778 3398 19014
rect 3634 18778 3676 19014
rect 3356 3654 3676 18778
rect 5948 87072 6268 87088
rect 5948 87008 5956 87072
rect 6020 87008 6036 87072
rect 6100 87008 6116 87072
rect 6180 87008 6196 87072
rect 6260 87008 6268 87072
rect 5948 85984 6268 87008
rect 5948 85920 5956 85984
rect 6020 85920 6036 85984
rect 6100 85920 6116 85984
rect 6180 85920 6196 85984
rect 6260 85920 6268 85984
rect 5948 84896 6268 85920
rect 5948 84832 5956 84896
rect 6020 84832 6036 84896
rect 6100 84832 6116 84896
rect 6180 84832 6196 84896
rect 6260 84832 6268 84896
rect 5948 83808 6268 84832
rect 5948 83744 5956 83808
rect 6020 83744 6036 83808
rect 6100 83744 6116 83808
rect 6180 83744 6196 83808
rect 6260 83744 6268 83808
rect 5948 82720 6268 83744
rect 5948 82656 5956 82720
rect 6020 82656 6036 82720
rect 6100 82656 6116 82720
rect 6180 82656 6196 82720
rect 6260 82656 6268 82720
rect 5948 81632 6268 82656
rect 5948 81568 5956 81632
rect 6020 81568 6036 81632
rect 6100 81568 6116 81632
rect 6180 81568 6196 81632
rect 6260 81568 6268 81632
rect 5948 80544 6268 81568
rect 5948 80480 5956 80544
rect 6020 80480 6036 80544
rect 6100 80480 6116 80544
rect 6180 80480 6196 80544
rect 6260 80480 6268 80544
rect 5948 79456 6268 80480
rect 5948 79392 5956 79456
rect 6020 79392 6036 79456
rect 6100 79392 6116 79456
rect 6180 79392 6196 79456
rect 6260 79392 6268 79456
rect 5948 78368 6268 79392
rect 5948 78304 5956 78368
rect 6020 78304 6036 78368
rect 6100 78304 6116 78368
rect 6180 78304 6196 78368
rect 6260 78304 6268 78368
rect 5948 77280 6268 78304
rect 5948 77216 5956 77280
rect 6020 77216 6036 77280
rect 6100 77216 6116 77280
rect 6180 77216 6196 77280
rect 6260 77216 6268 77280
rect 5948 76192 6268 77216
rect 5948 76128 5956 76192
rect 6020 76128 6036 76192
rect 6100 76128 6116 76192
rect 6180 76128 6196 76192
rect 6260 76128 6268 76192
rect 5948 76014 6268 76128
rect 5948 75778 5990 76014
rect 6226 75778 6268 76014
rect 5948 75104 6268 75778
rect 5948 75040 5956 75104
rect 6020 75040 6036 75104
rect 6100 75040 6116 75104
rect 6180 75040 6196 75104
rect 6260 75040 6268 75104
rect 5948 74016 6268 75040
rect 5948 73952 5956 74016
rect 6020 73952 6036 74016
rect 6100 73952 6116 74016
rect 6180 73952 6196 74016
rect 6260 73952 6268 74016
rect 5948 72928 6268 73952
rect 5948 72864 5956 72928
rect 6020 72864 6036 72928
rect 6100 72864 6116 72928
rect 6180 72864 6196 72928
rect 6260 72864 6268 72928
rect 5948 71840 6268 72864
rect 5948 71776 5956 71840
rect 6020 71776 6036 71840
rect 6100 71776 6116 71840
rect 6180 71776 6196 71840
rect 6260 71776 6268 71840
rect 5948 70752 6268 71776
rect 5948 70688 5956 70752
rect 6020 70688 6036 70752
rect 6100 70688 6116 70752
rect 6180 70688 6196 70752
rect 6260 70688 6268 70752
rect 5948 69664 6268 70688
rect 5948 69600 5956 69664
rect 6020 69600 6036 69664
rect 6100 69600 6116 69664
rect 6180 69600 6196 69664
rect 6260 69600 6268 69664
rect 5948 68576 6268 69600
rect 5948 68512 5956 68576
rect 6020 68512 6036 68576
rect 6100 68512 6116 68576
rect 6180 68512 6196 68576
rect 6260 68512 6268 68576
rect 5948 67488 6268 68512
rect 5948 67424 5956 67488
rect 6020 67424 6036 67488
rect 6100 67424 6116 67488
rect 6180 67424 6196 67488
rect 6260 67424 6268 67488
rect 5948 66400 6268 67424
rect 5948 66336 5956 66400
rect 6020 66336 6036 66400
rect 6100 66336 6116 66400
rect 6180 66336 6196 66400
rect 6260 66336 6268 66400
rect 5948 65312 6268 66336
rect 5948 65248 5956 65312
rect 6020 65248 6036 65312
rect 6100 65248 6116 65312
rect 6180 65248 6196 65312
rect 6260 65248 6268 65312
rect 5948 64224 6268 65248
rect 5948 64160 5956 64224
rect 6020 64160 6036 64224
rect 6100 64160 6116 64224
rect 6180 64160 6196 64224
rect 6260 64160 6268 64224
rect 5948 63136 6268 64160
rect 5948 63072 5956 63136
rect 6020 63072 6036 63136
rect 6100 63072 6116 63136
rect 6180 63072 6196 63136
rect 6260 63072 6268 63136
rect 5948 62048 6268 63072
rect 5948 61984 5956 62048
rect 6020 61984 6036 62048
rect 6100 61984 6116 62048
rect 6180 61984 6196 62048
rect 6260 61984 6268 62048
rect 5948 60960 6268 61984
rect 5948 60896 5956 60960
rect 6020 60896 6036 60960
rect 6100 60896 6116 60960
rect 6180 60896 6196 60960
rect 6260 60896 6268 60960
rect 5948 59872 6268 60896
rect 5948 59808 5956 59872
rect 6020 59808 6036 59872
rect 6100 59808 6116 59872
rect 6180 59808 6196 59872
rect 6260 59808 6268 59872
rect 5948 58784 6268 59808
rect 5948 58720 5956 58784
rect 6020 58720 6036 58784
rect 6100 58720 6116 58784
rect 6180 58720 6196 58784
rect 6260 58720 6268 58784
rect 5948 57696 6268 58720
rect 5948 57632 5956 57696
rect 6020 57632 6036 57696
rect 6100 57632 6116 57696
rect 6180 57632 6196 57696
rect 6260 57632 6268 57696
rect 5948 57014 6268 57632
rect 5948 56778 5990 57014
rect 6226 56778 6268 57014
rect 5948 56608 6268 56778
rect 5948 56544 5956 56608
rect 6020 56544 6036 56608
rect 6100 56544 6116 56608
rect 6180 56544 6196 56608
rect 6260 56544 6268 56608
rect 5948 55520 6268 56544
rect 5948 55456 5956 55520
rect 6020 55456 6036 55520
rect 6100 55456 6116 55520
rect 6180 55456 6196 55520
rect 6260 55456 6268 55520
rect 5948 54432 6268 55456
rect 5948 54368 5956 54432
rect 6020 54368 6036 54432
rect 6100 54368 6116 54432
rect 6180 54368 6196 54432
rect 6260 54368 6268 54432
rect 5948 53344 6268 54368
rect 5948 53280 5956 53344
rect 6020 53280 6036 53344
rect 6100 53280 6116 53344
rect 6180 53280 6196 53344
rect 6260 53280 6268 53344
rect 5948 52256 6268 53280
rect 5948 52192 5956 52256
rect 6020 52192 6036 52256
rect 6100 52192 6116 52256
rect 6180 52192 6196 52256
rect 6260 52192 6268 52256
rect 5948 51168 6268 52192
rect 5948 51104 5956 51168
rect 6020 51104 6036 51168
rect 6100 51104 6116 51168
rect 6180 51104 6196 51168
rect 6260 51104 6268 51168
rect 5948 50080 6268 51104
rect 5948 50016 5956 50080
rect 6020 50016 6036 50080
rect 6100 50016 6116 50080
rect 6180 50016 6196 50080
rect 6260 50016 6268 50080
rect 5948 48992 6268 50016
rect 5948 48928 5956 48992
rect 6020 48928 6036 48992
rect 6100 48928 6116 48992
rect 6180 48928 6196 48992
rect 6260 48928 6268 48992
rect 5948 47904 6268 48928
rect 5948 47840 5956 47904
rect 6020 47840 6036 47904
rect 6100 47840 6116 47904
rect 6180 47840 6196 47904
rect 6260 47840 6268 47904
rect 5948 46816 6268 47840
rect 5948 46752 5956 46816
rect 6020 46752 6036 46816
rect 6100 46752 6116 46816
rect 6180 46752 6196 46816
rect 6260 46752 6268 46816
rect 5948 45728 6268 46752
rect 5948 45664 5956 45728
rect 6020 45664 6036 45728
rect 6100 45664 6116 45728
rect 6180 45664 6196 45728
rect 6260 45664 6268 45728
rect 5948 44640 6268 45664
rect 5948 44576 5956 44640
rect 6020 44576 6036 44640
rect 6100 44576 6116 44640
rect 6180 44576 6196 44640
rect 6260 44576 6268 44640
rect 5948 43552 6268 44576
rect 5948 43488 5956 43552
rect 6020 43488 6036 43552
rect 6100 43488 6116 43552
rect 6180 43488 6196 43552
rect 6260 43488 6268 43552
rect 5948 42464 6268 43488
rect 5948 42400 5956 42464
rect 6020 42400 6036 42464
rect 6100 42400 6116 42464
rect 6180 42400 6196 42464
rect 6260 42400 6268 42464
rect 5948 41376 6268 42400
rect 5948 41312 5956 41376
rect 6020 41312 6036 41376
rect 6100 41312 6116 41376
rect 6180 41312 6196 41376
rect 6260 41312 6268 41376
rect 5948 40288 6268 41312
rect 5948 40224 5956 40288
rect 6020 40224 6036 40288
rect 6100 40224 6116 40288
rect 6180 40224 6196 40288
rect 6260 40224 6268 40288
rect 5948 39200 6268 40224
rect 5948 39136 5956 39200
rect 6020 39136 6036 39200
rect 6100 39136 6116 39200
rect 6180 39136 6196 39200
rect 6260 39136 6268 39200
rect 5948 38112 6268 39136
rect 5948 38048 5956 38112
rect 6020 38048 6036 38112
rect 6100 38048 6116 38112
rect 6180 38048 6196 38112
rect 6260 38048 6268 38112
rect 5948 38014 6268 38048
rect 5948 37778 5990 38014
rect 6226 37778 6268 38014
rect 5948 37024 6268 37778
rect 5948 36960 5956 37024
rect 6020 36960 6036 37024
rect 6100 36960 6116 37024
rect 6180 36960 6196 37024
rect 6260 36960 6268 37024
rect 5948 35936 6268 36960
rect 5948 35872 5956 35936
rect 6020 35872 6036 35936
rect 6100 35872 6116 35936
rect 6180 35872 6196 35936
rect 6260 35872 6268 35936
rect 5948 34848 6268 35872
rect 5948 34784 5956 34848
rect 6020 34784 6036 34848
rect 6100 34784 6116 34848
rect 6180 34784 6196 34848
rect 6260 34784 6268 34848
rect 5948 33760 6268 34784
rect 5948 33696 5956 33760
rect 6020 33696 6036 33760
rect 6100 33696 6116 33760
rect 6180 33696 6196 33760
rect 6260 33696 6268 33760
rect 5948 32672 6268 33696
rect 5948 32608 5956 32672
rect 6020 32608 6036 32672
rect 6100 32608 6116 32672
rect 6180 32608 6196 32672
rect 6260 32608 6268 32672
rect 5948 31584 6268 32608
rect 5948 31520 5956 31584
rect 6020 31520 6036 31584
rect 6100 31520 6116 31584
rect 6180 31520 6196 31584
rect 6260 31520 6268 31584
rect 5948 30496 6268 31520
rect 5948 30432 5956 30496
rect 6020 30432 6036 30496
rect 6100 30432 6116 30496
rect 6180 30432 6196 30496
rect 6260 30432 6268 30496
rect 5948 29408 6268 30432
rect 5948 29344 5956 29408
rect 6020 29344 6036 29408
rect 6100 29344 6116 29408
rect 6180 29344 6196 29408
rect 6260 29344 6268 29408
rect 5948 28320 6268 29344
rect 5948 28256 5956 28320
rect 6020 28256 6036 28320
rect 6100 28256 6116 28320
rect 6180 28256 6196 28320
rect 6260 28256 6268 28320
rect 5948 27232 6268 28256
rect 5948 27168 5956 27232
rect 6020 27168 6036 27232
rect 6100 27168 6116 27232
rect 6180 27168 6196 27232
rect 6260 27168 6268 27232
rect 5948 26144 6268 27168
rect 5948 26080 5956 26144
rect 6020 26080 6036 26144
rect 6100 26080 6116 26144
rect 6180 26080 6196 26144
rect 6260 26080 6268 26144
rect 5948 25056 6268 26080
rect 5948 24992 5956 25056
rect 6020 24992 6036 25056
rect 6100 24992 6116 25056
rect 6180 24992 6196 25056
rect 6260 24992 6268 25056
rect 5948 23968 6268 24992
rect 5948 23904 5956 23968
rect 6020 23904 6036 23968
rect 6100 23904 6116 23968
rect 6180 23904 6196 23968
rect 6260 23904 6268 23968
rect 5948 22880 6268 23904
rect 5948 22816 5956 22880
rect 6020 22816 6036 22880
rect 6100 22816 6116 22880
rect 6180 22816 6196 22880
rect 6260 22816 6268 22880
rect 5948 21792 6268 22816
rect 5948 21728 5956 21792
rect 6020 21728 6036 21792
rect 6100 21728 6116 21792
rect 6180 21728 6196 21792
rect 6260 21728 6268 21792
rect 5948 20704 6268 21728
rect 5948 20640 5956 20704
rect 6020 20640 6036 20704
rect 6100 20640 6116 20704
rect 6180 20640 6196 20704
rect 6260 20640 6268 20704
rect 5948 19616 6268 20640
rect 5948 19552 5956 19616
rect 6020 19552 6036 19616
rect 6100 19552 6116 19616
rect 6180 19552 6196 19616
rect 6260 19552 6268 19616
rect 5948 19014 6268 19552
rect 5948 18778 5990 19014
rect 6226 18778 6268 19014
rect 5948 18528 6268 18778
rect 5948 18464 5956 18528
rect 6020 18464 6036 18528
rect 6100 18464 6116 18528
rect 6180 18464 6196 18528
rect 6260 18464 6268 18528
rect 5948 17440 6268 18464
rect 5948 17376 5956 17440
rect 6020 17376 6036 17440
rect 6100 17376 6116 17440
rect 6180 17376 6196 17440
rect 6260 17376 6268 17440
rect 5948 16352 6268 17376
rect 5948 16288 5956 16352
rect 6020 16288 6036 16352
rect 6100 16288 6116 16352
rect 6180 16288 6196 16352
rect 6260 16288 6268 16352
rect 5948 15264 6268 16288
rect 5948 15200 5956 15264
rect 6020 15200 6036 15264
rect 6100 15200 6116 15264
rect 6180 15200 6196 15264
rect 6260 15200 6268 15264
rect 5948 14176 6268 15200
rect 5948 14112 5956 14176
rect 6020 14112 6036 14176
rect 6100 14112 6116 14176
rect 6180 14112 6196 14176
rect 6260 14112 6268 14176
rect 5948 13088 6268 14112
rect 5948 13024 5956 13088
rect 6020 13024 6036 13088
rect 6100 13024 6116 13088
rect 6180 13024 6196 13088
rect 6260 13024 6268 13088
rect 5948 12000 6268 13024
rect 5948 11936 5956 12000
rect 6020 11936 6036 12000
rect 6100 11936 6116 12000
rect 6180 11936 6196 12000
rect 6260 11936 6268 12000
rect 5948 10912 6268 11936
rect 5948 10848 5956 10912
rect 6020 10848 6036 10912
rect 6100 10848 6116 10912
rect 6180 10848 6196 10912
rect 6260 10848 6268 10912
rect 5948 9824 6268 10848
rect 5948 9760 5956 9824
rect 6020 9760 6036 9824
rect 6100 9760 6116 9824
rect 6180 9760 6196 9824
rect 6260 9760 6268 9824
rect 5948 8736 6268 9760
rect 5948 8672 5956 8736
rect 6020 8672 6036 8736
rect 6100 8672 6116 8736
rect 6180 8672 6196 8736
rect 6260 8672 6268 8736
rect 5948 7648 6268 8672
rect 5948 7584 5956 7648
rect 6020 7584 6036 7648
rect 6100 7584 6116 7648
rect 6180 7584 6196 7648
rect 6260 7584 6268 7648
rect 5948 7024 6268 7584
rect 6684 86528 7004 87088
rect 6684 86464 6692 86528
rect 6756 86464 6772 86528
rect 6836 86464 6852 86528
rect 6916 86464 6932 86528
rect 6996 86464 7004 86528
rect 6684 85440 7004 86464
rect 18716 87072 19036 88096
rect 18716 87008 18724 87072
rect 18788 87008 18804 87072
rect 18868 87008 18884 87072
rect 18948 87008 18964 87072
rect 19028 87008 19036 87072
rect 18716 85601 19036 87008
rect 19376 91354 19696 91396
rect 19376 91118 19418 91354
rect 19654 91118 19696 91354
rect 19376 88704 19696 91118
rect 19376 88640 19384 88704
rect 19448 88640 19464 88704
rect 19528 88640 19544 88704
rect 19608 88640 19624 88704
rect 19688 88640 19696 88704
rect 19376 87616 19696 88640
rect 19376 87552 19384 87616
rect 19448 87552 19464 87616
rect 19528 87552 19544 87616
rect 19608 87552 19624 87616
rect 19688 87552 19696 87616
rect 19376 86528 19696 87552
rect 19376 86464 19384 86528
rect 19448 86464 19464 86528
rect 19528 86464 19544 86528
rect 19608 86464 19624 86528
rect 19688 86464 19696 86528
rect 19376 85601 19696 86464
rect 37716 90694 38036 91396
rect 37716 90458 37758 90694
rect 37994 90458 38036 90694
rect 37716 89248 38036 90458
rect 37716 89184 37724 89248
rect 37788 89184 37804 89248
rect 37868 89184 37884 89248
rect 37948 89184 37964 89248
rect 38028 89184 38036 89248
rect 37716 88160 38036 89184
rect 37716 88096 37724 88160
rect 37788 88096 37804 88160
rect 37868 88096 37884 88160
rect 37948 88096 37964 88160
rect 38028 88096 38036 88160
rect 37716 87072 38036 88096
rect 37716 87008 37724 87072
rect 37788 87008 37804 87072
rect 37868 87008 37884 87072
rect 37948 87008 37964 87072
rect 38028 87008 38036 87072
rect 37716 85601 38036 87008
rect 38376 91354 38696 91396
rect 38376 91118 38418 91354
rect 38654 91118 38696 91354
rect 38376 88704 38696 91118
rect 38376 88640 38384 88704
rect 38448 88640 38464 88704
rect 38528 88640 38544 88704
rect 38608 88640 38624 88704
rect 38688 88640 38696 88704
rect 38376 87616 38696 88640
rect 38376 87552 38384 87616
rect 38448 87552 38464 87616
rect 38528 87552 38544 87616
rect 38608 87552 38624 87616
rect 38688 87552 38696 87616
rect 38376 86528 38696 87552
rect 38376 86464 38384 86528
rect 38448 86464 38464 86528
rect 38528 86464 38544 86528
rect 38608 86464 38624 86528
rect 38688 86464 38696 86528
rect 38376 85601 38696 86464
rect 56716 90694 57036 91396
rect 56716 90458 56758 90694
rect 56994 90458 57036 90694
rect 56716 89248 57036 90458
rect 56716 89184 56724 89248
rect 56788 89184 56804 89248
rect 56868 89184 56884 89248
rect 56948 89184 56964 89248
rect 57028 89184 57036 89248
rect 56716 88160 57036 89184
rect 56716 88096 56724 88160
rect 56788 88096 56804 88160
rect 56868 88096 56884 88160
rect 56948 88096 56964 88160
rect 57028 88096 57036 88160
rect 56716 87072 57036 88096
rect 56716 87008 56724 87072
rect 56788 87008 56804 87072
rect 56868 87008 56884 87072
rect 56948 87008 56964 87072
rect 57028 87008 57036 87072
rect 56716 85601 57036 87008
rect 57376 91354 57696 91396
rect 57376 91118 57418 91354
rect 57654 91118 57696 91354
rect 57376 88704 57696 91118
rect 57376 88640 57384 88704
rect 57448 88640 57464 88704
rect 57528 88640 57544 88704
rect 57608 88640 57624 88704
rect 57688 88640 57696 88704
rect 57376 87616 57696 88640
rect 57376 87552 57384 87616
rect 57448 87552 57464 87616
rect 57528 87552 57544 87616
rect 57608 87552 57624 87616
rect 57688 87552 57696 87616
rect 57376 86528 57696 87552
rect 57376 86464 57384 86528
rect 57448 86464 57464 86528
rect 57528 86464 57544 86528
rect 57608 86464 57624 86528
rect 57688 86464 57696 86528
rect 57376 85601 57696 86464
rect 75716 90694 76036 91396
rect 75716 90458 75758 90694
rect 75994 90458 76036 90694
rect 75716 89248 76036 90458
rect 75716 89184 75724 89248
rect 75788 89184 75804 89248
rect 75868 89184 75884 89248
rect 75948 89184 75964 89248
rect 76028 89184 76036 89248
rect 75716 88160 76036 89184
rect 75716 88096 75724 88160
rect 75788 88096 75804 88160
rect 75868 88096 75884 88160
rect 75948 88096 75964 88160
rect 76028 88096 76036 88160
rect 75716 87072 76036 88096
rect 75716 87008 75724 87072
rect 75788 87008 75804 87072
rect 75868 87008 75884 87072
rect 75948 87008 75964 87072
rect 76028 87008 76036 87072
rect 75716 85601 76036 87008
rect 76376 91354 76696 91396
rect 76376 91118 76418 91354
rect 76654 91118 76696 91354
rect 76376 88704 76696 91118
rect 90824 91354 91144 91396
rect 90824 91118 90866 91354
rect 91102 91118 91144 91354
rect 76376 88640 76384 88704
rect 76448 88640 76464 88704
rect 76528 88640 76544 88704
rect 76608 88640 76624 88704
rect 76688 88640 76696 88704
rect 76376 87616 76696 88640
rect 76376 87552 76384 87616
rect 76448 87552 76464 87616
rect 76528 87552 76544 87616
rect 76608 87552 76624 87616
rect 76688 87552 76696 87616
rect 76376 86528 76696 87552
rect 90164 90694 90484 90736
rect 90164 90458 90206 90694
rect 90442 90458 90484 90694
rect 76376 86464 76384 86528
rect 76448 86464 76464 86528
rect 76528 86464 76544 86528
rect 76608 86464 76624 86528
rect 76688 86464 76696 86528
rect 76376 85601 76696 86464
rect 87092 87072 87412 87088
rect 87092 87008 87100 87072
rect 87164 87008 87180 87072
rect 87244 87008 87260 87072
rect 87324 87008 87340 87072
rect 87404 87008 87412 87072
rect 87092 85984 87412 87008
rect 87092 85920 87100 85984
rect 87164 85920 87180 85984
rect 87244 85920 87260 85984
rect 87324 85920 87340 85984
rect 87404 85920 87412 85984
rect 6684 85376 6692 85440
rect 6756 85376 6772 85440
rect 6836 85376 6852 85440
rect 6916 85376 6932 85440
rect 6996 85376 7004 85440
rect 6684 84352 7004 85376
rect 6684 84288 6692 84352
rect 6756 84288 6772 84352
rect 6836 84288 6852 84352
rect 6916 84288 6932 84352
rect 6996 84288 7004 84352
rect 6684 83264 7004 84288
rect 87092 84896 87412 85920
rect 87092 84832 87100 84896
rect 87164 84832 87180 84896
rect 87244 84832 87260 84896
rect 87324 84832 87340 84896
rect 87404 84832 87412 84896
rect 87092 83808 87412 84832
rect 87092 83744 87100 83808
rect 87164 83744 87180 83808
rect 87244 83744 87260 83808
rect 87324 83744 87340 83808
rect 87404 83744 87412 83808
rect 6684 83200 6692 83264
rect 6756 83200 6772 83264
rect 6836 83200 6852 83264
rect 6916 83200 6932 83264
rect 6996 83200 7004 83264
rect 6684 82176 7004 83200
rect 11144 83030 11186 83266
rect 11422 83030 11464 83266
rect 45144 83030 45186 83266
rect 45422 83030 45464 83266
rect 48144 83030 48186 83266
rect 48422 83030 48464 83266
rect 82144 83030 82186 83266
rect 82422 83030 82464 83266
rect 87092 82720 87412 83744
rect 87092 82656 87100 82720
rect 87164 82656 87180 82720
rect 87244 82656 87260 82720
rect 87324 82656 87340 82720
rect 87404 82656 87412 82720
rect 10484 82370 10526 82606
rect 10762 82370 10804 82606
rect 44484 82370 44526 82606
rect 44762 82370 44804 82606
rect 47484 82370 47526 82606
rect 47762 82370 47804 82606
rect 81484 82370 81526 82606
rect 81762 82370 81804 82606
rect 6684 82112 6692 82176
rect 6756 82112 6772 82176
rect 6836 82112 6852 82176
rect 6916 82112 6932 82176
rect 6996 82112 7004 82176
rect 6684 81088 7004 82112
rect 6684 81024 6692 81088
rect 6756 81024 6772 81088
rect 6836 81024 6852 81088
rect 6916 81024 6932 81088
rect 6996 81024 7004 81088
rect 6684 80000 7004 81024
rect 6684 79936 6692 80000
rect 6756 79936 6772 80000
rect 6836 79936 6852 80000
rect 6916 79936 6932 80000
rect 6996 79936 7004 80000
rect 6684 78912 7004 79936
rect 6684 78848 6692 78912
rect 6756 78848 6772 78912
rect 6836 78848 6852 78912
rect 6916 78848 6932 78912
rect 6996 78848 7004 78912
rect 6684 77824 7004 78848
rect 6684 77760 6692 77824
rect 6756 77760 6772 77824
rect 6836 77760 6852 77824
rect 6916 77760 6932 77824
rect 6996 77760 7004 77824
rect 6684 76736 7004 77760
rect 6684 76672 6692 76736
rect 6756 76674 6772 76736
rect 6836 76674 6852 76736
rect 6916 76674 6932 76736
rect 6996 76672 7004 76736
rect 87092 81632 87412 82656
rect 87092 81568 87100 81632
rect 87164 81568 87180 81632
rect 87244 81568 87260 81632
rect 87324 81568 87340 81632
rect 87404 81568 87412 81632
rect 87092 80544 87412 81568
rect 87092 80480 87100 80544
rect 87164 80480 87180 80544
rect 87244 80480 87260 80544
rect 87324 80480 87340 80544
rect 87404 80480 87412 80544
rect 87092 79456 87412 80480
rect 87092 79392 87100 79456
rect 87164 79392 87180 79456
rect 87244 79392 87260 79456
rect 87324 79392 87340 79456
rect 87404 79392 87412 79456
rect 87092 78368 87412 79392
rect 87092 78304 87100 78368
rect 87164 78304 87180 78368
rect 87244 78304 87260 78368
rect 87324 78304 87340 78368
rect 87404 78304 87412 78368
rect 87092 77280 87412 78304
rect 87092 77216 87100 77280
rect 87164 77216 87180 77280
rect 87244 77216 87260 77280
rect 87324 77216 87340 77280
rect 87404 77216 87412 77280
rect 6684 76438 6726 76672
rect 6962 76438 7004 76672
rect 11144 76438 11186 76674
rect 11422 76438 11464 76674
rect 45144 76438 45186 76674
rect 45422 76438 45464 76674
rect 48144 76438 48186 76674
rect 48422 76438 48464 76674
rect 82144 76438 82186 76674
rect 82422 76438 82464 76674
rect 6684 75648 7004 76438
rect 87092 76192 87412 77216
rect 87092 76128 87100 76192
rect 87164 76128 87180 76192
rect 87244 76128 87260 76192
rect 87324 76128 87340 76192
rect 87404 76128 87412 76192
rect 87092 76014 87412 76128
rect 10484 75778 10526 76014
rect 10762 75778 10804 76014
rect 44484 75778 44526 76014
rect 44762 75778 44804 76014
rect 47484 75778 47526 76014
rect 47762 75778 47804 76014
rect 81484 75778 81526 76014
rect 81762 75778 81804 76014
rect 87092 75778 87134 76014
rect 87370 75778 87412 76014
rect 6684 75584 6692 75648
rect 6756 75584 6772 75648
rect 6836 75584 6852 75648
rect 6916 75584 6932 75648
rect 6996 75584 7004 75648
rect 6684 74560 7004 75584
rect 6684 74496 6692 74560
rect 6756 74496 6772 74560
rect 6836 74496 6852 74560
rect 6916 74496 6932 74560
rect 6996 74496 7004 74560
rect 6684 73472 7004 74496
rect 6684 73408 6692 73472
rect 6756 73408 6772 73472
rect 6836 73408 6852 73472
rect 6916 73408 6932 73472
rect 6996 73408 7004 73472
rect 6684 72384 7004 73408
rect 6684 72320 6692 72384
rect 6756 72320 6772 72384
rect 6836 72320 6852 72384
rect 6916 72320 6932 72384
rect 6996 72320 7004 72384
rect 6684 71296 7004 72320
rect 6684 71232 6692 71296
rect 6756 71232 6772 71296
rect 6836 71232 6852 71296
rect 6916 71232 6932 71296
rect 6996 71232 7004 71296
rect 6684 70208 7004 71232
rect 6684 70144 6692 70208
rect 6756 70144 6772 70208
rect 6836 70144 6852 70208
rect 6916 70144 6932 70208
rect 6996 70144 7004 70208
rect 6684 69120 7004 70144
rect 6684 69056 6692 69120
rect 6756 69056 6772 69120
rect 6836 69056 6852 69120
rect 6916 69056 6932 69120
rect 6996 69056 7004 69120
rect 6684 68032 7004 69056
rect 6684 67968 6692 68032
rect 6756 67968 6772 68032
rect 6836 67968 6852 68032
rect 6916 67968 6932 68032
rect 6996 67968 7004 68032
rect 6684 66944 7004 67968
rect 6684 66880 6692 66944
rect 6756 66880 6772 66944
rect 6836 66880 6852 66944
rect 6916 66880 6932 66944
rect 6996 66880 7004 66944
rect 6684 65856 7004 66880
rect 6684 65792 6692 65856
rect 6756 65792 6772 65856
rect 6836 65792 6852 65856
rect 6916 65792 6932 65856
rect 6996 65792 7004 65856
rect 6684 64768 7004 65792
rect 6684 64704 6692 64768
rect 6756 64704 6772 64768
rect 6836 64704 6852 64768
rect 6916 64704 6932 64768
rect 6996 64704 7004 64768
rect 6684 63680 7004 64704
rect 6684 63616 6692 63680
rect 6756 63616 6772 63680
rect 6836 63616 6852 63680
rect 6916 63616 6932 63680
rect 6996 63616 7004 63680
rect 6684 62592 7004 63616
rect 6684 62528 6692 62592
rect 6756 62528 6772 62592
rect 6836 62528 6852 62592
rect 6916 62528 6932 62592
rect 6996 62528 7004 62592
rect 6684 61504 7004 62528
rect 6684 61440 6692 61504
rect 6756 61440 6772 61504
rect 6836 61440 6852 61504
rect 6916 61440 6932 61504
rect 6996 61440 7004 61504
rect 6684 60416 7004 61440
rect 6684 60352 6692 60416
rect 6756 60352 6772 60416
rect 6836 60352 6852 60416
rect 6916 60352 6932 60416
rect 6996 60352 7004 60416
rect 6684 59328 7004 60352
rect 6684 59264 6692 59328
rect 6756 59264 6772 59328
rect 6836 59264 6852 59328
rect 6916 59264 6932 59328
rect 6996 59264 7004 59328
rect 6684 58240 7004 59264
rect 6684 58176 6692 58240
rect 6756 58176 6772 58240
rect 6836 58176 6852 58240
rect 6916 58176 6932 58240
rect 6996 58176 7004 58240
rect 6684 57674 7004 58176
rect 87092 75104 87412 75778
rect 87092 75040 87100 75104
rect 87164 75040 87180 75104
rect 87244 75040 87260 75104
rect 87324 75040 87340 75104
rect 87404 75040 87412 75104
rect 87092 74016 87412 75040
rect 87092 73952 87100 74016
rect 87164 73952 87180 74016
rect 87244 73952 87260 74016
rect 87324 73952 87340 74016
rect 87404 73952 87412 74016
rect 87092 72928 87412 73952
rect 87092 72864 87100 72928
rect 87164 72864 87180 72928
rect 87244 72864 87260 72928
rect 87324 72864 87340 72928
rect 87404 72864 87412 72928
rect 87092 71840 87412 72864
rect 87092 71776 87100 71840
rect 87164 71776 87180 71840
rect 87244 71776 87260 71840
rect 87324 71776 87340 71840
rect 87404 71776 87412 71840
rect 87092 70752 87412 71776
rect 87092 70688 87100 70752
rect 87164 70688 87180 70752
rect 87244 70688 87260 70752
rect 87324 70688 87340 70752
rect 87404 70688 87412 70752
rect 87092 69664 87412 70688
rect 87092 69600 87100 69664
rect 87164 69600 87180 69664
rect 87244 69600 87260 69664
rect 87324 69600 87340 69664
rect 87404 69600 87412 69664
rect 87092 68576 87412 69600
rect 87092 68512 87100 68576
rect 87164 68512 87180 68576
rect 87244 68512 87260 68576
rect 87324 68512 87340 68576
rect 87404 68512 87412 68576
rect 87092 67488 87412 68512
rect 87092 67424 87100 67488
rect 87164 67424 87180 67488
rect 87244 67424 87260 67488
rect 87324 67424 87340 67488
rect 87404 67424 87412 67488
rect 87092 66400 87412 67424
rect 87092 66336 87100 66400
rect 87164 66336 87180 66400
rect 87244 66336 87260 66400
rect 87324 66336 87340 66400
rect 87404 66336 87412 66400
rect 87092 65312 87412 66336
rect 87092 65248 87100 65312
rect 87164 65248 87180 65312
rect 87244 65248 87260 65312
rect 87324 65248 87340 65312
rect 87404 65248 87412 65312
rect 87092 64224 87412 65248
rect 87092 64160 87100 64224
rect 87164 64160 87180 64224
rect 87244 64160 87260 64224
rect 87324 64160 87340 64224
rect 87404 64160 87412 64224
rect 87092 63136 87412 64160
rect 87092 63072 87100 63136
rect 87164 63072 87180 63136
rect 87244 63072 87260 63136
rect 87324 63072 87340 63136
rect 87404 63072 87412 63136
rect 87092 62048 87412 63072
rect 87092 61984 87100 62048
rect 87164 61984 87180 62048
rect 87244 61984 87260 62048
rect 87324 61984 87340 62048
rect 87404 61984 87412 62048
rect 87092 60960 87412 61984
rect 87092 60896 87100 60960
rect 87164 60896 87180 60960
rect 87244 60896 87260 60960
rect 87324 60896 87340 60960
rect 87404 60896 87412 60960
rect 87092 59872 87412 60896
rect 87092 59808 87100 59872
rect 87164 59808 87180 59872
rect 87244 59808 87260 59872
rect 87324 59808 87340 59872
rect 87404 59808 87412 59872
rect 87092 58784 87412 59808
rect 87092 58720 87100 58784
rect 87164 58720 87180 58784
rect 87244 58720 87260 58784
rect 87324 58720 87340 58784
rect 87404 58720 87412 58784
rect 87092 57696 87412 58720
rect 6684 57438 6726 57674
rect 6962 57438 7004 57674
rect 11144 57438 11186 57674
rect 11422 57438 11464 57674
rect 45144 57438 45186 57674
rect 45422 57438 45464 57674
rect 48144 57438 48186 57674
rect 48422 57438 48464 57674
rect 82144 57438 82186 57674
rect 82422 57438 82464 57674
rect 87092 57632 87100 57696
rect 87164 57632 87180 57696
rect 87244 57632 87260 57696
rect 87324 57632 87340 57696
rect 87404 57632 87412 57696
rect 6684 57152 7004 57438
rect 6684 57088 6692 57152
rect 6756 57088 6772 57152
rect 6836 57088 6852 57152
rect 6916 57088 6932 57152
rect 6996 57088 7004 57152
rect 6684 56064 7004 57088
rect 87092 57014 87412 57632
rect 10484 56778 10526 57014
rect 10762 56778 10804 57014
rect 44484 56778 44526 57014
rect 44762 56778 44804 57014
rect 47484 56778 47526 57014
rect 47762 56778 47804 57014
rect 81484 56778 81526 57014
rect 81762 56778 81804 57014
rect 87092 56778 87134 57014
rect 87370 56778 87412 57014
rect 6684 56000 6692 56064
rect 6756 56000 6772 56064
rect 6836 56000 6852 56064
rect 6916 56000 6932 56064
rect 6996 56000 7004 56064
rect 6684 54976 7004 56000
rect 6684 54912 6692 54976
rect 6756 54912 6772 54976
rect 6836 54912 6852 54976
rect 6916 54912 6932 54976
rect 6996 54912 7004 54976
rect 6684 53888 7004 54912
rect 6684 53824 6692 53888
rect 6756 53824 6772 53888
rect 6836 53824 6852 53888
rect 6916 53824 6932 53888
rect 6996 53824 7004 53888
rect 6684 52800 7004 53824
rect 6684 52736 6692 52800
rect 6756 52736 6772 52800
rect 6836 52736 6852 52800
rect 6916 52736 6932 52800
rect 6996 52736 7004 52800
rect 6684 51712 7004 52736
rect 6684 51648 6692 51712
rect 6756 51648 6772 51712
rect 6836 51648 6852 51712
rect 6916 51648 6932 51712
rect 6996 51648 7004 51712
rect 6684 50624 7004 51648
rect 6684 50560 6692 50624
rect 6756 50560 6772 50624
rect 6836 50560 6852 50624
rect 6916 50560 6932 50624
rect 6996 50560 7004 50624
rect 6684 49536 7004 50560
rect 6684 49472 6692 49536
rect 6756 49472 6772 49536
rect 6836 49472 6852 49536
rect 6916 49472 6932 49536
rect 6996 49472 7004 49536
rect 6684 48448 7004 49472
rect 87092 56608 87412 56778
rect 87092 56544 87100 56608
rect 87164 56544 87180 56608
rect 87244 56544 87260 56608
rect 87324 56544 87340 56608
rect 87404 56544 87412 56608
rect 87092 55520 87412 56544
rect 87092 55456 87100 55520
rect 87164 55456 87180 55520
rect 87244 55456 87260 55520
rect 87324 55456 87340 55520
rect 87404 55456 87412 55520
rect 87092 54432 87412 55456
rect 87092 54368 87100 54432
rect 87164 54368 87180 54432
rect 87244 54368 87260 54432
rect 87324 54368 87340 54432
rect 87404 54368 87412 54432
rect 87092 53344 87412 54368
rect 87092 53280 87100 53344
rect 87164 53280 87180 53344
rect 87244 53280 87260 53344
rect 87324 53280 87340 53344
rect 87404 53280 87412 53344
rect 87092 52256 87412 53280
rect 87092 52192 87100 52256
rect 87164 52192 87180 52256
rect 87244 52192 87260 52256
rect 87324 52192 87340 52256
rect 87404 52192 87412 52256
rect 87092 51168 87412 52192
rect 87092 51104 87100 51168
rect 87164 51104 87180 51168
rect 87244 51104 87260 51168
rect 87324 51104 87340 51168
rect 87404 51104 87412 51168
rect 87092 50080 87412 51104
rect 87092 50016 87100 50080
rect 87164 50016 87180 50080
rect 87244 50016 87260 50080
rect 87324 50016 87340 50080
rect 87404 50016 87412 50080
rect 11144 49030 11186 49266
rect 11422 49030 11464 49266
rect 45144 49030 45186 49266
rect 45422 49030 45464 49266
rect 48144 49030 48186 49266
rect 48422 49030 48464 49266
rect 82144 49030 82186 49266
rect 82422 49030 82464 49266
rect 87092 48992 87412 50016
rect 87092 48928 87100 48992
rect 87164 48928 87180 48992
rect 87244 48928 87260 48992
rect 87324 48928 87340 48992
rect 87404 48928 87412 48992
rect 6684 48384 6692 48448
rect 6756 48384 6772 48448
rect 6836 48384 6852 48448
rect 6916 48384 6932 48448
rect 6996 48384 7004 48448
rect 6684 47360 7004 48384
rect 10484 48370 10526 48606
rect 10762 48370 10804 48606
rect 44484 48370 44526 48606
rect 44762 48370 44804 48606
rect 47484 48370 47526 48606
rect 47762 48370 47804 48606
rect 81484 48370 81526 48606
rect 81762 48370 81804 48606
rect 6684 47296 6692 47360
rect 6756 47296 6772 47360
rect 6836 47296 6852 47360
rect 6916 47296 6932 47360
rect 6996 47296 7004 47360
rect 6684 46272 7004 47296
rect 6684 46208 6692 46272
rect 6756 46208 6772 46272
rect 6836 46208 6852 46272
rect 6916 46208 6932 46272
rect 6996 46208 7004 46272
rect 6684 45184 7004 46208
rect 87092 47904 87412 48928
rect 87092 47840 87100 47904
rect 87164 47840 87180 47904
rect 87244 47840 87260 47904
rect 87324 47840 87340 47904
rect 87404 47840 87412 47904
rect 87092 46816 87412 47840
rect 87092 46752 87100 46816
rect 87164 46752 87180 46816
rect 87244 46752 87260 46816
rect 87324 46752 87340 46816
rect 87404 46752 87412 46816
rect 11144 45630 11186 45866
rect 11422 45630 11464 45866
rect 45144 45630 45186 45866
rect 45422 45630 45464 45866
rect 48144 45630 48186 45866
rect 48422 45630 48464 45866
rect 82144 45630 82186 45866
rect 82422 45630 82464 45866
rect 87092 45728 87412 46752
rect 87092 45664 87100 45728
rect 87164 45664 87180 45728
rect 87244 45664 87260 45728
rect 87324 45664 87340 45728
rect 87404 45664 87412 45728
rect 6684 45120 6692 45184
rect 6756 45120 6772 45184
rect 6836 45120 6852 45184
rect 6916 45120 6932 45184
rect 6996 45120 7004 45184
rect 6684 44096 7004 45120
rect 10484 44970 10526 45206
rect 10762 44970 10804 45206
rect 44484 44970 44526 45206
rect 44762 44970 44804 45206
rect 47484 44970 47526 45206
rect 47762 44970 47804 45206
rect 81484 44970 81526 45206
rect 81762 44970 81804 45206
rect 6684 44032 6692 44096
rect 6756 44032 6772 44096
rect 6836 44032 6852 44096
rect 6916 44032 6932 44096
rect 6996 44032 7004 44096
rect 6684 43008 7004 44032
rect 6684 42944 6692 43008
rect 6756 42944 6772 43008
rect 6836 42944 6852 43008
rect 6916 42944 6932 43008
rect 6996 42944 7004 43008
rect 6684 41920 7004 42944
rect 6684 41856 6692 41920
rect 6756 41856 6772 41920
rect 6836 41856 6852 41920
rect 6916 41856 6932 41920
rect 6996 41856 7004 41920
rect 6684 40832 7004 41856
rect 6684 40768 6692 40832
rect 6756 40768 6772 40832
rect 6836 40768 6852 40832
rect 6916 40768 6932 40832
rect 6996 40768 7004 40832
rect 6684 39744 7004 40768
rect 6684 39680 6692 39744
rect 6756 39680 6772 39744
rect 6836 39680 6852 39744
rect 6916 39680 6932 39744
rect 6996 39680 7004 39744
rect 6684 38674 7004 39680
rect 87092 44640 87412 45664
rect 87092 44576 87100 44640
rect 87164 44576 87180 44640
rect 87244 44576 87260 44640
rect 87324 44576 87340 44640
rect 87404 44576 87412 44640
rect 87092 43552 87412 44576
rect 87092 43488 87100 43552
rect 87164 43488 87180 43552
rect 87244 43488 87260 43552
rect 87324 43488 87340 43552
rect 87404 43488 87412 43552
rect 87092 42464 87412 43488
rect 87092 42400 87100 42464
rect 87164 42400 87180 42464
rect 87244 42400 87260 42464
rect 87324 42400 87340 42464
rect 87404 42400 87412 42464
rect 87092 41376 87412 42400
rect 87092 41312 87100 41376
rect 87164 41312 87180 41376
rect 87244 41312 87260 41376
rect 87324 41312 87340 41376
rect 87404 41312 87412 41376
rect 87092 40288 87412 41312
rect 87092 40224 87100 40288
rect 87164 40224 87180 40288
rect 87244 40224 87260 40288
rect 87324 40224 87340 40288
rect 87404 40224 87412 40288
rect 87092 39200 87412 40224
rect 87092 39136 87100 39200
rect 87164 39136 87180 39200
rect 87244 39136 87260 39200
rect 87324 39136 87340 39200
rect 87404 39136 87412 39200
rect 6684 38656 6726 38674
rect 6962 38656 7004 38674
rect 6684 38592 6692 38656
rect 6996 38592 7004 38656
rect 6684 38438 6726 38592
rect 6962 38438 7004 38592
rect 11144 38438 11186 38674
rect 11422 38438 11464 38674
rect 45144 38438 45186 38674
rect 45422 38438 45464 38674
rect 48144 38438 48186 38674
rect 48422 38438 48464 38674
rect 82144 38438 82186 38674
rect 82422 38438 82464 38674
rect 6684 37568 7004 38438
rect 87092 38112 87412 39136
rect 87092 38048 87100 38112
rect 87164 38048 87180 38112
rect 87244 38048 87260 38112
rect 87324 38048 87340 38112
rect 87404 38048 87412 38112
rect 87092 38014 87412 38048
rect 10484 37778 10526 38014
rect 10762 37778 10804 38014
rect 44484 37778 44526 38014
rect 44762 37778 44804 38014
rect 47484 37778 47526 38014
rect 47762 37778 47804 38014
rect 81484 37778 81526 38014
rect 81762 37778 81804 38014
rect 87092 37778 87134 38014
rect 87370 37778 87412 38014
rect 6684 37504 6692 37568
rect 6756 37504 6772 37568
rect 6836 37504 6852 37568
rect 6916 37504 6932 37568
rect 6996 37504 7004 37568
rect 6684 36480 7004 37504
rect 6684 36416 6692 36480
rect 6756 36416 6772 36480
rect 6836 36416 6852 36480
rect 6916 36416 6932 36480
rect 6996 36416 7004 36480
rect 6684 35392 7004 36416
rect 6684 35328 6692 35392
rect 6756 35328 6772 35392
rect 6836 35328 6852 35392
rect 6916 35328 6932 35392
rect 6996 35328 7004 35392
rect 6684 34304 7004 35328
rect 6684 34240 6692 34304
rect 6756 34240 6772 34304
rect 6836 34240 6852 34304
rect 6916 34240 6932 34304
rect 6996 34240 7004 34304
rect 6684 33216 7004 34240
rect 6684 33152 6692 33216
rect 6756 33152 6772 33216
rect 6836 33152 6852 33216
rect 6916 33152 6932 33216
rect 6996 33152 7004 33216
rect 6684 32128 7004 33152
rect 6684 32064 6692 32128
rect 6756 32064 6772 32128
rect 6836 32064 6852 32128
rect 6916 32064 6932 32128
rect 6996 32064 7004 32128
rect 6684 31040 7004 32064
rect 6684 30976 6692 31040
rect 6756 30976 6772 31040
rect 6836 30976 6852 31040
rect 6916 30976 6932 31040
rect 6996 30976 7004 31040
rect 6684 29952 7004 30976
rect 6684 29888 6692 29952
rect 6756 29888 6772 29952
rect 6836 29888 6852 29952
rect 6916 29888 6932 29952
rect 6996 29888 7004 29952
rect 6684 28864 7004 29888
rect 6684 28800 6692 28864
rect 6756 28800 6772 28864
rect 6836 28800 6852 28864
rect 6916 28800 6932 28864
rect 6996 28800 7004 28864
rect 6684 27776 7004 28800
rect 6684 27712 6692 27776
rect 6756 27712 6772 27776
rect 6836 27712 6852 27776
rect 6916 27712 6932 27776
rect 6996 27712 7004 27776
rect 6684 26688 7004 27712
rect 6684 26624 6692 26688
rect 6756 26624 6772 26688
rect 6836 26624 6852 26688
rect 6916 26624 6932 26688
rect 6996 26624 7004 26688
rect 6684 25600 7004 26624
rect 6684 25536 6692 25600
rect 6756 25536 6772 25600
rect 6836 25536 6852 25600
rect 6916 25536 6932 25600
rect 6996 25536 7004 25600
rect 6684 24512 7004 25536
rect 6684 24448 6692 24512
rect 6756 24448 6772 24512
rect 6836 24448 6852 24512
rect 6916 24448 6932 24512
rect 6996 24448 7004 24512
rect 6684 23424 7004 24448
rect 6684 23360 6692 23424
rect 6756 23360 6772 23424
rect 6836 23360 6852 23424
rect 6916 23360 6932 23424
rect 6996 23360 7004 23424
rect 6684 22336 7004 23360
rect 6684 22272 6692 22336
rect 6756 22272 6772 22336
rect 6836 22272 6852 22336
rect 6916 22272 6932 22336
rect 6996 22272 7004 22336
rect 6684 21248 7004 22272
rect 6684 21184 6692 21248
rect 6756 21184 6772 21248
rect 6836 21184 6852 21248
rect 6916 21184 6932 21248
rect 6996 21184 7004 21248
rect 6684 20160 7004 21184
rect 6684 20096 6692 20160
rect 6756 20096 6772 20160
rect 6836 20096 6852 20160
rect 6916 20096 6932 20160
rect 6996 20096 7004 20160
rect 6684 19674 7004 20096
rect 87092 37024 87412 37778
rect 87092 36960 87100 37024
rect 87164 36960 87180 37024
rect 87244 36960 87260 37024
rect 87324 36960 87340 37024
rect 87404 36960 87412 37024
rect 87092 35936 87412 36960
rect 87092 35872 87100 35936
rect 87164 35872 87180 35936
rect 87244 35872 87260 35936
rect 87324 35872 87340 35936
rect 87404 35872 87412 35936
rect 87092 34848 87412 35872
rect 87092 34784 87100 34848
rect 87164 34784 87180 34848
rect 87244 34784 87260 34848
rect 87324 34784 87340 34848
rect 87404 34784 87412 34848
rect 87092 33760 87412 34784
rect 87092 33696 87100 33760
rect 87164 33696 87180 33760
rect 87244 33696 87260 33760
rect 87324 33696 87340 33760
rect 87404 33696 87412 33760
rect 87092 32672 87412 33696
rect 87092 32608 87100 32672
rect 87164 32608 87180 32672
rect 87244 32608 87260 32672
rect 87324 32608 87340 32672
rect 87404 32608 87412 32672
rect 87092 31584 87412 32608
rect 87092 31520 87100 31584
rect 87164 31520 87180 31584
rect 87244 31520 87260 31584
rect 87324 31520 87340 31584
rect 87404 31520 87412 31584
rect 87092 30496 87412 31520
rect 87092 30432 87100 30496
rect 87164 30432 87180 30496
rect 87244 30432 87260 30496
rect 87324 30432 87340 30496
rect 87404 30432 87412 30496
rect 87092 29408 87412 30432
rect 87092 29344 87100 29408
rect 87164 29344 87180 29408
rect 87244 29344 87260 29408
rect 87324 29344 87340 29408
rect 87404 29344 87412 29408
rect 87092 28320 87412 29344
rect 87092 28256 87100 28320
rect 87164 28256 87180 28320
rect 87244 28256 87260 28320
rect 87324 28256 87340 28320
rect 87404 28256 87412 28320
rect 87092 27232 87412 28256
rect 87092 27168 87100 27232
rect 87164 27168 87180 27232
rect 87244 27168 87260 27232
rect 87324 27168 87340 27232
rect 87404 27168 87412 27232
rect 87092 26144 87412 27168
rect 87092 26080 87100 26144
rect 87164 26080 87180 26144
rect 87244 26080 87260 26144
rect 87324 26080 87340 26144
rect 87404 26080 87412 26144
rect 87092 25056 87412 26080
rect 87092 24992 87100 25056
rect 87164 24992 87180 25056
rect 87244 24992 87260 25056
rect 87324 24992 87340 25056
rect 87404 24992 87412 25056
rect 87092 23968 87412 24992
rect 87092 23904 87100 23968
rect 87164 23904 87180 23968
rect 87244 23904 87260 23968
rect 87324 23904 87340 23968
rect 87404 23904 87412 23968
rect 87092 22880 87412 23904
rect 87092 22816 87100 22880
rect 87164 22816 87180 22880
rect 87244 22816 87260 22880
rect 87324 22816 87340 22880
rect 87404 22816 87412 22880
rect 87092 21792 87412 22816
rect 87092 21728 87100 21792
rect 87164 21728 87180 21792
rect 87244 21728 87260 21792
rect 87324 21728 87340 21792
rect 87404 21728 87412 21792
rect 87092 20704 87412 21728
rect 87092 20640 87100 20704
rect 87164 20640 87180 20704
rect 87244 20640 87260 20704
rect 87324 20640 87340 20704
rect 87404 20640 87412 20704
rect 6684 19438 6726 19674
rect 6962 19438 7004 19674
rect 11144 19438 11186 19674
rect 11422 19438 11464 19674
rect 45144 19438 45186 19674
rect 45422 19438 45464 19674
rect 48144 19438 48186 19674
rect 48422 19438 48464 19674
rect 82144 19438 82186 19674
rect 82422 19438 82464 19674
rect 87092 19616 87412 20640
rect 87092 19552 87100 19616
rect 87164 19552 87180 19616
rect 87244 19552 87260 19616
rect 87324 19552 87340 19616
rect 87404 19552 87412 19616
rect 6684 19072 7004 19438
rect 6684 19008 6692 19072
rect 6756 19008 6772 19072
rect 6836 19008 6852 19072
rect 6916 19008 6932 19072
rect 6996 19008 7004 19072
rect 87092 19014 87412 19552
rect 6684 17984 7004 19008
rect 10484 18778 10526 19014
rect 10762 18778 10804 19014
rect 44484 18778 44526 19014
rect 44762 18778 44804 19014
rect 47484 18778 47526 19014
rect 47762 18778 47804 19014
rect 81484 18778 81526 19014
rect 81762 18778 81804 19014
rect 87092 18778 87134 19014
rect 87370 18778 87412 19014
rect 6684 17920 6692 17984
rect 6756 17920 6772 17984
rect 6836 17920 6852 17984
rect 6916 17920 6932 17984
rect 6996 17920 7004 17984
rect 6684 16896 7004 17920
rect 6684 16832 6692 16896
rect 6756 16832 6772 16896
rect 6836 16832 6852 16896
rect 6916 16832 6932 16896
rect 6996 16832 7004 16896
rect 6684 15808 7004 16832
rect 6684 15744 6692 15808
rect 6756 15744 6772 15808
rect 6836 15744 6852 15808
rect 6916 15744 6932 15808
rect 6996 15744 7004 15808
rect 6684 14720 7004 15744
rect 6684 14656 6692 14720
rect 6756 14656 6772 14720
rect 6836 14656 6852 14720
rect 6916 14656 6932 14720
rect 6996 14656 7004 14720
rect 6684 13632 7004 14656
rect 6684 13568 6692 13632
rect 6756 13568 6772 13632
rect 6836 13568 6852 13632
rect 6916 13568 6932 13632
rect 6996 13568 7004 13632
rect 6684 12544 7004 13568
rect 6684 12480 6692 12544
rect 6756 12480 6772 12544
rect 6836 12480 6852 12544
rect 6916 12480 6932 12544
rect 6996 12480 7004 12544
rect 6684 11456 7004 12480
rect 87092 18528 87412 18778
rect 87092 18464 87100 18528
rect 87164 18464 87180 18528
rect 87244 18464 87260 18528
rect 87324 18464 87340 18528
rect 87404 18464 87412 18528
rect 87092 17440 87412 18464
rect 87092 17376 87100 17440
rect 87164 17376 87180 17440
rect 87244 17376 87260 17440
rect 87324 17376 87340 17440
rect 87404 17376 87412 17440
rect 87092 16352 87412 17376
rect 87092 16288 87100 16352
rect 87164 16288 87180 16352
rect 87244 16288 87260 16352
rect 87324 16288 87340 16352
rect 87404 16288 87412 16352
rect 87092 15264 87412 16288
rect 87092 15200 87100 15264
rect 87164 15200 87180 15264
rect 87244 15200 87260 15264
rect 87324 15200 87340 15264
rect 87404 15200 87412 15264
rect 87092 14176 87412 15200
rect 87092 14112 87100 14176
rect 87164 14112 87180 14176
rect 87244 14112 87260 14176
rect 87324 14112 87340 14176
rect 87404 14112 87412 14176
rect 87092 13088 87412 14112
rect 87092 13024 87100 13088
rect 87164 13024 87180 13088
rect 87244 13024 87260 13088
rect 87324 13024 87340 13088
rect 87404 13024 87412 13088
rect 87092 12000 87412 13024
rect 87092 11936 87100 12000
rect 87164 11936 87180 12000
rect 87244 11936 87260 12000
rect 87324 11936 87340 12000
rect 87404 11936 87412 12000
rect 11144 11630 11186 11866
rect 11422 11630 11464 11866
rect 45144 11630 45186 11866
rect 45422 11630 45464 11866
rect 48144 11630 48186 11866
rect 48422 11630 48464 11866
rect 82144 11630 82186 11866
rect 82422 11630 82464 11866
rect 6684 11392 6692 11456
rect 6756 11392 6772 11456
rect 6836 11392 6852 11456
rect 6916 11392 6932 11456
rect 6996 11392 7004 11456
rect 6684 10368 7004 11392
rect 10484 10970 10526 11206
rect 10762 10970 10804 11206
rect 44484 10970 44526 11206
rect 44762 10970 44804 11206
rect 47484 10970 47526 11206
rect 47762 10970 47804 11206
rect 81484 10970 81526 11206
rect 81762 10970 81804 11206
rect 6684 10304 6692 10368
rect 6756 10304 6772 10368
rect 6836 10304 6852 10368
rect 6916 10304 6932 10368
rect 6996 10304 7004 10368
rect 6684 9280 7004 10304
rect 6684 9216 6692 9280
rect 6756 9216 6772 9280
rect 6836 9216 6852 9280
rect 6916 9216 6932 9280
rect 6996 9216 7004 9280
rect 6684 8192 7004 9216
rect 87092 10912 87412 11936
rect 87092 10848 87100 10912
rect 87164 10848 87180 10912
rect 87244 10848 87260 10912
rect 87324 10848 87340 10912
rect 87404 10848 87412 10912
rect 87092 9824 87412 10848
rect 87092 9760 87100 9824
rect 87164 9760 87180 9824
rect 87244 9760 87260 9824
rect 87324 9760 87340 9824
rect 87404 9760 87412 9824
rect 6684 8128 6692 8192
rect 6756 8128 6772 8192
rect 6836 8128 6852 8192
rect 6916 8128 6932 8192
rect 6996 8128 7004 8192
rect 6684 7104 7004 8128
rect 6684 7040 6692 7104
rect 6756 7040 6772 7104
rect 6836 7040 6852 7104
rect 6916 7040 6932 7104
rect 6996 7040 7004 7104
rect 6684 7024 7004 7040
rect 18716 7648 19036 8927
rect 18716 7584 18724 7648
rect 18788 7584 18804 7648
rect 18868 7584 18884 7648
rect 18948 7584 18964 7648
rect 19028 7584 19036 7648
rect 3356 3418 3398 3654
rect 3634 3418 3676 3654
rect 3356 3376 3676 3418
rect 18716 6560 19036 7584
rect 18716 6496 18724 6560
rect 18788 6496 18804 6560
rect 18868 6496 18884 6560
rect 18948 6496 18964 6560
rect 19028 6496 19036 6560
rect 18716 5472 19036 6496
rect 18716 5408 18724 5472
rect 18788 5408 18804 5472
rect 18868 5408 18884 5472
rect 18948 5408 18964 5472
rect 19028 5408 19036 5472
rect 18716 3654 19036 5408
rect 18716 3418 18758 3654
rect 18994 3418 19036 3654
rect 2696 2758 2738 2994
rect 2974 2758 3016 2994
rect 2696 2716 3016 2758
rect 18716 2716 19036 3418
rect 19376 7104 19696 8927
rect 19376 7040 19384 7104
rect 19448 7040 19464 7104
rect 19528 7040 19544 7104
rect 19608 7040 19624 7104
rect 19688 7040 19696 7104
rect 19376 6016 19696 7040
rect 19376 5952 19384 6016
rect 19448 5952 19464 6016
rect 19528 5952 19544 6016
rect 19608 5952 19624 6016
rect 19688 5952 19696 6016
rect 19376 4928 19696 5952
rect 19376 4864 19384 4928
rect 19448 4864 19464 4928
rect 19528 4864 19544 4928
rect 19608 4864 19624 4928
rect 19688 4864 19696 4928
rect 19376 2994 19696 4864
rect 19376 2758 19418 2994
rect 19654 2758 19696 2994
rect 19376 2716 19696 2758
rect 37716 7648 38036 8927
rect 37716 7584 37724 7648
rect 37788 7584 37804 7648
rect 37868 7584 37884 7648
rect 37948 7584 37964 7648
rect 38028 7584 38036 7648
rect 37716 6560 38036 7584
rect 37716 6496 37724 6560
rect 37788 6496 37804 6560
rect 37868 6496 37884 6560
rect 37948 6496 37964 6560
rect 38028 6496 38036 6560
rect 37716 5472 38036 6496
rect 37716 5408 37724 5472
rect 37788 5408 37804 5472
rect 37868 5408 37884 5472
rect 37948 5408 37964 5472
rect 38028 5408 38036 5472
rect 37716 3654 38036 5408
rect 37716 3418 37758 3654
rect 37994 3418 38036 3654
rect 37716 2716 38036 3418
rect 38376 7104 38696 8927
rect 38376 7040 38384 7104
rect 38448 7040 38464 7104
rect 38528 7040 38544 7104
rect 38608 7040 38624 7104
rect 38688 7040 38696 7104
rect 38376 6016 38696 7040
rect 38376 5952 38384 6016
rect 38448 5952 38464 6016
rect 38528 5952 38544 6016
rect 38608 5952 38624 6016
rect 38688 5952 38696 6016
rect 38376 4928 38696 5952
rect 38376 4864 38384 4928
rect 38448 4864 38464 4928
rect 38528 4864 38544 4928
rect 38608 4864 38624 4928
rect 38688 4864 38696 4928
rect 38376 2994 38696 4864
rect 38376 2758 38418 2994
rect 38654 2758 38696 2994
rect 38376 2716 38696 2758
rect 56716 7648 57036 8927
rect 56716 7584 56724 7648
rect 56788 7584 56804 7648
rect 56868 7584 56884 7648
rect 56948 7584 56964 7648
rect 57028 7584 57036 7648
rect 56716 6560 57036 7584
rect 56716 6496 56724 6560
rect 56788 6496 56804 6560
rect 56868 6496 56884 6560
rect 56948 6496 56964 6560
rect 57028 6496 57036 6560
rect 56716 5472 57036 6496
rect 56716 5408 56724 5472
rect 56788 5408 56804 5472
rect 56868 5408 56884 5472
rect 56948 5408 56964 5472
rect 57028 5408 57036 5472
rect 56716 3654 57036 5408
rect 56716 3418 56758 3654
rect 56994 3418 57036 3654
rect 56716 2716 57036 3418
rect 57376 7104 57696 8927
rect 57376 7040 57384 7104
rect 57448 7040 57464 7104
rect 57528 7040 57544 7104
rect 57608 7040 57624 7104
rect 57688 7040 57696 7104
rect 57376 6016 57696 7040
rect 57376 5952 57384 6016
rect 57448 5952 57464 6016
rect 57528 5952 57544 6016
rect 57608 5952 57624 6016
rect 57688 5952 57696 6016
rect 57376 4928 57696 5952
rect 57376 4864 57384 4928
rect 57448 4864 57464 4928
rect 57528 4864 57544 4928
rect 57608 4864 57624 4928
rect 57688 4864 57696 4928
rect 57376 2994 57696 4864
rect 57376 2758 57418 2994
rect 57654 2758 57696 2994
rect 57376 2716 57696 2758
rect 75716 7648 76036 8927
rect 75716 7584 75724 7648
rect 75788 7584 75804 7648
rect 75868 7584 75884 7648
rect 75948 7584 75964 7648
rect 76028 7584 76036 7648
rect 75716 6560 76036 7584
rect 75716 6496 75724 6560
rect 75788 6496 75804 6560
rect 75868 6496 75884 6560
rect 75948 6496 75964 6560
rect 76028 6496 76036 6560
rect 75716 5472 76036 6496
rect 75716 5408 75724 5472
rect 75788 5408 75804 5472
rect 75868 5408 75884 5472
rect 75948 5408 75964 5472
rect 76028 5408 76036 5472
rect 75716 3654 76036 5408
rect 75716 3418 75758 3654
rect 75994 3418 76036 3654
rect 75716 2716 76036 3418
rect 76376 7104 76696 8927
rect 76376 7040 76384 7104
rect 76448 7040 76464 7104
rect 76528 7040 76544 7104
rect 76608 7040 76624 7104
rect 76688 7040 76696 7104
rect 76376 6016 76696 7040
rect 87092 8736 87412 9760
rect 87092 8672 87100 8736
rect 87164 8672 87180 8736
rect 87244 8672 87260 8736
rect 87324 8672 87340 8736
rect 87404 8672 87412 8736
rect 87092 7648 87412 8672
rect 87092 7584 87100 7648
rect 87164 7584 87180 7648
rect 87244 7584 87260 7648
rect 87324 7584 87340 7648
rect 87404 7584 87412 7648
rect 87092 7024 87412 7584
rect 87828 86528 88148 87088
rect 87828 86464 87836 86528
rect 87900 86464 87916 86528
rect 87980 86464 87996 86528
rect 88060 86464 88076 86528
rect 88140 86464 88148 86528
rect 87828 85440 88148 86464
rect 87828 85376 87836 85440
rect 87900 85376 87916 85440
rect 87980 85376 87996 85440
rect 88060 85376 88076 85440
rect 88140 85376 88148 85440
rect 87828 84352 88148 85376
rect 87828 84288 87836 84352
rect 87900 84288 87916 84352
rect 87980 84288 87996 84352
rect 88060 84288 88076 84352
rect 88140 84288 88148 84352
rect 87828 83264 88148 84288
rect 87828 83200 87836 83264
rect 87900 83200 87916 83264
rect 87980 83200 87996 83264
rect 88060 83200 88076 83264
rect 88140 83200 88148 83264
rect 87828 82176 88148 83200
rect 87828 82112 87836 82176
rect 87900 82112 87916 82176
rect 87980 82112 87996 82176
rect 88060 82112 88076 82176
rect 88140 82112 88148 82176
rect 87828 81088 88148 82112
rect 87828 81024 87836 81088
rect 87900 81024 87916 81088
rect 87980 81024 87996 81088
rect 88060 81024 88076 81088
rect 88140 81024 88148 81088
rect 87828 80000 88148 81024
rect 87828 79936 87836 80000
rect 87900 79936 87916 80000
rect 87980 79936 87996 80000
rect 88060 79936 88076 80000
rect 88140 79936 88148 80000
rect 87828 78912 88148 79936
rect 87828 78848 87836 78912
rect 87900 78848 87916 78912
rect 87980 78848 87996 78912
rect 88060 78848 88076 78912
rect 88140 78848 88148 78912
rect 87828 77824 88148 78848
rect 87828 77760 87836 77824
rect 87900 77760 87916 77824
rect 87980 77760 87996 77824
rect 88060 77760 88076 77824
rect 88140 77760 88148 77824
rect 87828 76736 88148 77760
rect 87828 76672 87836 76736
rect 87900 76674 87916 76736
rect 87980 76674 87996 76736
rect 88060 76674 88076 76736
rect 88140 76672 88148 76736
rect 87828 76438 87870 76672
rect 88106 76438 88148 76672
rect 87828 75648 88148 76438
rect 87828 75584 87836 75648
rect 87900 75584 87916 75648
rect 87980 75584 87996 75648
rect 88060 75584 88076 75648
rect 88140 75584 88148 75648
rect 87828 74560 88148 75584
rect 87828 74496 87836 74560
rect 87900 74496 87916 74560
rect 87980 74496 87996 74560
rect 88060 74496 88076 74560
rect 88140 74496 88148 74560
rect 87828 73472 88148 74496
rect 87828 73408 87836 73472
rect 87900 73408 87916 73472
rect 87980 73408 87996 73472
rect 88060 73408 88076 73472
rect 88140 73408 88148 73472
rect 87828 72384 88148 73408
rect 87828 72320 87836 72384
rect 87900 72320 87916 72384
rect 87980 72320 87996 72384
rect 88060 72320 88076 72384
rect 88140 72320 88148 72384
rect 87828 71296 88148 72320
rect 87828 71232 87836 71296
rect 87900 71232 87916 71296
rect 87980 71232 87996 71296
rect 88060 71232 88076 71296
rect 88140 71232 88148 71296
rect 87828 70208 88148 71232
rect 87828 70144 87836 70208
rect 87900 70144 87916 70208
rect 87980 70144 87996 70208
rect 88060 70144 88076 70208
rect 88140 70144 88148 70208
rect 87828 69120 88148 70144
rect 87828 69056 87836 69120
rect 87900 69056 87916 69120
rect 87980 69056 87996 69120
rect 88060 69056 88076 69120
rect 88140 69056 88148 69120
rect 87828 68032 88148 69056
rect 87828 67968 87836 68032
rect 87900 67968 87916 68032
rect 87980 67968 87996 68032
rect 88060 67968 88076 68032
rect 88140 67968 88148 68032
rect 87828 66944 88148 67968
rect 87828 66880 87836 66944
rect 87900 66880 87916 66944
rect 87980 66880 87996 66944
rect 88060 66880 88076 66944
rect 88140 66880 88148 66944
rect 87828 65856 88148 66880
rect 87828 65792 87836 65856
rect 87900 65792 87916 65856
rect 87980 65792 87996 65856
rect 88060 65792 88076 65856
rect 88140 65792 88148 65856
rect 87828 64768 88148 65792
rect 87828 64704 87836 64768
rect 87900 64704 87916 64768
rect 87980 64704 87996 64768
rect 88060 64704 88076 64768
rect 88140 64704 88148 64768
rect 87828 63680 88148 64704
rect 87828 63616 87836 63680
rect 87900 63616 87916 63680
rect 87980 63616 87996 63680
rect 88060 63616 88076 63680
rect 88140 63616 88148 63680
rect 87828 62592 88148 63616
rect 87828 62528 87836 62592
rect 87900 62528 87916 62592
rect 87980 62528 87996 62592
rect 88060 62528 88076 62592
rect 88140 62528 88148 62592
rect 87828 61504 88148 62528
rect 87828 61440 87836 61504
rect 87900 61440 87916 61504
rect 87980 61440 87996 61504
rect 88060 61440 88076 61504
rect 88140 61440 88148 61504
rect 87828 60416 88148 61440
rect 87828 60352 87836 60416
rect 87900 60352 87916 60416
rect 87980 60352 87996 60416
rect 88060 60352 88076 60416
rect 88140 60352 88148 60416
rect 87828 59328 88148 60352
rect 87828 59264 87836 59328
rect 87900 59264 87916 59328
rect 87980 59264 87996 59328
rect 88060 59264 88076 59328
rect 88140 59264 88148 59328
rect 87828 58240 88148 59264
rect 87828 58176 87836 58240
rect 87900 58176 87916 58240
rect 87980 58176 87996 58240
rect 88060 58176 88076 58240
rect 88140 58176 88148 58240
rect 87828 57674 88148 58176
rect 87828 57438 87870 57674
rect 88106 57438 88148 57674
rect 87828 57152 88148 57438
rect 87828 57088 87836 57152
rect 87900 57088 87916 57152
rect 87980 57088 87996 57152
rect 88060 57088 88076 57152
rect 88140 57088 88148 57152
rect 87828 56064 88148 57088
rect 87828 56000 87836 56064
rect 87900 56000 87916 56064
rect 87980 56000 87996 56064
rect 88060 56000 88076 56064
rect 88140 56000 88148 56064
rect 87828 54976 88148 56000
rect 87828 54912 87836 54976
rect 87900 54912 87916 54976
rect 87980 54912 87996 54976
rect 88060 54912 88076 54976
rect 88140 54912 88148 54976
rect 87828 53888 88148 54912
rect 87828 53824 87836 53888
rect 87900 53824 87916 53888
rect 87980 53824 87996 53888
rect 88060 53824 88076 53888
rect 88140 53824 88148 53888
rect 87828 52800 88148 53824
rect 87828 52736 87836 52800
rect 87900 52736 87916 52800
rect 87980 52736 87996 52800
rect 88060 52736 88076 52800
rect 88140 52736 88148 52800
rect 87828 51712 88148 52736
rect 87828 51648 87836 51712
rect 87900 51648 87916 51712
rect 87980 51648 87996 51712
rect 88060 51648 88076 51712
rect 88140 51648 88148 51712
rect 87828 50624 88148 51648
rect 87828 50560 87836 50624
rect 87900 50560 87916 50624
rect 87980 50560 87996 50624
rect 88060 50560 88076 50624
rect 88140 50560 88148 50624
rect 87828 49536 88148 50560
rect 87828 49472 87836 49536
rect 87900 49472 87916 49536
rect 87980 49472 87996 49536
rect 88060 49472 88076 49536
rect 88140 49472 88148 49536
rect 87828 48448 88148 49472
rect 87828 48384 87836 48448
rect 87900 48384 87916 48448
rect 87980 48384 87996 48448
rect 88060 48384 88076 48448
rect 88140 48384 88148 48448
rect 87828 47360 88148 48384
rect 87828 47296 87836 47360
rect 87900 47296 87916 47360
rect 87980 47296 87996 47360
rect 88060 47296 88076 47360
rect 88140 47296 88148 47360
rect 87828 46272 88148 47296
rect 87828 46208 87836 46272
rect 87900 46208 87916 46272
rect 87980 46208 87996 46272
rect 88060 46208 88076 46272
rect 88140 46208 88148 46272
rect 87828 45184 88148 46208
rect 87828 45120 87836 45184
rect 87900 45120 87916 45184
rect 87980 45120 87996 45184
rect 88060 45120 88076 45184
rect 88140 45120 88148 45184
rect 87828 44096 88148 45120
rect 87828 44032 87836 44096
rect 87900 44032 87916 44096
rect 87980 44032 87996 44096
rect 88060 44032 88076 44096
rect 88140 44032 88148 44096
rect 87828 43008 88148 44032
rect 87828 42944 87836 43008
rect 87900 42944 87916 43008
rect 87980 42944 87996 43008
rect 88060 42944 88076 43008
rect 88140 42944 88148 43008
rect 87828 41920 88148 42944
rect 87828 41856 87836 41920
rect 87900 41856 87916 41920
rect 87980 41856 87996 41920
rect 88060 41856 88076 41920
rect 88140 41856 88148 41920
rect 87828 40832 88148 41856
rect 87828 40768 87836 40832
rect 87900 40768 87916 40832
rect 87980 40768 87996 40832
rect 88060 40768 88076 40832
rect 88140 40768 88148 40832
rect 87828 39744 88148 40768
rect 87828 39680 87836 39744
rect 87900 39680 87916 39744
rect 87980 39680 87996 39744
rect 88060 39680 88076 39744
rect 88140 39680 88148 39744
rect 87828 38674 88148 39680
rect 87828 38656 87870 38674
rect 88106 38656 88148 38674
rect 87828 38592 87836 38656
rect 88140 38592 88148 38656
rect 87828 38438 87870 38592
rect 88106 38438 88148 38592
rect 87828 37568 88148 38438
rect 87828 37504 87836 37568
rect 87900 37504 87916 37568
rect 87980 37504 87996 37568
rect 88060 37504 88076 37568
rect 88140 37504 88148 37568
rect 87828 36480 88148 37504
rect 87828 36416 87836 36480
rect 87900 36416 87916 36480
rect 87980 36416 87996 36480
rect 88060 36416 88076 36480
rect 88140 36416 88148 36480
rect 87828 35392 88148 36416
rect 87828 35328 87836 35392
rect 87900 35328 87916 35392
rect 87980 35328 87996 35392
rect 88060 35328 88076 35392
rect 88140 35328 88148 35392
rect 87828 34304 88148 35328
rect 87828 34240 87836 34304
rect 87900 34240 87916 34304
rect 87980 34240 87996 34304
rect 88060 34240 88076 34304
rect 88140 34240 88148 34304
rect 87828 33216 88148 34240
rect 87828 33152 87836 33216
rect 87900 33152 87916 33216
rect 87980 33152 87996 33216
rect 88060 33152 88076 33216
rect 88140 33152 88148 33216
rect 87828 32128 88148 33152
rect 87828 32064 87836 32128
rect 87900 32064 87916 32128
rect 87980 32064 87996 32128
rect 88060 32064 88076 32128
rect 88140 32064 88148 32128
rect 87828 31040 88148 32064
rect 87828 30976 87836 31040
rect 87900 30976 87916 31040
rect 87980 30976 87996 31040
rect 88060 30976 88076 31040
rect 88140 30976 88148 31040
rect 87828 29952 88148 30976
rect 87828 29888 87836 29952
rect 87900 29888 87916 29952
rect 87980 29888 87996 29952
rect 88060 29888 88076 29952
rect 88140 29888 88148 29952
rect 87828 28864 88148 29888
rect 87828 28800 87836 28864
rect 87900 28800 87916 28864
rect 87980 28800 87996 28864
rect 88060 28800 88076 28864
rect 88140 28800 88148 28864
rect 87828 27776 88148 28800
rect 87828 27712 87836 27776
rect 87900 27712 87916 27776
rect 87980 27712 87996 27776
rect 88060 27712 88076 27776
rect 88140 27712 88148 27776
rect 87828 26688 88148 27712
rect 87828 26624 87836 26688
rect 87900 26624 87916 26688
rect 87980 26624 87996 26688
rect 88060 26624 88076 26688
rect 88140 26624 88148 26688
rect 87828 25600 88148 26624
rect 87828 25536 87836 25600
rect 87900 25536 87916 25600
rect 87980 25536 87996 25600
rect 88060 25536 88076 25600
rect 88140 25536 88148 25600
rect 87828 24512 88148 25536
rect 87828 24448 87836 24512
rect 87900 24448 87916 24512
rect 87980 24448 87996 24512
rect 88060 24448 88076 24512
rect 88140 24448 88148 24512
rect 87828 23424 88148 24448
rect 87828 23360 87836 23424
rect 87900 23360 87916 23424
rect 87980 23360 87996 23424
rect 88060 23360 88076 23424
rect 88140 23360 88148 23424
rect 87828 22336 88148 23360
rect 87828 22272 87836 22336
rect 87900 22272 87916 22336
rect 87980 22272 87996 22336
rect 88060 22272 88076 22336
rect 88140 22272 88148 22336
rect 87828 21248 88148 22272
rect 87828 21184 87836 21248
rect 87900 21184 87916 21248
rect 87980 21184 87996 21248
rect 88060 21184 88076 21248
rect 88140 21184 88148 21248
rect 87828 20160 88148 21184
rect 87828 20096 87836 20160
rect 87900 20096 87916 20160
rect 87980 20096 87996 20160
rect 88060 20096 88076 20160
rect 88140 20096 88148 20160
rect 87828 19674 88148 20096
rect 87828 19438 87870 19674
rect 88106 19438 88148 19674
rect 87828 19072 88148 19438
rect 87828 19008 87836 19072
rect 87900 19008 87916 19072
rect 87980 19008 87996 19072
rect 88060 19008 88076 19072
rect 88140 19008 88148 19072
rect 87828 17984 88148 19008
rect 87828 17920 87836 17984
rect 87900 17920 87916 17984
rect 87980 17920 87996 17984
rect 88060 17920 88076 17984
rect 88140 17920 88148 17984
rect 87828 16896 88148 17920
rect 87828 16832 87836 16896
rect 87900 16832 87916 16896
rect 87980 16832 87996 16896
rect 88060 16832 88076 16896
rect 88140 16832 88148 16896
rect 87828 15808 88148 16832
rect 87828 15744 87836 15808
rect 87900 15744 87916 15808
rect 87980 15744 87996 15808
rect 88060 15744 88076 15808
rect 88140 15744 88148 15808
rect 87828 14720 88148 15744
rect 87828 14656 87836 14720
rect 87900 14656 87916 14720
rect 87980 14656 87996 14720
rect 88060 14656 88076 14720
rect 88140 14656 88148 14720
rect 87828 13632 88148 14656
rect 87828 13568 87836 13632
rect 87900 13568 87916 13632
rect 87980 13568 87996 13632
rect 88060 13568 88076 13632
rect 88140 13568 88148 13632
rect 87828 12544 88148 13568
rect 87828 12480 87836 12544
rect 87900 12480 87916 12544
rect 87980 12480 87996 12544
rect 88060 12480 88076 12544
rect 88140 12480 88148 12544
rect 87828 11456 88148 12480
rect 87828 11392 87836 11456
rect 87900 11392 87916 11456
rect 87980 11392 87996 11456
rect 88060 11392 88076 11456
rect 88140 11392 88148 11456
rect 87828 10368 88148 11392
rect 87828 10304 87836 10368
rect 87900 10304 87916 10368
rect 87980 10304 87996 10368
rect 88060 10304 88076 10368
rect 88140 10304 88148 10368
rect 87828 9280 88148 10304
rect 87828 9216 87836 9280
rect 87900 9216 87916 9280
rect 87980 9216 87996 9280
rect 88060 9216 88076 9280
rect 88140 9216 88148 9280
rect 87828 8192 88148 9216
rect 87828 8128 87836 8192
rect 87900 8128 87916 8192
rect 87980 8128 87996 8192
rect 88060 8128 88076 8192
rect 88140 8128 88148 8192
rect 87828 7104 88148 8128
rect 87828 7040 87836 7104
rect 87900 7040 87916 7104
rect 87980 7040 87996 7104
rect 88060 7040 88076 7104
rect 88140 7040 88148 7104
rect 87828 7024 88148 7040
rect 90164 76014 90484 90458
rect 90164 75778 90206 76014
rect 90442 75778 90484 76014
rect 90164 57014 90484 75778
rect 90164 56778 90206 57014
rect 90442 56778 90484 57014
rect 90164 38014 90484 56778
rect 90164 37778 90206 38014
rect 90442 37778 90484 38014
rect 90164 19014 90484 37778
rect 90164 18778 90206 19014
rect 90442 18778 90484 19014
rect 76376 5952 76384 6016
rect 76448 5952 76464 6016
rect 76528 5952 76544 6016
rect 76608 5952 76624 6016
rect 76688 5952 76696 6016
rect 76376 4928 76696 5952
rect 76376 4864 76384 4928
rect 76448 4864 76464 4928
rect 76528 4864 76544 4928
rect 76608 4864 76624 4928
rect 76688 4864 76696 4928
rect 76376 2994 76696 4864
rect 90164 3654 90484 18778
rect 90164 3418 90206 3654
rect 90442 3418 90484 3654
rect 90164 3376 90484 3418
rect 90824 76674 91144 91118
rect 90824 76438 90866 76674
rect 91102 76438 91144 76674
rect 90824 57674 91144 76438
rect 90824 57438 90866 57674
rect 91102 57438 91144 57674
rect 90824 38674 91144 57438
rect 90824 38438 90866 38674
rect 91102 38438 91144 38674
rect 90824 19674 91144 38438
rect 90824 19438 90866 19674
rect 91102 19438 91144 19674
rect 76376 2758 76418 2994
rect 76654 2758 76696 2994
rect 76376 2716 76696 2758
rect 90824 2994 91144 19438
rect 90824 2758 90866 2994
rect 91102 2758 91144 2994
rect 90824 2716 91144 2758
<< via4 >>
rect 2738 91118 2974 91354
rect 2738 76438 2974 76674
rect 2738 57438 2974 57674
rect 2738 38438 2974 38674
rect 2738 19438 2974 19674
rect 3398 90458 3634 90694
rect 18758 90458 18994 90694
rect 3398 75778 3634 76014
rect 3398 56778 3634 57014
rect 3398 37778 3634 38014
rect 3398 18778 3634 19014
rect 5990 75778 6226 76014
rect 5990 56778 6226 57014
rect 5990 37778 6226 38014
rect 5990 18778 6226 19014
rect 19418 91118 19654 91354
rect 37758 90458 37994 90694
rect 38418 91118 38654 91354
rect 56758 90458 56994 90694
rect 57418 91118 57654 91354
rect 75758 90458 75994 90694
rect 76418 91118 76654 91354
rect 90866 91118 91102 91354
rect 90206 90458 90442 90694
rect 11186 83030 11422 83266
rect 45186 83030 45422 83266
rect 48186 83030 48422 83266
rect 82186 83030 82422 83266
rect 10526 82370 10762 82606
rect 44526 82370 44762 82606
rect 47526 82370 47762 82606
rect 81526 82370 81762 82606
rect 6726 76672 6756 76674
rect 6756 76672 6772 76674
rect 6772 76672 6836 76674
rect 6836 76672 6852 76674
rect 6852 76672 6916 76674
rect 6916 76672 6932 76674
rect 6932 76672 6962 76674
rect 6726 76438 6962 76672
rect 11186 76438 11422 76674
rect 45186 76438 45422 76674
rect 48186 76438 48422 76674
rect 82186 76438 82422 76674
rect 10526 75778 10762 76014
rect 44526 75778 44762 76014
rect 47526 75778 47762 76014
rect 81526 75778 81762 76014
rect 87134 75778 87370 76014
rect 6726 57438 6962 57674
rect 11186 57438 11422 57674
rect 45186 57438 45422 57674
rect 48186 57438 48422 57674
rect 82186 57438 82422 57674
rect 10526 56778 10762 57014
rect 44526 56778 44762 57014
rect 47526 56778 47762 57014
rect 81526 56778 81762 57014
rect 87134 56778 87370 57014
rect 11186 49030 11422 49266
rect 45186 49030 45422 49266
rect 48186 49030 48422 49266
rect 82186 49030 82422 49266
rect 10526 48370 10762 48606
rect 44526 48370 44762 48606
rect 47526 48370 47762 48606
rect 81526 48370 81762 48606
rect 11186 45630 11422 45866
rect 45186 45630 45422 45866
rect 48186 45630 48422 45866
rect 82186 45630 82422 45866
rect 10526 44970 10762 45206
rect 44526 44970 44762 45206
rect 47526 44970 47762 45206
rect 81526 44970 81762 45206
rect 6726 38656 6962 38674
rect 6726 38592 6756 38656
rect 6756 38592 6772 38656
rect 6772 38592 6836 38656
rect 6836 38592 6852 38656
rect 6852 38592 6916 38656
rect 6916 38592 6932 38656
rect 6932 38592 6962 38656
rect 6726 38438 6962 38592
rect 11186 38438 11422 38674
rect 45186 38438 45422 38674
rect 48186 38438 48422 38674
rect 82186 38438 82422 38674
rect 10526 37778 10762 38014
rect 44526 37778 44762 38014
rect 47526 37778 47762 38014
rect 81526 37778 81762 38014
rect 87134 37778 87370 38014
rect 6726 19438 6962 19674
rect 11186 19438 11422 19674
rect 45186 19438 45422 19674
rect 48186 19438 48422 19674
rect 82186 19438 82422 19674
rect 10526 18778 10762 19014
rect 44526 18778 44762 19014
rect 47526 18778 47762 19014
rect 81526 18778 81762 19014
rect 87134 18778 87370 19014
rect 11186 11630 11422 11866
rect 45186 11630 45422 11866
rect 48186 11630 48422 11866
rect 82186 11630 82422 11866
rect 10526 10970 10762 11206
rect 44526 10970 44762 11206
rect 47526 10970 47762 11206
rect 81526 10970 81762 11206
rect 3398 3418 3634 3654
rect 18758 3418 18994 3654
rect 2738 2758 2974 2994
rect 19418 2758 19654 2994
rect 37758 3418 37994 3654
rect 38418 2758 38654 2994
rect 56758 3418 56994 3654
rect 57418 2758 57654 2994
rect 75758 3418 75994 3654
rect 87870 76672 87900 76674
rect 87900 76672 87916 76674
rect 87916 76672 87980 76674
rect 87980 76672 87996 76674
rect 87996 76672 88060 76674
rect 88060 76672 88076 76674
rect 88076 76672 88106 76674
rect 87870 76438 88106 76672
rect 87870 57438 88106 57674
rect 87870 38656 88106 38674
rect 87870 38592 87900 38656
rect 87900 38592 87916 38656
rect 87916 38592 87980 38656
rect 87980 38592 87996 38656
rect 87996 38592 88060 38656
rect 88060 38592 88076 38656
rect 88076 38592 88106 38656
rect 87870 38438 88106 38592
rect 87870 19438 88106 19674
rect 90206 75778 90442 76014
rect 90206 56778 90442 57014
rect 90206 37778 90442 38014
rect 90206 18778 90442 19014
rect 90206 3418 90442 3654
rect 90866 76438 91102 76674
rect 90866 57438 91102 57674
rect 90866 38438 91102 38674
rect 90866 19438 91102 19674
rect 76418 2758 76654 2994
rect 90866 2758 91102 2994
<< metal5 >>
rect 2696 91354 91144 91396
rect 2696 91118 2738 91354
rect 2974 91118 19418 91354
rect 19654 91118 38418 91354
rect 38654 91118 57418 91354
rect 57654 91118 76418 91354
rect 76654 91118 90866 91354
rect 91102 91118 91144 91354
rect 2696 91076 91144 91118
rect 3356 90694 90484 90736
rect 3356 90458 3398 90694
rect 3634 90458 18758 90694
rect 18994 90458 37758 90694
rect 37994 90458 56758 90694
rect 56994 90458 75758 90694
rect 75994 90458 90206 90694
rect 90442 90458 90484 90694
rect 3356 90416 90484 90458
rect 11162 83266 11446 83308
rect 11162 83030 11186 83266
rect 11422 83030 11446 83266
rect 11162 82988 11446 83030
rect 45162 83266 45446 83308
rect 45162 83030 45186 83266
rect 45422 83030 45446 83266
rect 45162 82988 45446 83030
rect 48162 83266 48446 83308
rect 48162 83030 48186 83266
rect 48422 83030 48446 83266
rect 48162 82988 48446 83030
rect 82162 83266 82446 83308
rect 82162 83030 82186 83266
rect 82422 83030 82446 83266
rect 82162 82988 82446 83030
rect 10502 82606 10786 82648
rect 10502 82370 10526 82606
rect 10762 82370 10786 82606
rect 10502 82328 10786 82370
rect 44502 82606 44786 82648
rect 44502 82370 44526 82606
rect 44762 82370 44786 82606
rect 44502 82328 44786 82370
rect 47502 82606 47786 82648
rect 47502 82370 47526 82606
rect 47762 82370 47786 82606
rect 47502 82328 47786 82370
rect 81502 82606 81786 82648
rect 81502 82370 81526 82606
rect 81762 82370 81786 82606
rect 81502 82328 81786 82370
rect 2696 76674 91144 76716
rect 2696 76438 2738 76674
rect 2974 76438 6726 76674
rect 6962 76438 11186 76674
rect 11422 76438 45186 76674
rect 45422 76438 48186 76674
rect 48422 76438 82186 76674
rect 82422 76438 87870 76674
rect 88106 76438 90866 76674
rect 91102 76438 91144 76674
rect 2696 76396 91144 76438
rect 2696 76014 91144 76056
rect 2696 75778 3398 76014
rect 3634 75778 5990 76014
rect 6226 75778 10526 76014
rect 10762 75778 44526 76014
rect 44762 75778 47526 76014
rect 47762 75778 81526 76014
rect 81762 75778 87134 76014
rect 87370 75778 90206 76014
rect 90442 75778 91144 76014
rect 2696 75736 91144 75778
rect 2696 57674 91144 57716
rect 2696 57438 2738 57674
rect 2974 57438 6726 57674
rect 6962 57438 11186 57674
rect 11422 57438 45186 57674
rect 45422 57438 48186 57674
rect 48422 57438 82186 57674
rect 82422 57438 87870 57674
rect 88106 57438 90866 57674
rect 91102 57438 91144 57674
rect 2696 57396 91144 57438
rect 2696 57014 91144 57056
rect 2696 56778 3398 57014
rect 3634 56778 5990 57014
rect 6226 56778 10526 57014
rect 10762 56778 44526 57014
rect 44762 56778 47526 57014
rect 47762 56778 81526 57014
rect 81762 56778 87134 57014
rect 87370 56778 90206 57014
rect 90442 56778 91144 57014
rect 2696 56736 91144 56778
rect 11162 49266 11446 49308
rect 11162 49030 11186 49266
rect 11422 49030 11446 49266
rect 11162 48988 11446 49030
rect 45162 49266 45446 49308
rect 45162 49030 45186 49266
rect 45422 49030 45446 49266
rect 45162 48988 45446 49030
rect 48162 49266 48446 49308
rect 48162 49030 48186 49266
rect 48422 49030 48446 49266
rect 48162 48988 48446 49030
rect 82162 49266 82446 49308
rect 82162 49030 82186 49266
rect 82422 49030 82446 49266
rect 82162 48988 82446 49030
rect 10502 48606 10786 48648
rect 10502 48370 10526 48606
rect 10762 48370 10786 48606
rect 10502 48328 10786 48370
rect 44502 48606 44786 48648
rect 44502 48370 44526 48606
rect 44762 48370 44786 48606
rect 44502 48328 44786 48370
rect 47502 48606 47786 48648
rect 47502 48370 47526 48606
rect 47762 48370 47786 48606
rect 47502 48328 47786 48370
rect 81502 48606 81786 48648
rect 81502 48370 81526 48606
rect 81762 48370 81786 48606
rect 81502 48328 81786 48370
rect 11162 45866 11446 45908
rect 11162 45630 11186 45866
rect 11422 45630 11446 45866
rect 11162 45588 11446 45630
rect 45162 45866 45446 45908
rect 45162 45630 45186 45866
rect 45422 45630 45446 45866
rect 45162 45588 45446 45630
rect 48162 45866 48446 45908
rect 48162 45630 48186 45866
rect 48422 45630 48446 45866
rect 48162 45588 48446 45630
rect 82162 45866 82446 45908
rect 82162 45630 82186 45866
rect 82422 45630 82446 45866
rect 82162 45588 82446 45630
rect 10502 45206 10786 45248
rect 10502 44970 10526 45206
rect 10762 44970 10786 45206
rect 10502 44928 10786 44970
rect 44502 45206 44786 45248
rect 44502 44970 44526 45206
rect 44762 44970 44786 45206
rect 44502 44928 44786 44970
rect 47502 45206 47786 45248
rect 47502 44970 47526 45206
rect 47762 44970 47786 45206
rect 47502 44928 47786 44970
rect 81502 45206 81786 45248
rect 81502 44970 81526 45206
rect 81762 44970 81786 45206
rect 81502 44928 81786 44970
rect 2696 38674 91144 38716
rect 2696 38438 2738 38674
rect 2974 38438 6726 38674
rect 6962 38438 11186 38674
rect 11422 38438 45186 38674
rect 45422 38438 48186 38674
rect 48422 38438 82186 38674
rect 82422 38438 87870 38674
rect 88106 38438 90866 38674
rect 91102 38438 91144 38674
rect 2696 38396 91144 38438
rect 2696 38014 91144 38056
rect 2696 37778 3398 38014
rect 3634 37778 5990 38014
rect 6226 37778 10526 38014
rect 10762 37778 44526 38014
rect 44762 37778 47526 38014
rect 47762 37778 81526 38014
rect 81762 37778 87134 38014
rect 87370 37778 90206 38014
rect 90442 37778 91144 38014
rect 2696 37736 91144 37778
rect 2696 19674 91144 19716
rect 2696 19438 2738 19674
rect 2974 19438 6726 19674
rect 6962 19438 11186 19674
rect 11422 19438 45186 19674
rect 45422 19438 48186 19674
rect 48422 19438 82186 19674
rect 82422 19438 87870 19674
rect 88106 19438 90866 19674
rect 91102 19438 91144 19674
rect 2696 19396 91144 19438
rect 2696 19014 91144 19056
rect 2696 18778 3398 19014
rect 3634 18778 5990 19014
rect 6226 18778 10526 19014
rect 10762 18778 44526 19014
rect 44762 18778 47526 19014
rect 47762 18778 81526 19014
rect 81762 18778 87134 19014
rect 87370 18778 90206 19014
rect 90442 18778 91144 19014
rect 2696 18736 91144 18778
rect 11162 11866 11446 11908
rect 11162 11630 11186 11866
rect 11422 11630 11446 11866
rect 11162 11588 11446 11630
rect 45162 11866 45446 11908
rect 45162 11630 45186 11866
rect 45422 11630 45446 11866
rect 45162 11588 45446 11630
rect 48162 11866 48446 11908
rect 48162 11630 48186 11866
rect 48422 11630 48446 11866
rect 48162 11588 48446 11630
rect 82162 11866 82446 11908
rect 82162 11630 82186 11866
rect 82422 11630 82446 11866
rect 82162 11588 82446 11630
rect 10502 11206 10786 11248
rect 10502 10970 10526 11206
rect 10762 10970 10786 11206
rect 10502 10928 10786 10970
rect 44502 11206 44786 11248
rect 44502 10970 44526 11206
rect 44762 10970 44786 11206
rect 44502 10928 44786 10970
rect 47502 11206 47786 11248
rect 47502 10970 47526 11206
rect 47762 10970 47786 11206
rect 47502 10928 47786 10970
rect 81502 11206 81786 11248
rect 81502 10970 81526 11206
rect 81762 10970 81786 11206
rect 81502 10928 81786 10970
rect 3356 3654 90484 3696
rect 3356 3418 3398 3654
rect 3634 3418 18758 3654
rect 18994 3418 37758 3654
rect 37994 3418 56758 3654
rect 56994 3418 75758 3654
rect 75994 3418 90206 3654
rect 90442 3418 90484 3654
rect 3356 3376 90484 3418
rect 2696 2994 91144 3036
rect 2696 2758 2738 2994
rect 2974 2758 19418 2994
rect 19654 2758 38418 2994
rect 38654 2758 57418 2994
rect 57654 2758 76418 2994
rect 76654 2758 90866 2994
rect 91102 2758 91144 2994
rect 2696 2716 91144 2758
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 18001
transform 1 0 88136 0 -1 48416
box -38 -48 222 592
use fpgacell  cell0
timestamp 0
transform 1 0 10000 0 1 10000
box 0 0 37000 37000
use fpgacell  cell1
timestamp 0
transform 1 0 47000 0 1 10000
box 0 0 37000 37000
use fpgacell  cell2
timestamp 0
transform 1 0 10000 0 1 47400
box 0 0 37000 37000
use fpgacell  cell3
timestamp 0
transform 1 0 47000 0 1 47400
box 0 0 37000 37000
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 18001
transform -1 0 30636 0 1 86496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 18001
transform -1 0 7636 0 -1 54944
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 18001
transform 1 0 30728 0 1 86496
box -38 -48 1878 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3
timestamp 1636986456
transform 1 0 5152 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1636986456
transform 1 0 6256 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp 18001
transform 1 0 7360 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1636986456
transform 1 0 7544 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1636986456
transform 1 0 8648 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp 18001
transform 1 0 9752 0 1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1636986456
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1636986456
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 18001
transform 1 0 12328 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_96
timestamp 18001
transform 1 0 13708 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 18001
transform 1 0 14904 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_123
timestamp 18001
transform 1 0 16192 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_130
timestamp 18001
transform 1 0 16836 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 18001
transform 1 0 17572 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_145
timestamp 18001
transform 1 0 18216 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_153
timestamp 18001
transform 1 0 18952 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_158
timestamp 18001
transform 1 0 19412 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 18001
transform 1 0 20056 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_169
timestamp 18001
transform 1 0 20424 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_179
timestamp 18001
transform 1 0 21344 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_187
timestamp 18001
transform 1 0 22080 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 18001
transform 1 0 22632 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_197
timestamp 18001
transform 1 0 23000 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_207
timestamp 18001
transform 1 0 23920 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_214
timestamp 18001
transform 1 0 24564 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 18001
transform 1 0 25300 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_229
timestamp 18001
transform 1 0 25944 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_237
timestamp 18001
transform 1 0 26680 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_242
timestamp 18001
transform 1 0 27140 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 18001
transform 1 0 27784 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_253
timestamp 18001
transform 1 0 28152 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_263
timestamp 18001
transform 1 0 29072 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_271
timestamp 18001
transform 1 0 29808 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 18001
transform 1 0 30360 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_281
timestamp 18001
transform 1 0 30728 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_290
timestamp 18001
transform 1 0 31556 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_297
timestamp 18001
transform 1 0 32200 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 18001
transform 1 0 32936 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_312
timestamp 18001
transform 1 0 33580 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_320
timestamp 18001
transform 1 0 34316 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_325
timestamp 18001
transform 1 0 34776 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_332
timestamp 18001
transform 1 0 35420 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_337
timestamp 18001
transform 1 0 35880 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_346
timestamp 18001
transform 1 0 36708 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_354
timestamp 18001
transform 1 0 37444 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_360
timestamp 18001
transform 1 0 37996 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_365
timestamp 18001
transform 1 0 38456 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_374
timestamp 18001
transform 1 0 39284 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_381
timestamp 18001
transform 1 0 39928 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_389
timestamp 18001
transform 1 0 40664 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_396
timestamp 18001
transform 1 0 41308 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_404
timestamp 18001
transform 1 0 42044 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_410
timestamp 18001
transform 1 0 42596 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_417
timestamp 18001
transform 1 0 43240 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_421
timestamp 18001
transform 1 0 43608 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_437
timestamp 18001
transform 1 0 45080 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_445
timestamp 18001
transform 1 0 45816 0 1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_459
timestamp 1636986456
transform 1 0 47104 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_471
timestamp 18001
transform 1 0 48208 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_475
timestamp 18001
transform 1 0 48576 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_477
timestamp 1636986456
transform 1 0 48760 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_489
timestamp 1636986456
transform 1 0 49864 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_501
timestamp 18001
transform 1 0 50968 0 1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_505
timestamp 1636986456
transform 1 0 51336 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_517
timestamp 18001
transform 1 0 52440 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_522
timestamp 18001
transform 1 0 52900 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_530
timestamp 18001
transform 1 0 53636 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_537
timestamp 18001
transform 1 0 54280 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_543
timestamp 18001
transform 1 0 54832 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_551
timestamp 18001
transform 1 0 55568 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_557
timestamp 18001
transform 1 0 56120 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_561
timestamp 18001
transform 1 0 56488 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_571
timestamp 18001
transform 1 0 57408 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_579
timestamp 18001
transform 1 0 58144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_585
timestamp 18001
transform 1 0 58696 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_593
timestamp 18001
transform 1 0 59432 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_601
timestamp 18001
transform 1 0 60168 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_606
timestamp 18001
transform 1 0 60628 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_614
timestamp 18001
transform 1 0 61364 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_621
timestamp 18001
transform 1 0 62008 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_627
timestamp 18001
transform 1 0 62560 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_635
timestamp 18001
transform 1 0 63296 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_641
timestamp 18001
transform 1 0 63848 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_645
timestamp 18001
transform 1 0 64216 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_655
timestamp 18001
transform 1 0 65136 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_663
timestamp 18001
transform 1 0 65872 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_669
timestamp 18001
transform 1 0 66424 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_677
timestamp 18001
transform 1 0 67160 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_685
timestamp 18001
transform 1 0 67896 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_689
timestamp 18001
transform 1 0 68264 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_697
timestamp 18001
transform 1 0 69000 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_704
timestamp 18001
transform 1 0 69644 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_710
timestamp 18001
transform 1 0 70196 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_718
timestamp 18001
transform 1 0 70932 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_724
timestamp 18001
transform 1 0 71484 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_729
timestamp 18001
transform 1 0 71944 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_738
timestamp 18001
transform 1 0 72772 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_746
timestamp 18001
transform 1 0 73508 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_752
timestamp 18001
transform 1 0 74060 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_760
timestamp 18001
transform 1 0 74796 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_768
timestamp 18001
transform 1 0 75532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_773
timestamp 18001
transform 1 0 75992 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_781
timestamp 18001
transform 1 0 76728 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_788
timestamp 18001
transform 1 0 77372 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_794
timestamp 18001
transform 1 0 77924 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_802
timestamp 18001
transform 1 0 78660 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_809
timestamp 18001
transform 1 0 79304 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_813
timestamp 18001
transform 1 0 79672 0 1 4896
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_823
timestamp 1636986456
transform 1 0 80592 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_835
timestamp 18001
transform 1 0 81696 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_839
timestamp 18001
transform 1 0 82064 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_851
timestamp 1636986456
transform 1 0 83168 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_863
timestamp 18001
transform 1 0 84272 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_867
timestamp 18001
transform 1 0 84640 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_869
timestamp 1636986456
transform 1 0 84824 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_881
timestamp 1636986456
transform 1 0 85928 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_893
timestamp 18001
transform 1 0 87032 0 1 4896
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_897
timestamp 1636986456
transform 1 0 87400 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_909
timestamp 18001
transform 1 0 88504 0 1 4896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1636986456
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1636986456
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1636986456
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1636986456
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 18001
transform 1 0 9568 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 18001
transform 1 0 9936 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1636986456
transform 1 0 10120 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1636986456
transform 1 0 11224 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1636986456
transform 1 0 12328 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1636986456
transform 1 0 13432 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 18001
transform 1 0 14536 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 18001
transform 1 0 15088 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1636986456
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1636986456
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1636986456
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1636986456
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 18001
transform 1 0 19688 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 18001
transform 1 0 20240 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1636986456
transform 1 0 20424 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1636986456
transform 1 0 21528 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1636986456
transform 1 0 22632 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1636986456
transform 1 0 23736 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 18001
transform 1 0 24840 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 18001
transform 1 0 25392 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1636986456
transform 1 0 25576 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1636986456
transform 1 0 26680 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1636986456
transform 1 0 27784 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1636986456
transform 1 0 28888 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 18001
transform 1 0 29992 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 18001
transform 1 0 30544 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1636986456
transform 1 0 30728 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1636986456
transform 1 0 31832 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1636986456
transform 1 0 32936 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1636986456
transform 1 0 34040 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 18001
transform 1 0 35144 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 18001
transform 1 0 35696 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1636986456
transform 1 0 35880 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1636986456
transform 1 0 36984 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1636986456
transform 1 0 38088 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1636986456
transform 1 0 39192 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 18001
transform 1 0 40296 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 18001
transform 1 0 40848 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1636986456
transform 1 0 41032 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_405
timestamp 1636986456
transform 1 0 42136 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_417
timestamp 1636986456
transform 1 0 43240 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_429
timestamp 1636986456
transform 1 0 44344 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 18001
transform 1 0 45448 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 18001
transform 1 0 46000 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_449
timestamp 1636986456
transform 1 0 46184 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_461
timestamp 1636986456
transform 1 0 47288 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_473
timestamp 1636986456
transform 1 0 48392 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_485
timestamp 1636986456
transform 1 0 49496 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_497
timestamp 18001
transform 1 0 50600 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 18001
transform 1 0 51152 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_505
timestamp 1636986456
transform 1 0 51336 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_517
timestamp 1636986456
transform 1 0 52440 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_529
timestamp 1636986456
transform 1 0 53544 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_541
timestamp 1636986456
transform 1 0 54648 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_553
timestamp 18001
transform 1 0 55752 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_559
timestamp 18001
transform 1 0 56304 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_561
timestamp 1636986456
transform 1 0 56488 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_573
timestamp 1636986456
transform 1 0 57592 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_585
timestamp 1636986456
transform 1 0 58696 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_597
timestamp 1636986456
transform 1 0 59800 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_609
timestamp 18001
transform 1 0 60904 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_615
timestamp 18001
transform 1 0 61456 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_617
timestamp 1636986456
transform 1 0 61640 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_629
timestamp 1636986456
transform 1 0 62744 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_641
timestamp 1636986456
transform 1 0 63848 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_653
timestamp 1636986456
transform 1 0 64952 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_665
timestamp 18001
transform 1 0 66056 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_671
timestamp 18001
transform 1 0 66608 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_673
timestamp 1636986456
transform 1 0 66792 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_685
timestamp 1636986456
transform 1 0 67896 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_697
timestamp 1636986456
transform 1 0 69000 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_709
timestamp 1636986456
transform 1 0 70104 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_721
timestamp 18001
transform 1 0 71208 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_727
timestamp 18001
transform 1 0 71760 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_729
timestamp 1636986456
transform 1 0 71944 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_741
timestamp 1636986456
transform 1 0 73048 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_753
timestamp 1636986456
transform 1 0 74152 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_765
timestamp 1636986456
transform 1 0 75256 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_777
timestamp 18001
transform 1 0 76360 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_783
timestamp 18001
transform 1 0 76912 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_785
timestamp 1636986456
transform 1 0 77096 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_797
timestamp 1636986456
transform 1 0 78200 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_809
timestamp 1636986456
transform 1 0 79304 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_821
timestamp 1636986456
transform 1 0 80408 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_833
timestamp 18001
transform 1 0 81512 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_839
timestamp 18001
transform 1 0 82064 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_851
timestamp 1636986456
transform 1 0 83168 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_863
timestamp 1636986456
transform 1 0 84272 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_875
timestamp 1636986456
transform 1 0 85376 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_887
timestamp 18001
transform 1 0 86480 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_895
timestamp 18001
transform 1 0 87216 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_897
timestamp 1636986456
transform 1 0 87400 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_909
timestamp 18001
transform 1 0 88504 0 -1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1636986456
transform 1 0 5152 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1636986456
transform 1 0 6256 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 18001
transform 1 0 7360 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1636986456
transform 1 0 7544 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1636986456
transform 1 0 8648 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1636986456
transform 1 0 9752 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1636986456
transform 1 0 10856 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 18001
transform 1 0 11960 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 18001
transform 1 0 12512 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1636986456
transform 1 0 12696 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1636986456
transform 1 0 13800 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1636986456
transform 1 0 14904 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1636986456
transform 1 0 16008 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 18001
transform 1 0 17112 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 18001
transform 1 0 17664 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1636986456
transform 1 0 17848 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1636986456
transform 1 0 18952 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1636986456
transform 1 0 20056 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1636986456
transform 1 0 21160 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 18001
transform 1 0 22264 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 18001
transform 1 0 22816 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1636986456
transform 1 0 23000 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1636986456
transform 1 0 24104 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1636986456
transform 1 0 25208 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1636986456
transform 1 0 26312 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 18001
transform 1 0 27416 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 18001
transform 1 0 27968 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1636986456
transform 1 0 28152 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1636986456
transform 1 0 29256 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1636986456
transform 1 0 30360 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1636986456
transform 1 0 31464 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 18001
transform 1 0 32568 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 18001
transform 1 0 33120 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1636986456
transform 1 0 33304 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1636986456
transform 1 0 34408 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1636986456
transform 1 0 35512 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1636986456
transform 1 0 36616 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 18001
transform 1 0 37720 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 18001
transform 1 0 38272 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1636986456
transform 1 0 38456 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1636986456
transform 1 0 39560 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1636986456
transform 1 0 40664 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_401
timestamp 1636986456
transform 1 0 41768 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 18001
transform 1 0 42872 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 18001
transform 1 0 43424 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 1636986456
transform 1 0 43608 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 1636986456
transform 1 0 44712 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_445
timestamp 1636986456
transform 1 0 45816 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_457
timestamp 1636986456
transform 1 0 46920 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_469
timestamp 18001
transform 1 0 48024 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 18001
transform 1 0 48576 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_477
timestamp 1636986456
transform 1 0 48760 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_489
timestamp 1636986456
transform 1 0 49864 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_501
timestamp 1636986456
transform 1 0 50968 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_513
timestamp 1636986456
transform 1 0 52072 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_525
timestamp 18001
transform 1 0 53176 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_531
timestamp 18001
transform 1 0 53728 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_533
timestamp 1636986456
transform 1 0 53912 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_545
timestamp 1636986456
transform 1 0 55016 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_557
timestamp 1636986456
transform 1 0 56120 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_569
timestamp 1636986456
transform 1 0 57224 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_581
timestamp 18001
transform 1 0 58328 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_587
timestamp 18001
transform 1 0 58880 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_589
timestamp 1636986456
transform 1 0 59064 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_601
timestamp 1636986456
transform 1 0 60168 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_613
timestamp 1636986456
transform 1 0 61272 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_625
timestamp 1636986456
transform 1 0 62376 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_637
timestamp 18001
transform 1 0 63480 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_643
timestamp 18001
transform 1 0 64032 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_645
timestamp 1636986456
transform 1 0 64216 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_657
timestamp 1636986456
transform 1 0 65320 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_669
timestamp 1636986456
transform 1 0 66424 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_681
timestamp 1636986456
transform 1 0 67528 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_693
timestamp 18001
transform 1 0 68632 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_699
timestamp 18001
transform 1 0 69184 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_701
timestamp 1636986456
transform 1 0 69368 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_713
timestamp 1636986456
transform 1 0 70472 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_725
timestamp 1636986456
transform 1 0 71576 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_737
timestamp 1636986456
transform 1 0 72680 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_749
timestamp 18001
transform 1 0 73784 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_755
timestamp 18001
transform 1 0 74336 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_757
timestamp 1636986456
transform 1 0 74520 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_769
timestamp 1636986456
transform 1 0 75624 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_781
timestamp 1636986456
transform 1 0 76728 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_793
timestamp 1636986456
transform 1 0 77832 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_805
timestamp 18001
transform 1 0 78936 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_811
timestamp 18001
transform 1 0 79488 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_813
timestamp 1636986456
transform 1 0 79672 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_825
timestamp 1636986456
transform 1 0 80776 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_837
timestamp 1636986456
transform 1 0 81880 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_849
timestamp 1636986456
transform 1 0 82984 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_861
timestamp 18001
transform 1 0 84088 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_867
timestamp 18001
transform 1 0 84640 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_869
timestamp 1636986456
transform 1 0 84824 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_881
timestamp 1636986456
transform 1 0 85928 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_893
timestamp 1636986456
transform 1 0 87032 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_905
timestamp 18001
transform 1 0 88136 0 1 5984
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1636986456
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1636986456
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1636986456
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1636986456
transform 1 0 8464 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 18001
transform 1 0 9568 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 18001
transform 1 0 9936 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1636986456
transform 1 0 10120 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1636986456
transform 1 0 11224 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1636986456
transform 1 0 12328 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1636986456
transform 1 0 13432 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 18001
transform 1 0 14536 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 18001
transform 1 0 15088 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1636986456
transform 1 0 15272 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1636986456
transform 1 0 16376 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1636986456
transform 1 0 17480 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1636986456
transform 1 0 18584 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 18001
transform 1 0 19688 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 18001
transform 1 0 20240 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1636986456
transform 1 0 20424 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1636986456
transform 1 0 21528 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1636986456
transform 1 0 22632 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1636986456
transform 1 0 23736 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 18001
transform 1 0 24840 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 18001
transform 1 0 25392 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1636986456
transform 1 0 25576 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1636986456
transform 1 0 26680 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1636986456
transform 1 0 27784 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1636986456
transform 1 0 28888 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 18001
transform 1 0 29992 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 18001
transform 1 0 30544 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1636986456
transform 1 0 30728 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1636986456
transform 1 0 31832 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1636986456
transform 1 0 32936 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1636986456
transform 1 0 34040 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 18001
transform 1 0 35144 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 18001
transform 1 0 35696 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1636986456
transform 1 0 35880 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1636986456
transform 1 0 36984 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1636986456
transform 1 0 38088 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1636986456
transform 1 0 39192 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 18001
transform 1 0 40296 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 18001
transform 1 0 40848 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1636986456
transform 1 0 41032 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1636986456
transform 1 0 42136 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1636986456
transform 1 0 43240 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1636986456
transform 1 0 44344 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 18001
transform 1 0 45448 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 18001
transform 1 0 46000 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1636986456
transform 1 0 46184 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1636986456
transform 1 0 47288 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1636986456
transform 1 0 48392 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_485
timestamp 1636986456
transform 1 0 49496 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 18001
transform 1 0 50600 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 18001
transform 1 0 51152 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_505
timestamp 1636986456
transform 1 0 51336 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_517
timestamp 1636986456
transform 1 0 52440 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_529
timestamp 1636986456
transform 1 0 53544 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_541
timestamp 1636986456
transform 1 0 54648 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_553
timestamp 18001
transform 1 0 55752 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_559
timestamp 18001
transform 1 0 56304 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_561
timestamp 1636986456
transform 1 0 56488 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_573
timestamp 1636986456
transform 1 0 57592 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_585
timestamp 1636986456
transform 1 0 58696 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_597
timestamp 1636986456
transform 1 0 59800 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_609
timestamp 18001
transform 1 0 60904 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_615
timestamp 18001
transform 1 0 61456 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_617
timestamp 1636986456
transform 1 0 61640 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_629
timestamp 1636986456
transform 1 0 62744 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_641
timestamp 1636986456
transform 1 0 63848 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_653
timestamp 1636986456
transform 1 0 64952 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_665
timestamp 18001
transform 1 0 66056 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_671
timestamp 18001
transform 1 0 66608 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_673
timestamp 1636986456
transform 1 0 66792 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_685
timestamp 1636986456
transform 1 0 67896 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_697
timestamp 1636986456
transform 1 0 69000 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_709
timestamp 1636986456
transform 1 0 70104 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_721
timestamp 18001
transform 1 0 71208 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_727
timestamp 18001
transform 1 0 71760 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_729
timestamp 1636986456
transform 1 0 71944 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_741
timestamp 1636986456
transform 1 0 73048 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_753
timestamp 1636986456
transform 1 0 74152 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_765
timestamp 1636986456
transform 1 0 75256 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_777
timestamp 18001
transform 1 0 76360 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_783
timestamp 18001
transform 1 0 76912 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_785
timestamp 1636986456
transform 1 0 77096 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_797
timestamp 1636986456
transform 1 0 78200 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_809
timestamp 1636986456
transform 1 0 79304 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_821
timestamp 1636986456
transform 1 0 80408 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_833
timestamp 18001
transform 1 0 81512 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_839
timestamp 18001
transform 1 0 82064 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_841
timestamp 1636986456
transform 1 0 82248 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_853
timestamp 1636986456
transform 1 0 83352 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_865
timestamp 1636986456
transform 1 0 84456 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_877
timestamp 1636986456
transform 1 0 85560 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_889
timestamp 18001
transform 1 0 86664 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_895
timestamp 18001
transform 1 0 87216 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_897
timestamp 1636986456
transform 1 0 87400 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_909
timestamp 18001
transform 1 0 88504 0 -1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1636986456
transform 1 0 5152 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1636986456
transform 1 0 6256 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 18001
transform 1 0 7360 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1636986456
transform 1 0 7544 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1636986456
transform 1 0 8648 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_53
timestamp 18001
transform 1 0 9752 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_57
timestamp 1636986456
transform 1 0 10120 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_69
timestamp 1636986456
transform 1 0 11224 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_81
timestamp 18001
transform 1 0 12328 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1636986456
transform 1 0 12696 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1636986456
transform 1 0 13800 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_109
timestamp 18001
transform 1 0 14904 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_113
timestamp 1636986456
transform 1 0 15272 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_125
timestamp 1636986456
transform 1 0 16376 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_137
timestamp 18001
transform 1 0 17480 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1636986456
transform 1 0 17848 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1636986456
transform 1 0 18952 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_165
timestamp 18001
transform 1 0 20056 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_169
timestamp 1636986456
transform 1 0 20424 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_181
timestamp 1636986456
transform 1 0 21528 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_193
timestamp 18001
transform 1 0 22632 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1636986456
transform 1 0 23000 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1636986456
transform 1 0 24104 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_221
timestamp 18001
transform 1 0 25208 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_225
timestamp 1636986456
transform 1 0 25576 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_237
timestamp 1636986456
transform 1 0 26680 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_249
timestamp 18001
transform 1 0 27784 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1636986456
transform 1 0 28152 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1636986456
transform 1 0 29256 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_277
timestamp 18001
transform 1 0 30360 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_281
timestamp 1636986456
transform 1 0 30728 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_293
timestamp 1636986456
transform 1 0 31832 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_305
timestamp 18001
transform 1 0 32936 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1636986456
transform 1 0 33304 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1636986456
transform 1 0 34408 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_333
timestamp 18001
transform 1 0 35512 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_337
timestamp 1636986456
transform 1 0 35880 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_349
timestamp 1636986456
transform 1 0 36984 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_361
timestamp 18001
transform 1 0 38088 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1636986456
transform 1 0 38456 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1636986456
transform 1 0 39560 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_389
timestamp 18001
transform 1 0 40664 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_393
timestamp 1636986456
transform 1 0 41032 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_405
timestamp 1636986456
transform 1 0 42136 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_417
timestamp 18001
transform 1 0 43240 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1636986456
transform 1 0 43608 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1636986456
transform 1 0 44712 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_445
timestamp 18001
transform 1 0 45816 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_449
timestamp 1636986456
transform 1 0 46184 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_461
timestamp 1636986456
transform 1 0 47288 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_473
timestamp 18001
transform 1 0 48392 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1636986456
transform 1 0 48760 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1636986456
transform 1 0 49864 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_501
timestamp 18001
transform 1 0 50968 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_505
timestamp 1636986456
transform 1 0 51336 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_517
timestamp 1636986456
transform 1 0 52440 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_529
timestamp 18001
transform 1 0 53544 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_533
timestamp 1636986456
transform 1 0 53912 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_545
timestamp 1636986456
transform 1 0 55016 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_557
timestamp 18001
transform 1 0 56120 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_561
timestamp 1636986456
transform 1 0 56488 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_573
timestamp 1636986456
transform 1 0 57592 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_585
timestamp 18001
transform 1 0 58696 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_589
timestamp 1636986456
transform 1 0 59064 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_601
timestamp 1636986456
transform 1 0 60168 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_613
timestamp 18001
transform 1 0 61272 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_617
timestamp 1636986456
transform 1 0 61640 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_629
timestamp 1636986456
transform 1 0 62744 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_641
timestamp 18001
transform 1 0 63848 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_645
timestamp 1636986456
transform 1 0 64216 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_657
timestamp 1636986456
transform 1 0 65320 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_669
timestamp 18001
transform 1 0 66424 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_673
timestamp 1636986456
transform 1 0 66792 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_685
timestamp 1636986456
transform 1 0 67896 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_697
timestamp 18001
transform 1 0 69000 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_701
timestamp 1636986456
transform 1 0 69368 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_713
timestamp 1636986456
transform 1 0 70472 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_725
timestamp 18001
transform 1 0 71576 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_729
timestamp 1636986456
transform 1 0 71944 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_741
timestamp 1636986456
transform 1 0 73048 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_753
timestamp 18001
transform 1 0 74152 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_757
timestamp 1636986456
transform 1 0 74520 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_769
timestamp 1636986456
transform 1 0 75624 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_781
timestamp 18001
transform 1 0 76728 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_785
timestamp 1636986456
transform 1 0 77096 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_797
timestamp 1636986456
transform 1 0 78200 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_809
timestamp 18001
transform 1 0 79304 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_813
timestamp 1636986456
transform 1 0 79672 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_825
timestamp 1636986456
transform 1 0 80776 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_837
timestamp 18001
transform 1 0 81880 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_841
timestamp 1636986456
transform 1 0 82248 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_853
timestamp 1636986456
transform 1 0 83352 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_865
timestamp 18001
transform 1 0 84456 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_869
timestamp 1636986456
transform 1 0 84824 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_881
timestamp 1636986456
transform 1 0 85928 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_893
timestamp 18001
transform 1 0 87032 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_897
timestamp 1636986456
transform 1 0 87400 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_909
timestamp 18001
transform 1 0 88504 0 1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1636986456
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1636986456
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_27
timestamp 18001
transform 1 0 7360 0 -1 8160
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_885
timestamp 1636986456
transform 1 0 86296 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_897
timestamp 1636986456
transform 1 0 87400 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_909
timestamp 18001
transform 1 0 88504 0 -1 8160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1636986456
transform 1 0 5152 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1636986456
transform 1 0 6256 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 18001
transform 1 0 7360 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_29
timestamp 18001
transform 1 0 7544 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_885
timestamp 1636986456
transform 1 0 86296 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_897
timestamp 1636986456
transform 1 0 87400 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_909
timestamp 18001
transform 1 0 88504 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1636986456
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1636986456
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_27
timestamp 18001
transform 1 0 7360 0 -1 9248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_885
timestamp 1636986456
transform 1 0 86296 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_897
timestamp 1636986456
transform 1 0 87400 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_909
timestamp 18001
transform 1 0 88504 0 -1 9248
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1636986456
transform 1 0 5152 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1636986456
transform 1 0 6256 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 18001
transform 1 0 7360 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_29
timestamp 18001
transform 1 0 7544 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_885
timestamp 1636986456
transform 1 0 86296 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_897
timestamp 1636986456
transform 1 0 87400 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_909
timestamp 18001
transform 1 0 88504 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1636986456
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1636986456
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_27
timestamp 18001
transform 1 0 7360 0 -1 10336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_885
timestamp 1636986456
transform 1 0 86296 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_897
timestamp 1636986456
transform 1 0 87400 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_909
timestamp 18001
transform 1 0 88504 0 -1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1636986456
transform 1 0 5152 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1636986456
transform 1 0 6256 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 18001
transform 1 0 7360 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_29
timestamp 18001
transform 1 0 7544 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_885
timestamp 1636986456
transform 1 0 86296 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_897
timestamp 1636986456
transform 1 0 87400 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_909
timestamp 18001
transform 1 0 88504 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1636986456
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1636986456
transform 1 0 6256 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_27
timestamp 18001
transform 1 0 7360 0 -1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_885
timestamp 1636986456
transform 1 0 86296 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_897
timestamp 1636986456
transform 1 0 87400 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_909
timestamp 18001
transform 1 0 88504 0 -1 11424
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1636986456
transform 1 0 5152 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1636986456
transform 1 0 6256 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 18001
transform 1 0 7360 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_29
timestamp 18001
transform 1 0 7544 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_885
timestamp 1636986456
transform 1 0 86296 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_897
timestamp 1636986456
transform 1 0 87400 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_909
timestamp 18001
transform 1 0 88504 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1636986456
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1636986456
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_27
timestamp 18001
transform 1 0 7360 0 -1 12512
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_885
timestamp 1636986456
transform 1 0 86296 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_897
timestamp 1636986456
transform 1 0 87400 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_909
timestamp 18001
transform 1 0 88504 0 -1 12512
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1636986456
transform 1 0 5152 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1636986456
transform 1 0 6256 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 18001
transform 1 0 7360 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_29
timestamp 18001
transform 1 0 7544 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_885
timestamp 1636986456
transform 1 0 86296 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_897
timestamp 1636986456
transform 1 0 87400 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_909
timestamp 18001
transform 1 0 88504 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1636986456
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1636986456
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_27
timestamp 18001
transform 1 0 7360 0 -1 13600
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_885
timestamp 1636986456
transform 1 0 86296 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_897
timestamp 1636986456
transform 1 0 87400 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_909
timestamp 18001
transform 1 0 88504 0 -1 13600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1636986456
transform 1 0 5152 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1636986456
transform 1 0 6256 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 18001
transform 1 0 7360 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_29
timestamp 18001
transform 1 0 7544 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_885
timestamp 1636986456
transform 1 0 86296 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_897
timestamp 1636986456
transform 1 0 87400 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_909
timestamp 18001
transform 1 0 88504 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_6
timestamp 1636986456
transform 1 0 5428 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_18
timestamp 1636986456
transform 1 0 6532 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_885
timestamp 1636986456
transform 1 0 86296 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_897
timestamp 18001
transform 1 0 87400 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_905
timestamp 18001
transform 1 0 88136 0 -1 14688
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_6
timestamp 1636986456
transform 1 0 5428 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_18
timestamp 18001
transform 1 0 6532 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_26
timestamp 18001
transform 1 0 7268 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_29
timestamp 18001
transform 1 0 7544 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_885
timestamp 1636986456
transform 1 0 86296 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_897
timestamp 18001
transform 1 0 87400 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_905
timestamp 18001
transform 1 0 88136 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1636986456
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1636986456
transform 1 0 6256 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_27
timestamp 18001
transform 1 0 7360 0 -1 15776
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_885
timestamp 1636986456
transform 1 0 86296 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_897
timestamp 1636986456
transform 1 0 87400 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_909
timestamp 18001
transform 1 0 88504 0 -1 15776
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_6
timestamp 1636986456
transform 1 0 5428 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_18
timestamp 18001
transform 1 0 6532 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 18001
transform 1 0 7268 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_29
timestamp 18001
transform 1 0 7544 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_885
timestamp 1636986456
transform 1 0 86296 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_897
timestamp 18001
transform 1 0 87400 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_905
timestamp 18001
transform 1 0 88136 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1636986456
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1636986456
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_27
timestamp 18001
transform 1 0 7360 0 -1 16864
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_885
timestamp 1636986456
transform 1 0 86296 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_897
timestamp 1636986456
transform 1 0 87400 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_909
timestamp 18001
transform 1 0 88504 0 -1 16864
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_6
timestamp 1636986456
transform 1 0 5428 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_18
timestamp 18001
transform 1 0 6532 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 18001
transform 1 0 7268 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_29
timestamp 18001
transform 1 0 7544 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_885
timestamp 1636986456
transform 1 0 86296 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_897
timestamp 18001
transform 1 0 87400 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_905
timestamp 18001
transform 1 0 88136 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1636986456
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1636986456
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_27
timestamp 18001
transform 1 0 7360 0 -1 17952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_885
timestamp 1636986456
transform 1 0 86296 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_897
timestamp 1636986456
transform 1 0 87400 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_909
timestamp 18001
transform 1 0 88504 0 -1 17952
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_6
timestamp 1636986456
transform 1 0 5428 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_18
timestamp 18001
transform 1 0 6532 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_26
timestamp 18001
transform 1 0 7268 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_29
timestamp 18001
transform 1 0 7544 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_885
timestamp 1636986456
transform 1 0 86296 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_897
timestamp 18001
transform 1 0 87400 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_905
timestamp 18001
transform 1 0 88136 0 1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1636986456
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1636986456
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_27
timestamp 18001
transform 1 0 7360 0 -1 19040
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_885
timestamp 1636986456
transform 1 0 86296 0 -1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_897
timestamp 1636986456
transform 1 0 87400 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_909
timestamp 18001
transform 1 0 88504 0 -1 19040
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1636986456
transform 1 0 5152 0 1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1636986456
transform 1 0 6256 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 18001
transform 1 0 7360 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_29
timestamp 18001
transform 1 0 7544 0 1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_885
timestamp 1636986456
transform 1 0 86296 0 1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_897
timestamp 1636986456
transform 1 0 87400 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_909
timestamp 18001
transform 1 0 88504 0 1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_6
timestamp 1636986456
transform 1 0 5428 0 -1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_18
timestamp 1636986456
transform 1 0 6532 0 -1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_885
timestamp 1636986456
transform 1 0 86296 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_897
timestamp 18001
transform 1 0 87400 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_905
timestamp 18001
transform 1 0 88136 0 -1 20128
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_6
timestamp 1636986456
transform 1 0 5428 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_18
timestamp 18001
transform 1 0 6532 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_26
timestamp 18001
transform 1 0 7268 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_29
timestamp 18001
transform 1 0 7544 0 1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_885
timestamp 1636986456
transform 1 0 86296 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_897
timestamp 18001
transform 1 0 87400 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_905
timestamp 18001
transform 1 0 88136 0 1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1636986456
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1636986456
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_27
timestamp 18001
transform 1 0 7360 0 -1 21216
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_885
timestamp 1636986456
transform 1 0 86296 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_897
timestamp 1636986456
transform 1 0 87400 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_909
timestamp 18001
transform 1 0 88504 0 -1 21216
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_6
timestamp 1636986456
transform 1 0 5428 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_18
timestamp 18001
transform 1 0 6532 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_26
timestamp 18001
transform 1 0 7268 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_29
timestamp 18001
transform 1 0 7544 0 1 21216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_885
timestamp 1636986456
transform 1 0 86296 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_897
timestamp 18001
transform 1 0 87400 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_905
timestamp 18001
transform 1 0 88136 0 1 21216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1636986456
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1636986456
transform 1 0 6256 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_27
timestamp 18001
transform 1 0 7360 0 -1 22304
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_885
timestamp 1636986456
transform 1 0 86296 0 -1 22304
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_897
timestamp 1636986456
transform 1 0 87400 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_909
timestamp 18001
transform 1 0 88504 0 -1 22304
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_6
timestamp 1636986456
transform 1 0 5428 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_18
timestamp 18001
transform 1 0 6532 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_26
timestamp 18001
transform 1 0 7268 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_29
timestamp 18001
transform 1 0 7544 0 1 22304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_885
timestamp 1636986456
transform 1 0 86296 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_897
timestamp 18001
transform 1 0 87400 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_905
timestamp 18001
transform 1 0 88136 0 1 22304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1636986456
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1636986456
transform 1 0 6256 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_27
timestamp 18001
transform 1 0 7360 0 -1 23392
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_885
timestamp 1636986456
transform 1 0 86296 0 -1 23392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_897
timestamp 1636986456
transform 1 0 87400 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_909
timestamp 18001
transform 1 0 88504 0 -1 23392
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_6
timestamp 1636986456
transform 1 0 5428 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_18
timestamp 18001
transform 1 0 6532 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_26
timestamp 18001
transform 1 0 7268 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_29
timestamp 18001
transform 1 0 7544 0 1 23392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_885
timestamp 1636986456
transform 1 0 86296 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_897
timestamp 18001
transform 1 0 87400 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_905
timestamp 18001
transform 1 0 88136 0 1 23392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1636986456
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1636986456
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_27
timestamp 18001
transform 1 0 7360 0 -1 24480
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_885
timestamp 1636986456
transform 1 0 86296 0 -1 24480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_897
timestamp 1636986456
transform 1 0 87400 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_909
timestamp 18001
transform 1 0 88504 0 -1 24480
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1636986456
transform 1 0 5152 0 1 24480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1636986456
transform 1 0 6256 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 18001
transform 1 0 7360 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_29
timestamp 18001
transform 1 0 7544 0 1 24480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_885
timestamp 1636986456
transform 1 0 86296 0 1 24480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_897
timestamp 1636986456
transform 1 0 87400 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_909
timestamp 18001
transform 1 0 88504 0 1 24480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_6
timestamp 1636986456
transform 1 0 5428 0 -1 25568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_18
timestamp 1636986456
transform 1 0 6532 0 -1 25568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_885
timestamp 1636986456
transform 1 0 86296 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_897
timestamp 18001
transform 1 0 87400 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_905
timestamp 18001
transform 1 0 88136 0 -1 25568
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_6
timestamp 1636986456
transform 1 0 5428 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_18
timestamp 18001
transform 1 0 6532 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_26
timestamp 18001
transform 1 0 7268 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_29
timestamp 18001
transform 1 0 7544 0 1 25568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_885
timestamp 1636986456
transform 1 0 86296 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_897
timestamp 18001
transform 1 0 87400 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_905
timestamp 18001
transform 1 0 88136 0 1 25568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1636986456
transform 1 0 5152 0 -1 26656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1636986456
transform 1 0 6256 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_27
timestamp 18001
transform 1 0 7360 0 -1 26656
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_885
timestamp 1636986456
transform 1 0 86296 0 -1 26656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_897
timestamp 1636986456
transform 1 0 87400 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_909
timestamp 18001
transform 1 0 88504 0 -1 26656
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_6
timestamp 1636986456
transform 1 0 5428 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_18
timestamp 18001
transform 1 0 6532 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_26
timestamp 18001
transform 1 0 7268 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_29
timestamp 18001
transform 1 0 7544 0 1 26656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_885
timestamp 1636986456
transform 1 0 86296 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_897
timestamp 18001
transform 1 0 87400 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_905
timestamp 18001
transform 1 0 88136 0 1 26656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1636986456
transform 1 0 5152 0 -1 27744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1636986456
transform 1 0 6256 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_27
timestamp 18001
transform 1 0 7360 0 -1 27744
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_885
timestamp 1636986456
transform 1 0 86296 0 -1 27744
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_897
timestamp 1636986456
transform 1 0 87400 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_909
timestamp 18001
transform 1 0 88504 0 -1 27744
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_6
timestamp 1636986456
transform 1 0 5428 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_18
timestamp 18001
transform 1 0 6532 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_26
timestamp 18001
transform 1 0 7268 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_29
timestamp 18001
transform 1 0 7544 0 1 27744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_885
timestamp 1636986456
transform 1 0 86296 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_897
timestamp 18001
transform 1 0 87400 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_905
timestamp 18001
transform 1 0 88136 0 1 27744
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1636986456
transform 1 0 5152 0 -1 28832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1636986456
transform 1 0 6256 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_27
timestamp 18001
transform 1 0 7360 0 -1 28832
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_885
timestamp 1636986456
transform 1 0 86296 0 -1 28832
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_897
timestamp 1636986456
transform 1 0 87400 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_909
timestamp 18001
transform 1 0 88504 0 -1 28832
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_7
timestamp 1636986456
transform 1 0 5520 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_19
timestamp 18001
transform 1 0 6624 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 18001
transform 1 0 7360 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_44_29
timestamp 18001
transform 1 0 7544 0 1 28832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_885
timestamp 1636986456
transform 1 0 86296 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_897
timestamp 18001
transform 1 0 87400 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_905
timestamp 18001
transform 1 0 88136 0 1 28832
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1636986456
transform 1 0 5152 0 -1 29920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1636986456
transform 1 0 6256 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_27
timestamp 18001
transform 1 0 7360 0 -1 29920
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_885
timestamp 1636986456
transform 1 0 86296 0 -1 29920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_897
timestamp 1636986456
transform 1 0 87400 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_909
timestamp 18001
transform 1 0 88504 0 -1 29920
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1636986456
transform 1 0 5152 0 1 29920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1636986456
transform 1 0 6256 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 18001
transform 1 0 7360 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_46_29
timestamp 18001
transform 1 0 7544 0 1 29920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_885
timestamp 1636986456
transform 1 0 86296 0 1 29920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_897
timestamp 1636986456
transform 1 0 87400 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_909
timestamp 18001
transform 1 0 88504 0 1 29920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_7
timestamp 1636986456
transform 1 0 5520 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_19
timestamp 18001
transform 1 0 6624 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_27
timestamp 18001
transform 1 0 7360 0 -1 31008
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_885
timestamp 1636986456
transform 1 0 86296 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_897
timestamp 18001
transform 1 0 87400 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_905
timestamp 18001
transform 1 0 88136 0 -1 31008
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_7
timestamp 1636986456
transform 1 0 5520 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_19
timestamp 18001
transform 1 0 6624 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 18001
transform 1 0 7360 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_48_29
timestamp 18001
transform 1 0 7544 0 1 31008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_885
timestamp 1636986456
transform 1 0 86296 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_897
timestamp 18001
transform 1 0 87400 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_905
timestamp 18001
transform 1 0 88136 0 1 31008
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1636986456
transform 1 0 5152 0 -1 32096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1636986456
transform 1 0 6256 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_27
timestamp 18001
transform 1 0 7360 0 -1 32096
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_885
timestamp 1636986456
transform 1 0 86296 0 -1 32096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_897
timestamp 1636986456
transform 1 0 87400 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_909
timestamp 18001
transform 1 0 88504 0 -1 32096
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_7
timestamp 1636986456
transform 1 0 5520 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_19
timestamp 18001
transform 1 0 6624 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 18001
transform 1 0 7360 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_50_29
timestamp 18001
transform 1 0 7544 0 1 32096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_885
timestamp 1636986456
transform 1 0 86296 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_897
timestamp 18001
transform 1 0 87400 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_905
timestamp 18001
transform 1 0 88136 0 1 32096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1636986456
transform 1 0 5152 0 -1 33184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1636986456
transform 1 0 6256 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_27
timestamp 18001
transform 1 0 7360 0 -1 33184
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_885
timestamp 1636986456
transform 1 0 86296 0 -1 33184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_897
timestamp 1636986456
transform 1 0 87400 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_909
timestamp 18001
transform 1 0 88504 0 -1 33184
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_7
timestamp 1636986456
transform 1 0 5520 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_19
timestamp 18001
transform 1 0 6624 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 18001
transform 1 0 7360 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_52_29
timestamp 18001
transform 1 0 7544 0 1 33184
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_885
timestamp 1636986456
transform 1 0 86296 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_897
timestamp 18001
transform 1 0 87400 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_905
timestamp 18001
transform 1 0 88136 0 1 33184
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_6
timestamp 1636986456
transform 1 0 5428 0 -1 34272
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_18
timestamp 1636986456
transform 1 0 6532 0 -1 34272
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_885
timestamp 1636986456
transform 1 0 86296 0 -1 34272
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_897
timestamp 1636986456
transform 1 0 87400 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_909
timestamp 18001
transform 1 0 88504 0 -1 34272
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_7
timestamp 1636986456
transform 1 0 5520 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_19
timestamp 18001
transform 1 0 6624 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 18001
transform 1 0 7360 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_54_29
timestamp 18001
transform 1 0 7544 0 1 34272
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_885
timestamp 1636986456
transform 1 0 86296 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_897
timestamp 18001
transform 1 0 87400 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_905
timestamp 18001
transform 1 0 88136 0 1 34272
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1636986456
transform 1 0 5152 0 -1 35360
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1636986456
transform 1 0 6256 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_55_27
timestamp 18001
transform 1 0 7360 0 -1 35360
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_885
timestamp 1636986456
transform 1 0 86296 0 -1 35360
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_897
timestamp 1636986456
transform 1 0 87400 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_909
timestamp 18001
transform 1 0 88504 0 -1 35360
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1636986456
transform 1 0 5152 0 1 35360
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1636986456
transform 1 0 6256 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 18001
transform 1 0 7360 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_56_29
timestamp 18001
transform 1 0 7544 0 1 35360
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_885
timestamp 1636986456
transform 1 0 86296 0 1 35360
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_897
timestamp 1636986456
transform 1 0 87400 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_909
timestamp 18001
transform 1 0 88504 0 1 35360
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_7
timestamp 1636986456
transform 1 0 5520 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_19
timestamp 18001
transform 1 0 6624 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_27
timestamp 18001
transform 1 0 7360 0 -1 36448
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_885
timestamp 1636986456
transform 1 0 86296 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_897
timestamp 18001
transform 1 0 87400 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_905
timestamp 18001
transform 1 0 88136 0 -1 36448
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_58_7
timestamp 1636986456
transform 1 0 5520 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_19
timestamp 18001
transform 1 0 6624 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 18001
transform 1 0 7360 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_58_29
timestamp 18001
transform 1 0 7544 0 1 36448
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_885
timestamp 1636986456
transform 1 0 86296 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_897
timestamp 18001
transform 1 0 87400 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_905
timestamp 18001
transform 1 0 88136 0 1 36448
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1636986456
transform 1 0 5152 0 -1 37536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1636986456
transform 1 0 6256 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_59_27
timestamp 18001
transform 1 0 7360 0 -1 37536
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_885
timestamp 1636986456
transform 1 0 86296 0 -1 37536
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_897
timestamp 1636986456
transform 1 0 87400 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_909
timestamp 18001
transform 1 0 88504 0 -1 37536
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_7
timestamp 1636986456
transform 1 0 5520 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_19
timestamp 18001
transform 1 0 6624 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 18001
transform 1 0 7360 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_60_29
timestamp 18001
transform 1 0 7544 0 1 37536
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_885
timestamp 1636986456
transform 1 0 86296 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_897
timestamp 18001
transform 1 0 87400 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_905
timestamp 18001
transform 1 0 88136 0 1 37536
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1636986456
transform 1 0 5152 0 -1 38624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1636986456
transform 1 0 6256 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_27
timestamp 18001
transform 1 0 7360 0 -1 38624
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_885
timestamp 1636986456
transform 1 0 86296 0 -1 38624
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_897
timestamp 1636986456
transform 1 0 87400 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_909
timestamp 18001
transform 1 0 88504 0 -1 38624
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_7
timestamp 1636986456
transform 1 0 5520 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_19
timestamp 18001
transform 1 0 6624 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 18001
transform 1 0 7360 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_62_29
timestamp 18001
transform 1 0 7544 0 1 38624
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_885
timestamp 1636986456
transform 1 0 86296 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_897
timestamp 18001
transform 1 0 87400 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_905
timestamp 18001
transform 1 0 88136 0 1 38624
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1636986456
transform 1 0 5152 0 -1 39712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1636986456
transform 1 0 6256 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_63_27
timestamp 18001
transform 1 0 7360 0 -1 39712
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_885
timestamp 1636986456
transform 1 0 86296 0 -1 39712
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_897
timestamp 1636986456
transform 1 0 87400 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_909
timestamp 18001
transform 1 0 88504 0 -1 39712
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_7
timestamp 1636986456
transform 1 0 5520 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_19
timestamp 18001
transform 1 0 6624 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 18001
transform 1 0 7360 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_64_29
timestamp 18001
transform 1 0 7544 0 1 39712
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_885
timestamp 1636986456
transform 1 0 86296 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_897
timestamp 18001
transform 1 0 87400 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_903
timestamp 18001
transform 1 0 87952 0 1 39712
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 1636986456
transform 1 0 5152 0 -1 40800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_15
timestamp 1636986456
transform 1 0 6256 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_65_27
timestamp 18001
transform 1 0 7360 0 -1 40800
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_65_885
timestamp 1636986456
transform 1 0 86296 0 -1 40800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_897
timestamp 1636986456
transform 1 0 87400 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_65_909
timestamp 18001
transform 1 0 88504 0 -1 40800
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_3
timestamp 1636986456
transform 1 0 5152 0 1 40800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_15
timestamp 1636986456
transform 1 0 6256 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 18001
transform 1 0 7360 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_66_29
timestamp 18001
transform 1 0 7544 0 1 40800
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_885
timestamp 1636986456
transform 1 0 86296 0 1 40800
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_897
timestamp 1636986456
transform 1 0 87400 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_909
timestamp 18001
transform 1 0 88504 0 1 40800
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_7
timestamp 1636986456
transform 1 0 5520 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_19
timestamp 18001
transform 1 0 6624 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_27
timestamp 18001
transform 1 0 7360 0 -1 41888
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_67_885
timestamp 1636986456
transform 1 0 86296 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_897
timestamp 18001
transform 1 0 87400 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_905
timestamp 18001
transform 1 0 88136 0 -1 41888
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_68_7
timestamp 1636986456
transform 1 0 5520 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_19
timestamp 18001
transform 1 0 6624 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 18001
transform 1 0 7360 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_68_29
timestamp 18001
transform 1 0 7544 0 1 41888
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_885
timestamp 1636986456
transform 1 0 86296 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_897
timestamp 18001
transform 1 0 87400 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_905
timestamp 18001
transform 1 0 88136 0 1 41888
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_6
timestamp 1636986456
transform 1 0 5428 0 -1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_18
timestamp 1636986456
transform 1 0 6532 0 -1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_885
timestamp 1636986456
transform 1 0 86296 0 -1 42976
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_897
timestamp 1636986456
transform 1 0 87400 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_69_909
timestamp 18001
transform 1 0 88504 0 -1 42976
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_7
timestamp 1636986456
transform 1 0 5520 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_19
timestamp 18001
transform 1 0 6624 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 18001
transform 1 0 7360 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_70_29
timestamp 18001
transform 1 0 7544 0 1 42976
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_885
timestamp 1636986456
transform 1 0 86296 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_70_897
timestamp 18001
transform 1 0 87400 0 1 42976
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_71_3
timestamp 1636986456
transform 1 0 5152 0 -1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 1636986456
transform 1 0 6256 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_71_27
timestamp 18001
transform 1 0 7360 0 -1 44064
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_71_885
timestamp 1636986456
transform 1 0 86296 0 -1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_897
timestamp 1636986456
transform 1 0 87400 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_909
timestamp 18001
transform 1 0 88504 0 -1 44064
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_6
timestamp 1636986456
transform 1 0 5428 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_18
timestamp 18001
transform 1 0 6532 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_26
timestamp 18001
transform 1 0 7268 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_72_29
timestamp 18001
transform 1 0 7544 0 1 44064
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_885
timestamp 1636986456
transform 1 0 86296 0 1 44064
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_897
timestamp 1636986456
transform 1 0 87400 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_909
timestamp 18001
transform 1 0 88504 0 1 44064
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_6
timestamp 1636986456
transform 1 0 5428 0 -1 45152
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_18
timestamp 1636986456
transform 1 0 6532 0 -1 45152
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_885
timestamp 1636986456
transform 1 0 86296 0 -1 45152
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_897
timestamp 1636986456
transform 1 0 87400 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_73_909
timestamp 18001
transform 1 0 88504 0 -1 45152
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1636986456
transform 1 0 5152 0 1 45152
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1636986456
transform 1 0 6256 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 18001
transform 1 0 7360 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_74_29
timestamp 18001
transform 1 0 7544 0 1 45152
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_885
timestamp 1636986456
transform 1 0 86296 0 1 45152
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_897
timestamp 1636986456
transform 1 0 87400 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_909
timestamp 18001
transform 1 0 88504 0 1 45152
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_6
timestamp 1636986456
transform 1 0 5428 0 -1 46240
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_18
timestamp 1636986456
transform 1 0 6532 0 -1 46240
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_885
timestamp 1636986456
transform 1 0 86296 0 -1 46240
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_897
timestamp 1636986456
transform 1 0 87400 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_75_909
timestamp 18001
transform 1 0 88504 0 -1 46240
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_3
timestamp 1636986456
transform 1 0 5152 0 1 46240
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_15
timestamp 1636986456
transform 1 0 6256 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 18001
transform 1 0 7360 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_76_29
timestamp 18001
transform 1 0 7544 0 1 46240
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_885
timestamp 1636986456
transform 1 0 86296 0 1 46240
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_897
timestamp 1636986456
transform 1 0 87400 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_909
timestamp 18001
transform 1 0 88504 0 1 46240
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_9
timestamp 1636986456
transform 1 0 5704 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_21
timestamp 18001
transform 1 0 6808 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_77_29
timestamp 18001
transform 1 0 7544 0 -1 47328
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_885
timestamp 1636986456
transform 1 0 86296 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_897
timestamp 18001
transform 1 0 87400 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_77_905
timestamp 18001
transform 1 0 88136 0 -1 47328
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1636986456
transform 1 0 5152 0 1 47328
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1636986456
transform 1 0 6256 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 18001
transform 1 0 7360 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_78_29
timestamp 18001
transform 1 0 7544 0 1 47328
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_885
timestamp 1636986456
transform 1 0 86296 0 1 47328
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_897
timestamp 1636986456
transform 1 0 87400 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_909
timestamp 18001
transform 1 0 88504 0 1 47328
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_3
timestamp 1636986456
transform 1 0 5152 0 -1 48416
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 1636986456
transform 1 0 6256 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_27
timestamp 18001
transform 1 0 7360 0 -1 48416
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_79_885
timestamp 1636986456
transform 1 0 86296 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_897
timestamp 18001
transform 1 0 87400 0 -1 48416
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_80_3
timestamp 1636986456
transform 1 0 5152 0 1 48416
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_15
timestamp 1636986456
transform 1 0 6256 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 18001
transform 1 0 7360 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_80_29
timestamp 18001
transform 1 0 7544 0 1 48416
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_885
timestamp 1636986456
transform 1 0 86296 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_897
timestamp 18001
transform 1 0 87400 0 1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_905
timestamp 18001
transform 1 0 88136 0 1 48416
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_81_3
timestamp 1636986456
transform 1 0 5152 0 -1 49504
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1636986456
transform 1 0 6256 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_81_27
timestamp 18001
transform 1 0 7360 0 -1 49504
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_81_885
timestamp 1636986456
transform 1 0 86296 0 -1 49504
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_897
timestamp 1636986456
transform 1 0 87400 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_81_909
timestamp 18001
transform 1 0 88504 0 -1 49504
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_6
timestamp 1636986456
transform 1 0 5428 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_18
timestamp 18001
transform 1 0 6532 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_26
timestamp 18001
transform 1 0 7268 0 1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_82_29
timestamp 18001
transform 1 0 7544 0 1 49504
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_885
timestamp 1636986456
transform 1 0 86296 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_897
timestamp 18001
transform 1 0 87400 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_905
timestamp 18001
transform 1 0 88136 0 1 49504
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_83_3
timestamp 1636986456
transform 1 0 5152 0 -1 50592
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_15
timestamp 1636986456
transform 1 0 6256 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_83_27
timestamp 18001
transform 1 0 7360 0 -1 50592
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_83_885
timestamp 1636986456
transform 1 0 86296 0 -1 50592
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_897
timestamp 1636986456
transform 1 0 87400 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_83_909
timestamp 18001
transform 1 0 88504 0 -1 50592
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_84_3
timestamp 1636986456
transform 1 0 5152 0 1 50592
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_15
timestamp 1636986456
transform 1 0 6256 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 18001
transform 1 0 7360 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_84_29
timestamp 18001
transform 1 0 7544 0 1 50592
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_885
timestamp 1636986456
transform 1 0 86296 0 1 50592
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_897
timestamp 1636986456
transform 1 0 87400 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_909
timestamp 18001
transform 1 0 88504 0 1 50592
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_6
timestamp 1636986456
transform 1 0 5428 0 -1 51680
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_18
timestamp 1636986456
transform 1 0 6532 0 -1 51680
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_885
timestamp 1636986456
transform 1 0 86296 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_897
timestamp 18001
transform 1 0 87400 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_85_905
timestamp 18001
transform 1 0 88136 0 -1 51680
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_86_3
timestamp 1636986456
transform 1 0 5152 0 1 51680
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_15
timestamp 1636986456
transform 1 0 6256 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 18001
transform 1 0 7360 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_86_29
timestamp 18001
transform 1 0 7544 0 1 51680
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_885
timestamp 1636986456
transform 1 0 86296 0 1 51680
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_897
timestamp 1636986456
transform 1 0 87400 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_909
timestamp 18001
transform 1 0 88504 0 1 51680
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_6
timestamp 1636986456
transform 1 0 5428 0 -1 52768
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_18
timestamp 1636986456
transform 1 0 6532 0 -1 52768
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_885
timestamp 1636986456
transform 1 0 86296 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_897
timestamp 18001
transform 1 0 87400 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_87_905
timestamp 18001
transform 1 0 88136 0 -1 52768
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_88_6
timestamp 1636986456
transform 1 0 5428 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_18
timestamp 18001
transform 1 0 6532 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_88_26
timestamp 18001
transform 1 0 7268 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_88_29
timestamp 18001
transform 1 0 7544 0 1 52768
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_885
timestamp 1636986456
transform 1 0 86296 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_897
timestamp 18001
transform 1 0 87400 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_88_905
timestamp 18001
transform 1 0 88136 0 1 52768
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_89_6
timestamp 1636986456
transform 1 0 5428 0 -1 53856
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_18
timestamp 1636986456
transform 1 0 6532 0 -1 53856
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_885
timestamp 1636986456
transform 1 0 86296 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_89_897
timestamp 18001
transform 1 0 87400 0 -1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_89_905
timestamp 18001
transform 1 0 88136 0 -1 53856
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_90_6
timestamp 1636986456
transform 1 0 5428 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_90_18
timestamp 18001
transform 1 0 6532 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_90_26
timestamp 18001
transform 1 0 7268 0 1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_90_29
timestamp 18001
transform 1 0 7544 0 1 53856
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_885
timestamp 1636986456
transform 1 0 86296 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_90_897
timestamp 18001
transform 1 0 87400 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_90_905
timestamp 18001
transform 1 0 88136 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_91_3
timestamp 18001
transform 1 0 5152 0 -1 54944
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_9
timestamp 18001
transform 1 0 5704 0 -1 54944
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_885
timestamp 1636986456
transform 1 0 86296 0 -1 54944
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_897
timestamp 1636986456
transform 1 0 87400 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_91_909
timestamp 18001
transform 1 0 88504 0 -1 54944
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_92_6
timestamp 1636986456
transform 1 0 5428 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_18
timestamp 18001
transform 1 0 6532 0 1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_92_26
timestamp 18001
transform 1 0 7268 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_92_29
timestamp 18001
transform 1 0 7544 0 1 54944
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_885
timestamp 1636986456
transform 1 0 86296 0 1 54944
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_897
timestamp 1636986456
transform 1 0 87400 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_909
timestamp 18001
transform 1 0 88504 0 1 54944
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_6
timestamp 1636986456
transform 1 0 5428 0 -1 56032
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_18
timestamp 1636986456
transform 1 0 6532 0 -1 56032
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_885
timestamp 1636986456
transform 1 0 86296 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_897
timestamp 18001
transform 1 0 87400 0 -1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_93_905
timestamp 18001
transform 1 0 88136 0 -1 56032
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_94_3
timestamp 1636986456
transform 1 0 5152 0 1 56032
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_15
timestamp 1636986456
transform 1 0 6256 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_27
timestamp 18001
transform 1 0 7360 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_94_29
timestamp 18001
transform 1 0 7544 0 1 56032
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_885
timestamp 1636986456
transform 1 0 86296 0 1 56032
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_897
timestamp 1636986456
transform 1 0 87400 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_909
timestamp 18001
transform 1 0 88504 0 1 56032
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_6
timestamp 1636986456
transform 1 0 5428 0 -1 57120
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_18
timestamp 1636986456
transform 1 0 6532 0 -1 57120
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_885
timestamp 1636986456
transform 1 0 86296 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_95_897
timestamp 18001
transform 1 0 87400 0 -1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_95_905
timestamp 18001
transform 1 0 88136 0 -1 57120
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_96_3
timestamp 1636986456
transform 1 0 5152 0 1 57120
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_15
timestamp 1636986456
transform 1 0 6256 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_96_27
timestamp 18001
transform 1 0 7360 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_96_29
timestamp 18001
transform 1 0 7544 0 1 57120
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_885
timestamp 1636986456
transform 1 0 86296 0 1 57120
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_897
timestamp 1636986456
transform 1 0 87400 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_96_909
timestamp 18001
transform 1 0 88504 0 1 57120
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_6
timestamp 1636986456
transform 1 0 5428 0 -1 58208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_18
timestamp 1636986456
transform 1 0 6532 0 -1 58208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_885
timestamp 1636986456
transform 1 0 86296 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_897
timestamp 18001
transform 1 0 87400 0 -1 58208
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_97_905
timestamp 18001
transform 1 0 88136 0 -1 58208
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_98_3
timestamp 1636986456
transform 1 0 5152 0 1 58208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_15
timestamp 1636986456
transform 1 0 6256 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_27
timestamp 18001
transform 1 0 7360 0 1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_98_29
timestamp 18001
transform 1 0 7544 0 1 58208
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_885
timestamp 1636986456
transform 1 0 86296 0 1 58208
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_897
timestamp 1636986456
transform 1 0 87400 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_909
timestamp 18001
transform 1 0 88504 0 1 58208
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_6
timestamp 1636986456
transform 1 0 5428 0 -1 59296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_18
timestamp 1636986456
transform 1 0 6532 0 -1 59296
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_885
timestamp 1636986456
transform 1 0 86296 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_897
timestamp 18001
transform 1 0 87400 0 -1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_99_905
timestamp 18001
transform 1 0 88136 0 -1 59296
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_100_6
timestamp 1636986456
transform 1 0 5428 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_18
timestamp 18001
transform 1 0 6532 0 1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_100_26
timestamp 18001
transform 1 0 7268 0 1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_100_29
timestamp 18001
transform 1 0 7544 0 1 59296
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_885
timestamp 1636986456
transform 1 0 86296 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_897
timestamp 18001
transform 1 0 87400 0 1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_100_905
timestamp 18001
transform 1 0 88136 0 1 59296
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_3
timestamp 1636986456
transform 1 0 5152 0 -1 60384
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_15
timestamp 1636986456
transform 1 0 6256 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_27
timestamp 18001
transform 1 0 7360 0 -1 60384
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_885
timestamp 1636986456
transform 1 0 86296 0 -1 60384
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_897
timestamp 1636986456
transform 1 0 87400 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_101_909
timestamp 18001
transform 1 0 88504 0 -1 60384
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_102_3
timestamp 1636986456
transform 1 0 5152 0 1 60384
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_15
timestamp 1636986456
transform 1 0 6256 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_102_27
timestamp 18001
transform 1 0 7360 0 1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_102_29
timestamp 18001
transform 1 0 7544 0 1 60384
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_102_885
timestamp 1636986456
transform 1 0 86296 0 1 60384
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_102_897
timestamp 1636986456
transform 1 0 87400 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_102_909
timestamp 18001
transform 1 0 88504 0 1 60384
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_103_6
timestamp 1636986456
transform 1 0 5428 0 -1 61472
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_18
timestamp 1636986456
transform 1 0 6532 0 -1 61472
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_103_885
timestamp 1636986456
transform 1 0 86296 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_103_897
timestamp 18001
transform 1 0 87400 0 -1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_103_905
timestamp 18001
transform 1 0 88136 0 -1 61472
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_104_3
timestamp 1636986456
transform 1 0 5152 0 1 61472
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_15
timestamp 1636986456
transform 1 0 6256 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_104_27
timestamp 18001
transform 1 0 7360 0 1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_104_29
timestamp 18001
transform 1 0 7544 0 1 61472
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_104_885
timestamp 1636986456
transform 1 0 86296 0 1 61472
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_104_897
timestamp 1636986456
transform 1 0 87400 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_104_909
timestamp 18001
transform 1 0 88504 0 1 61472
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_105_6
timestamp 1636986456
transform 1 0 5428 0 -1 62560
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_18
timestamp 1636986456
transform 1 0 6532 0 -1 62560
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_105_885
timestamp 1636986456
transform 1 0 86296 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_105_897
timestamp 18001
transform 1 0 87400 0 -1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_105_905
timestamp 18001
transform 1 0 88136 0 -1 62560
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_106_3
timestamp 1636986456
transform 1 0 5152 0 1 62560
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_15
timestamp 1636986456
transform 1 0 6256 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_106_27
timestamp 18001
transform 1 0 7360 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_106_29
timestamp 18001
transform 1 0 7544 0 1 62560
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_106_885
timestamp 1636986456
transform 1 0 86296 0 1 62560
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_106_897
timestamp 1636986456
transform 1 0 87400 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_106_909
timestamp 18001
transform 1 0 88504 0 1 62560
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_107_6
timestamp 1636986456
transform 1 0 5428 0 -1 63648
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_18
timestamp 1636986456
transform 1 0 6532 0 -1 63648
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_107_885
timestamp 1636986456
transform 1 0 86296 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_897
timestamp 18001
transform 1 0 87400 0 -1 63648
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_107_905
timestamp 18001
transform 1 0 88136 0 -1 63648
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_108_3
timestamp 1636986456
transform 1 0 5152 0 1 63648
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_15
timestamp 1636986456
transform 1 0 6256 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_108_27
timestamp 18001
transform 1 0 7360 0 1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_108_29
timestamp 18001
transform 1 0 7544 0 1 63648
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_108_885
timestamp 1636986456
transform 1 0 86296 0 1 63648
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_108_897
timestamp 1636986456
transform 1 0 87400 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_108_909
timestamp 18001
transform 1 0 88504 0 1 63648
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_109_6
timestamp 1636986456
transform 1 0 5428 0 -1 64736
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_18
timestamp 1636986456
transform 1 0 6532 0 -1 64736
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_109_885
timestamp 1636986456
transform 1 0 86296 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_109_897
timestamp 18001
transform 1 0 87400 0 -1 64736
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_109_905
timestamp 18001
transform 1 0 88136 0 -1 64736
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_110_6
timestamp 1636986456
transform 1 0 5428 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_110_18
timestamp 18001
transform 1 0 6532 0 1 64736
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_110_26
timestamp 18001
transform 1 0 7268 0 1 64736
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_110_29
timestamp 18001
transform 1 0 7544 0 1 64736
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_110_885
timestamp 1636986456
transform 1 0 86296 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_110_897
timestamp 18001
transform 1 0 87400 0 1 64736
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_110_905
timestamp 18001
transform 1 0 88136 0 1 64736
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_111_3
timestamp 1636986456
transform 1 0 5152 0 -1 65824
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_15
timestamp 1636986456
transform 1 0 6256 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_111_27
timestamp 18001
transform 1 0 7360 0 -1 65824
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_111_885
timestamp 1636986456
transform 1 0 86296 0 -1 65824
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_111_897
timestamp 1636986456
transform 1 0 87400 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_111_909
timestamp 18001
transform 1 0 88504 0 -1 65824
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_112_3
timestamp 1636986456
transform 1 0 5152 0 1 65824
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_15
timestamp 1636986456
transform 1 0 6256 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_112_27
timestamp 18001
transform 1 0 7360 0 1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_112_29
timestamp 18001
transform 1 0 7544 0 1 65824
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_112_885
timestamp 1636986456
transform 1 0 86296 0 1 65824
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_112_897
timestamp 1636986456
transform 1 0 87400 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_112_909
timestamp 18001
transform 1 0 88504 0 1 65824
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_113_7
timestamp 1636986456
transform 1 0 5520 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_113_19
timestamp 18001
transform 1 0 6624 0 -1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_113_27
timestamp 18001
transform 1 0 7360 0 -1 66912
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_113_885
timestamp 1636986456
transform 1 0 86296 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_113_897
timestamp 18001
transform 1 0 87400 0 -1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_113_905
timestamp 18001
transform 1 0 88136 0 -1 66912
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_114_3
timestamp 1636986456
transform 1 0 5152 0 1 66912
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_15
timestamp 1636986456
transform 1 0 6256 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_114_27
timestamp 18001
transform 1 0 7360 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_114_29
timestamp 18001
transform 1 0 7544 0 1 66912
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_114_885
timestamp 1636986456
transform 1 0 86296 0 1 66912
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_114_897
timestamp 1636986456
transform 1 0 87400 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_114_909
timestamp 18001
transform 1 0 88504 0 1 66912
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_115_7
timestamp 1636986456
transform 1 0 5520 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_115_19
timestamp 18001
transform 1 0 6624 0 -1 68000
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_115_27
timestamp 18001
transform 1 0 7360 0 -1 68000
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_115_885
timestamp 1636986456
transform 1 0 86296 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_115_897
timestamp 18001
transform 1 0 87400 0 -1 68000
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_115_905
timestamp 18001
transform 1 0 88136 0 -1 68000
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_116_3
timestamp 1636986456
transform 1 0 5152 0 1 68000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_15
timestamp 1636986456
transform 1 0 6256 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_116_27
timestamp 18001
transform 1 0 7360 0 1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_116_29
timestamp 18001
transform 1 0 7544 0 1 68000
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_116_885
timestamp 1636986456
transform 1 0 86296 0 1 68000
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_116_897
timestamp 1636986456
transform 1 0 87400 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_116_909
timestamp 18001
transform 1 0 88504 0 1 68000
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_117_7
timestamp 1636986456
transform 1 0 5520 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_117_19
timestamp 18001
transform 1 0 6624 0 -1 69088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_117_27
timestamp 18001
transform 1 0 7360 0 -1 69088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_117_885
timestamp 1636986456
transform 1 0 86296 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_117_897
timestamp 18001
transform 1 0 87400 0 -1 69088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_117_905
timestamp 18001
transform 1 0 88136 0 -1 69088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_118_3
timestamp 1636986456
transform 1 0 5152 0 1 69088
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_118_15
timestamp 1636986456
transform 1 0 6256 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_118_27
timestamp 18001
transform 1 0 7360 0 1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_118_29
timestamp 18001
transform 1 0 7544 0 1 69088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_118_885
timestamp 1636986456
transform 1 0 86296 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_118_897
timestamp 18001
transform 1 0 87400 0 1 69088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_118_905
timestamp 18001
transform 1 0 88136 0 1 69088
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_119_7
timestamp 1636986456
transform 1 0 5520 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_119_19
timestamp 18001
transform 1 0 6624 0 -1 70176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_119_27
timestamp 18001
transform 1 0 7360 0 -1 70176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_119_885
timestamp 1636986456
transform 1 0 86296 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_119_897
timestamp 18001
transform 1 0 87400 0 -1 70176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_119_905
timestamp 18001
transform 1 0 88136 0 -1 70176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_120_7
timestamp 1636986456
transform 1 0 5520 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_120_19
timestamp 18001
transform 1 0 6624 0 1 70176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_120_27
timestamp 18001
transform 1 0 7360 0 1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_120_29
timestamp 18001
transform 1 0 7544 0 1 70176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_120_885
timestamp 1636986456
transform 1 0 86296 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_120_897
timestamp 18001
transform 1 0 87400 0 1 70176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_120_905
timestamp 18001
transform 1 0 88136 0 1 70176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_121_3
timestamp 1636986456
transform 1 0 5152 0 -1 71264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_15
timestamp 1636986456
transform 1 0 6256 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_121_27
timestamp 18001
transform 1 0 7360 0 -1 71264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_121_885
timestamp 1636986456
transform 1 0 86296 0 -1 71264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_121_897
timestamp 1636986456
transform 1 0 87400 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_121_909
timestamp 18001
transform 1 0 88504 0 -1 71264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_122_3
timestamp 1636986456
transform 1 0 5152 0 1 71264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_15
timestamp 1636986456
transform 1 0 6256 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_122_27
timestamp 18001
transform 1 0 7360 0 1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_122_29
timestamp 18001
transform 1 0 7544 0 1 71264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_122_885
timestamp 1636986456
transform 1 0 86296 0 1 71264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_122_897
timestamp 1636986456
transform 1 0 87400 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_122_909
timestamp 18001
transform 1 0 88504 0 1 71264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_123_7
timestamp 1636986456
transform 1 0 5520 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_123_19
timestamp 18001
transform 1 0 6624 0 -1 72352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_123_27
timestamp 18001
transform 1 0 7360 0 -1 72352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_123_885
timestamp 1636986456
transform 1 0 86296 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_123_897
timestamp 18001
transform 1 0 87400 0 -1 72352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_123_905
timestamp 18001
transform 1 0 88136 0 -1 72352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_124_3
timestamp 1636986456
transform 1 0 5152 0 1 72352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_15
timestamp 1636986456
transform 1 0 6256 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_124_27
timestamp 18001
transform 1 0 7360 0 1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_124_29
timestamp 18001
transform 1 0 7544 0 1 72352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_124_885
timestamp 1636986456
transform 1 0 86296 0 1 72352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_124_897
timestamp 1636986456
transform 1 0 87400 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_124_909
timestamp 18001
transform 1 0 88504 0 1 72352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_125_7
timestamp 1636986456
transform 1 0 5520 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_125_19
timestamp 18001
transform 1 0 6624 0 -1 73440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_125_27
timestamp 18001
transform 1 0 7360 0 -1 73440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_125_885
timestamp 1636986456
transform 1 0 86296 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_125_897
timestamp 18001
transform 1 0 87400 0 -1 73440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_125_905
timestamp 18001
transform 1 0 88136 0 -1 73440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_126_3
timestamp 1636986456
transform 1 0 5152 0 1 73440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_15
timestamp 1636986456
transform 1 0 6256 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_126_27
timestamp 18001
transform 1 0 7360 0 1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_126_29
timestamp 18001
transform 1 0 7544 0 1 73440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_126_885
timestamp 1636986456
transform 1 0 86296 0 1 73440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_126_897
timestamp 1636986456
transform 1 0 87400 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_126_909
timestamp 18001
transform 1 0 88504 0 1 73440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_127_7
timestamp 1636986456
transform 1 0 5520 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_127_19
timestamp 18001
transform 1 0 6624 0 -1 74528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_127_27
timestamp 18001
transform 1 0 7360 0 -1 74528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_127_885
timestamp 1636986456
transform 1 0 86296 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_127_897
timestamp 18001
transform 1 0 87400 0 -1 74528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_127_905
timestamp 18001
transform 1 0 88136 0 -1 74528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_128_3
timestamp 1636986456
transform 1 0 5152 0 1 74528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_15
timestamp 1636986456
transform 1 0 6256 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_128_27
timestamp 18001
transform 1 0 7360 0 1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_128_29
timestamp 18001
transform 1 0 7544 0 1 74528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_128_885
timestamp 1636986456
transform 1 0 86296 0 1 74528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_128_897
timestamp 1636986456
transform 1 0 87400 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_128_909
timestamp 18001
transform 1 0 88504 0 1 74528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_129_7
timestamp 1636986456
transform 1 0 5520 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_129_19
timestamp 18001
transform 1 0 6624 0 -1 75616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_129_27
timestamp 18001
transform 1 0 7360 0 -1 75616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_129_885
timestamp 1636986456
transform 1 0 86296 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_129_897
timestamp 18001
transform 1 0 87400 0 -1 75616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_129_905
timestamp 18001
transform 1 0 88136 0 -1 75616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_130_7
timestamp 1636986456
transform 1 0 5520 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_130_19
timestamp 18001
transform 1 0 6624 0 1 75616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_130_27
timestamp 18001
transform 1 0 7360 0 1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_130_29
timestamp 18001
transform 1 0 7544 0 1 75616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_130_885
timestamp 1636986456
transform 1 0 86296 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_130_897
timestamp 18001
transform 1 0 87400 0 1 75616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_130_905
timestamp 18001
transform 1 0 88136 0 1 75616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_131_3
timestamp 1636986456
transform 1 0 5152 0 -1 76704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_15
timestamp 1636986456
transform 1 0 6256 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_131_27
timestamp 18001
transform 1 0 7360 0 -1 76704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_131_885
timestamp 1636986456
transform 1 0 86296 0 -1 76704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_131_897
timestamp 1636986456
transform 1 0 87400 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_131_909
timestamp 18001
transform 1 0 88504 0 -1 76704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_132_3
timestamp 1636986456
transform 1 0 5152 0 1 76704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_15
timestamp 1636986456
transform 1 0 6256 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_132_27
timestamp 18001
transform 1 0 7360 0 1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_132_29
timestamp 18001
transform 1 0 7544 0 1 76704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_132_885
timestamp 1636986456
transform 1 0 86296 0 1 76704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_132_897
timestamp 1636986456
transform 1 0 87400 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_132_909
timestamp 18001
transform 1 0 88504 0 1 76704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_133_7
timestamp 1636986456
transform 1 0 5520 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_133_19
timestamp 18001
transform 1 0 6624 0 -1 77792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_133_27
timestamp 18001
transform 1 0 7360 0 -1 77792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_133_885
timestamp 1636986456
transform 1 0 86296 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_133_897
timestamp 18001
transform 1 0 87400 0 -1 77792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_134_3
timestamp 1636986456
transform 1 0 5152 0 1 77792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_15
timestamp 1636986456
transform 1 0 6256 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_134_27
timestamp 18001
transform 1 0 7360 0 1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_134_29
timestamp 18001
transform 1 0 7544 0 1 77792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_134_885
timestamp 1636986456
transform 1 0 86296 0 1 77792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_134_897
timestamp 1636986456
transform 1 0 87400 0 1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_134_909
timestamp 18001
transform 1 0 88504 0 1 77792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_135_7
timestamp 1636986456
transform 1 0 5520 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_135_19
timestamp 18001
transform 1 0 6624 0 -1 78880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_135_27
timestamp 18001
transform 1 0 7360 0 -1 78880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_135_885
timestamp 1636986456
transform 1 0 86296 0 -1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_135_897
timestamp 18001
transform 1 0 87400 0 -1 78880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_135_905
timestamp 18001
transform 1 0 88136 0 -1 78880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_136_3
timestamp 1636986456
transform 1 0 5152 0 1 78880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_15
timestamp 1636986456
transform 1 0 6256 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_136_27
timestamp 18001
transform 1 0 7360 0 1 78880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_136_29
timestamp 18001
transform 1 0 7544 0 1 78880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_136_885
timestamp 1636986456
transform 1 0 86296 0 1 78880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_136_897
timestamp 1636986456
transform 1 0 87400 0 1 78880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_136_909
timestamp 18001
transform 1 0 88504 0 1 78880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_137_7
timestamp 1636986456
transform 1 0 5520 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_137_19
timestamp 18001
transform 1 0 6624 0 -1 79968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_137_27
timestamp 18001
transform 1 0 7360 0 -1 79968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_137_885
timestamp 1636986456
transform 1 0 86296 0 -1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_137_897
timestamp 18001
transform 1 0 87400 0 -1 79968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_137_905
timestamp 18001
transform 1 0 88136 0 -1 79968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_138_3
timestamp 1636986456
transform 1 0 5152 0 1 79968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_15
timestamp 1636986456
transform 1 0 6256 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_138_27
timestamp 18001
transform 1 0 7360 0 1 79968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_138_29
timestamp 18001
transform 1 0 7544 0 1 79968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_138_885
timestamp 1636986456
transform 1 0 86296 0 1 79968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_138_897
timestamp 1636986456
transform 1 0 87400 0 1 79968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_138_909
timestamp 18001
transform 1 0 88504 0 1 79968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_139_7
timestamp 1636986456
transform 1 0 5520 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_139_19
timestamp 18001
transform 1 0 6624 0 -1 81056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_139_27
timestamp 18001
transform 1 0 7360 0 -1 81056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_139_885
timestamp 1636986456
transform 1 0 86296 0 -1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_139_897
timestamp 18001
transform 1 0 87400 0 -1 81056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_140_3
timestamp 1636986456
transform 1 0 5152 0 1 81056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_15
timestamp 1636986456
transform 1 0 6256 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_140_27
timestamp 18001
transform 1 0 7360 0 1 81056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_140_29
timestamp 18001
transform 1 0 7544 0 1 81056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_140_885
timestamp 1636986456
transform 1 0 86296 0 1 81056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_140_897
timestamp 1636986456
transform 1 0 87400 0 1 81056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_140_909
timestamp 18001
transform 1 0 88504 0 1 81056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_141_3
timestamp 1636986456
transform 1 0 5152 0 -1 82144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_15
timestamp 1636986456
transform 1 0 6256 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_141_27
timestamp 18001
transform 1 0 7360 0 -1 82144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_141_885
timestamp 1636986456
transform 1 0 86296 0 -1 82144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_141_897
timestamp 1636986456
transform 1 0 87400 0 -1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_141_909
timestamp 18001
transform 1 0 88504 0 -1 82144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_142_3
timestamp 1636986456
transform 1 0 5152 0 1 82144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_15
timestamp 1636986456
transform 1 0 6256 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_142_27
timestamp 18001
transform 1 0 7360 0 1 82144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_142_29
timestamp 18001
transform 1 0 7544 0 1 82144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_142_885
timestamp 1636986456
transform 1 0 86296 0 1 82144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_142_897
timestamp 1636986456
transform 1 0 87400 0 1 82144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_142_909
timestamp 18001
transform 1 0 88504 0 1 82144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_143_3
timestamp 1636986456
transform 1 0 5152 0 -1 83232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_15
timestamp 1636986456
transform 1 0 6256 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_143_27
timestamp 18001
transform 1 0 7360 0 -1 83232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_143_885
timestamp 1636986456
transform 1 0 86296 0 -1 83232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_143_897
timestamp 1636986456
transform 1 0 87400 0 -1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_143_909
timestamp 18001
transform 1 0 88504 0 -1 83232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_144_3
timestamp 1636986456
transform 1 0 5152 0 1 83232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_15
timestamp 1636986456
transform 1 0 6256 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_144_27
timestamp 18001
transform 1 0 7360 0 1 83232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_144_29
timestamp 18001
transform 1 0 7544 0 1 83232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_144_885
timestamp 1636986456
transform 1 0 86296 0 1 83232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_144_897
timestamp 1636986456
transform 1 0 87400 0 1 83232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_144_909
timestamp 18001
transform 1 0 88504 0 1 83232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_145_3
timestamp 1636986456
transform 1 0 5152 0 -1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_15
timestamp 1636986456
transform 1 0 6256 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_145_27
timestamp 18001
transform 1 0 7360 0 -1 84320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_145_885
timestamp 1636986456
transform 1 0 86296 0 -1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_145_897
timestamp 1636986456
transform 1 0 87400 0 -1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_145_909
timestamp 18001
transform 1 0 88504 0 -1 84320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_146_3
timestamp 1636986456
transform 1 0 5152 0 1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_15
timestamp 1636986456
transform 1 0 6256 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_146_27
timestamp 18001
transform 1 0 7360 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_146_29
timestamp 18001
transform 1 0 7544 0 1 84320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_146_885
timestamp 1636986456
transform 1 0 86296 0 1 84320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_146_897
timestamp 1636986456
transform 1 0 87400 0 1 84320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_146_909
timestamp 18001
transform 1 0 88504 0 1 84320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_147_3
timestamp 1636986456
transform 1 0 5152 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_15
timestamp 1636986456
transform 1 0 6256 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_147_27
timestamp 18001
transform 1 0 7360 0 -1 85408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_147_885
timestamp 1636986456
transform 1 0 86296 0 -1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_147_897
timestamp 1636986456
transform 1 0 87400 0 -1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_147_909
timestamp 18001
transform 1 0 88504 0 -1 85408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_148_3
timestamp 1636986456
transform 1 0 5152 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_15
timestamp 1636986456
transform 1 0 6256 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_148_27
timestamp 18001
transform 1 0 7360 0 1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_148_29
timestamp 18001
transform 1 0 7544 0 1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_148_885
timestamp 1636986456
transform 1 0 86296 0 1 85408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_148_897
timestamp 1636986456
transform 1 0 87400 0 1 85408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_148_909
timestamp 18001
transform 1 0 88504 0 1 85408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_149_3
timestamp 1636986456
transform 1 0 5152 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_15
timestamp 1636986456
transform 1 0 6256 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_149_27
timestamp 18001
transform 1 0 7360 0 -1 86496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_149_885
timestamp 1636986456
transform 1 0 86296 0 -1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_149_897
timestamp 1636986456
transform 1 0 87400 0 -1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_149_909
timestamp 18001
transform 1 0 88504 0 -1 86496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_150_3
timestamp 1636986456
transform 1 0 5152 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_15
timestamp 1636986456
transform 1 0 6256 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_150_27
timestamp 18001
transform 1 0 7360 0 1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_29
timestamp 1636986456
transform 1 0 7544 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_41
timestamp 1636986456
transform 1 0 8648 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_150_53
timestamp 18001
transform 1 0 9752 0 1 86496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_150_57
timestamp 1636986456
transform 1 0 10120 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_69
timestamp 1636986456
transform 1 0 11224 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_150_81
timestamp 18001
transform 1 0 12328 0 1 86496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_150_85
timestamp 1636986456
transform 1 0 12696 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_97
timestamp 1636986456
transform 1 0 13800 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_150_109
timestamp 18001
transform 1 0 14904 0 1 86496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_150_113
timestamp 1636986456
transform 1 0 15272 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_125
timestamp 1636986456
transform 1 0 16376 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_150_137
timestamp 18001
transform 1 0 17480 0 1 86496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_150_141
timestamp 1636986456
transform 1 0 17848 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_153
timestamp 1636986456
transform 1 0 18952 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_150_165
timestamp 18001
transform 1 0 20056 0 1 86496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_150_169
timestamp 1636986456
transform 1 0 20424 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_181
timestamp 1636986456
transform 1 0 21528 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_150_193
timestamp 18001
transform 1 0 22632 0 1 86496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_150_197
timestamp 1636986456
transform 1 0 23000 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_209
timestamp 1636986456
transform 1 0 24104 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_150_221
timestamp 18001
transform 1 0 25208 0 1 86496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_150_225
timestamp 1636986456
transform 1 0 25576 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_237
timestamp 1636986456
transform 1 0 26680 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_150_249
timestamp 18001
transform 1 0 27784 0 1 86496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_150_253
timestamp 18001
transform 1 0 28152 0 1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_259
timestamp 18001
transform 1 0 28704 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_150_301
timestamp 18001
transform 1 0 32568 0 1 86496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_150_307
timestamp 18001
transform 1 0 33120 0 1 86496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_150_309
timestamp 1636986456
transform 1 0 33304 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_321
timestamp 1636986456
transform 1 0 34408 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_150_333
timestamp 18001
transform 1 0 35512 0 1 86496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_150_337
timestamp 1636986456
transform 1 0 35880 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_349
timestamp 1636986456
transform 1 0 36984 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_150_361
timestamp 18001
transform 1 0 38088 0 1 86496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_150_365
timestamp 1636986456
transform 1 0 38456 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_377
timestamp 1636986456
transform 1 0 39560 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_150_389
timestamp 18001
transform 1 0 40664 0 1 86496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_150_393
timestamp 1636986456
transform 1 0 41032 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_405
timestamp 1636986456
transform 1 0 42136 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_150_417
timestamp 18001
transform 1 0 43240 0 1 86496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_150_421
timestamp 1636986456
transform 1 0 43608 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_433
timestamp 1636986456
transform 1 0 44712 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_150_445
timestamp 18001
transform 1 0 45816 0 1 86496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_150_449
timestamp 1636986456
transform 1 0 46184 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_461
timestamp 1636986456
transform 1 0 47288 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_150_473
timestamp 18001
transform 1 0 48392 0 1 86496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_150_477
timestamp 18001
transform 1 0 48760 0 1 86496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_150_485
timestamp 18001
transform 1 0 49496 0 1 86496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_150_505
timestamp 1636986456
transform 1 0 51336 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_517
timestamp 1636986456
transform 1 0 52440 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_150_529
timestamp 18001
transform 1 0 53544 0 1 86496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_150_533
timestamp 1636986456
transform 1 0 53912 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_545
timestamp 1636986456
transform 1 0 55016 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_150_557
timestamp 18001
transform 1 0 56120 0 1 86496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_150_561
timestamp 1636986456
transform 1 0 56488 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_573
timestamp 1636986456
transform 1 0 57592 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_150_585
timestamp 18001
transform 1 0 58696 0 1 86496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_150_589
timestamp 1636986456
transform 1 0 59064 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_601
timestamp 1636986456
transform 1 0 60168 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_150_613
timestamp 18001
transform 1 0 61272 0 1 86496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_150_617
timestamp 1636986456
transform 1 0 61640 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_629
timestamp 1636986456
transform 1 0 62744 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_150_641
timestamp 18001
transform 1 0 63848 0 1 86496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_150_645
timestamp 1636986456
transform 1 0 64216 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_657
timestamp 1636986456
transform 1 0 65320 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_150_669
timestamp 18001
transform 1 0 66424 0 1 86496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_150_673
timestamp 1636986456
transform 1 0 66792 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_685
timestamp 1636986456
transform 1 0 67896 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_150_697
timestamp 18001
transform 1 0 69000 0 1 86496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_150_701
timestamp 1636986456
transform 1 0 69368 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_713
timestamp 1636986456
transform 1 0 70472 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_150_725
timestamp 18001
transform 1 0 71576 0 1 86496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_150_729
timestamp 1636986456
transform 1 0 71944 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_741
timestamp 1636986456
transform 1 0 73048 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_150_753
timestamp 18001
transform 1 0 74152 0 1 86496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_150_757
timestamp 1636986456
transform 1 0 74520 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_769
timestamp 1636986456
transform 1 0 75624 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_150_781
timestamp 18001
transform 1 0 76728 0 1 86496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_150_785
timestamp 1636986456
transform 1 0 77096 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_797
timestamp 1636986456
transform 1 0 78200 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_150_809
timestamp 18001
transform 1 0 79304 0 1 86496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_150_813
timestamp 1636986456
transform 1 0 79672 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_825
timestamp 1636986456
transform 1 0 80776 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_150_837
timestamp 18001
transform 1 0 81880 0 1 86496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_150_841
timestamp 1636986456
transform 1 0 82248 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_853
timestamp 1636986456
transform 1 0 83352 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_150_865
timestamp 18001
transform 1 0 84456 0 1 86496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_150_869
timestamp 1636986456
transform 1 0 84824 0 1 86496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_150_881
timestamp 1636986456
transform 1 0 85928 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_150_893
timestamp 18001
transform 1 0 87032 0 1 86496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_150_897
timestamp 1636986456
transform 1 0 87400 0 1 86496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_150_909
timestamp 18001
transform 1 0 88504 0 1 86496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_151_3
timestamp 1636986456
transform 1 0 5152 0 -1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_15
timestamp 1636986456
transform 1 0 6256 0 -1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_27
timestamp 1636986456
transform 1 0 7360 0 -1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_39
timestamp 1636986456
transform 1 0 8464 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_151_51
timestamp 18001
transform 1 0 9568 0 -1 87584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_151_55
timestamp 18001
transform 1 0 9936 0 -1 87584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_151_57
timestamp 1636986456
transform 1 0 10120 0 -1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_69
timestamp 1636986456
transform 1 0 11224 0 -1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_81
timestamp 1636986456
transform 1 0 12328 0 -1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_93
timestamp 1636986456
transform 1 0 13432 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_151_105
timestamp 18001
transform 1 0 14536 0 -1 87584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_111
timestamp 18001
transform 1 0 15088 0 -1 87584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_151_113
timestamp 1636986456
transform 1 0 15272 0 -1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_125
timestamp 1636986456
transform 1 0 16376 0 -1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_137
timestamp 1636986456
transform 1 0 17480 0 -1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_149
timestamp 1636986456
transform 1 0 18584 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_151_161
timestamp 18001
transform 1 0 19688 0 -1 87584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_167
timestamp 18001
transform 1 0 20240 0 -1 87584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_151_169
timestamp 1636986456
transform 1 0 20424 0 -1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_181
timestamp 1636986456
transform 1 0 21528 0 -1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_193
timestamp 1636986456
transform 1 0 22632 0 -1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_205
timestamp 1636986456
transform 1 0 23736 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_151_217
timestamp 18001
transform 1 0 24840 0 -1 87584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_223
timestamp 18001
transform 1 0 25392 0 -1 87584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_151_225
timestamp 1636986456
transform 1 0 25576 0 -1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_237
timestamp 1636986456
transform 1 0 26680 0 -1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_249
timestamp 1636986456
transform 1 0 27784 0 -1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_261
timestamp 1636986456
transform 1 0 28888 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_151_273
timestamp 18001
transform 1 0 29992 0 -1 87584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_279
timestamp 18001
transform 1 0 30544 0 -1 87584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_151_281
timestamp 1636986456
transform 1 0 30728 0 -1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_293
timestamp 1636986456
transform 1 0 31832 0 -1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_305
timestamp 1636986456
transform 1 0 32936 0 -1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_317
timestamp 1636986456
transform 1 0 34040 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_151_329
timestamp 18001
transform 1 0 35144 0 -1 87584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_335
timestamp 18001
transform 1 0 35696 0 -1 87584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_151_337
timestamp 1636986456
transform 1 0 35880 0 -1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_349
timestamp 1636986456
transform 1 0 36984 0 -1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_361
timestamp 1636986456
transform 1 0 38088 0 -1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_373
timestamp 1636986456
transform 1 0 39192 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_151_385
timestamp 18001
transform 1 0 40296 0 -1 87584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_391
timestamp 18001
transform 1 0 40848 0 -1 87584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_151_393
timestamp 1636986456
transform 1 0 41032 0 -1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_405
timestamp 1636986456
transform 1 0 42136 0 -1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_417
timestamp 1636986456
transform 1 0 43240 0 -1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_429
timestamp 1636986456
transform 1 0 44344 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_151_441
timestamp 18001
transform 1 0 45448 0 -1 87584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_447
timestamp 18001
transform 1 0 46000 0 -1 87584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_151_449
timestamp 1636986456
transform 1 0 46184 0 -1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_461
timestamp 1636986456
transform 1 0 47288 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_151_473
timestamp 18001
transform 1 0 48392 0 -1 87584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_151_481
timestamp 18001
transform 1 0 49128 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_151_498
timestamp 18001
transform 1 0 50692 0 -1 87584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_151_505
timestamp 1636986456
transform 1 0 51336 0 -1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_517
timestamp 1636986456
transform 1 0 52440 0 -1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_529
timestamp 1636986456
transform 1 0 53544 0 -1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_541
timestamp 1636986456
transform 1 0 54648 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_151_553
timestamp 18001
transform 1 0 55752 0 -1 87584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_559
timestamp 18001
transform 1 0 56304 0 -1 87584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_151_561
timestamp 1636986456
transform 1 0 56488 0 -1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_573
timestamp 1636986456
transform 1 0 57592 0 -1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_585
timestamp 1636986456
transform 1 0 58696 0 -1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_597
timestamp 1636986456
transform 1 0 59800 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_151_609
timestamp 18001
transform 1 0 60904 0 -1 87584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_615
timestamp 18001
transform 1 0 61456 0 -1 87584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_151_617
timestamp 1636986456
transform 1 0 61640 0 -1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_629
timestamp 1636986456
transform 1 0 62744 0 -1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_641
timestamp 1636986456
transform 1 0 63848 0 -1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_653
timestamp 1636986456
transform 1 0 64952 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_151_665
timestamp 18001
transform 1 0 66056 0 -1 87584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_671
timestamp 18001
transform 1 0 66608 0 -1 87584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_151_673
timestamp 1636986456
transform 1 0 66792 0 -1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_685
timestamp 1636986456
transform 1 0 67896 0 -1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_697
timestamp 1636986456
transform 1 0 69000 0 -1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_709
timestamp 1636986456
transform 1 0 70104 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_151_721
timestamp 18001
transform 1 0 71208 0 -1 87584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_727
timestamp 18001
transform 1 0 71760 0 -1 87584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_151_729
timestamp 1636986456
transform 1 0 71944 0 -1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_741
timestamp 1636986456
transform 1 0 73048 0 -1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_753
timestamp 1636986456
transform 1 0 74152 0 -1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_765
timestamp 1636986456
transform 1 0 75256 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_151_777
timestamp 18001
transform 1 0 76360 0 -1 87584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_783
timestamp 18001
transform 1 0 76912 0 -1 87584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_151_785
timestamp 1636986456
transform 1 0 77096 0 -1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_797
timestamp 1636986456
transform 1 0 78200 0 -1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_809
timestamp 1636986456
transform 1 0 79304 0 -1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_821
timestamp 1636986456
transform 1 0 80408 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_151_833
timestamp 18001
transform 1 0 81512 0 -1 87584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_839
timestamp 18001
transform 1 0 82064 0 -1 87584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_151_841
timestamp 1636986456
transform 1 0 82248 0 -1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_853
timestamp 1636986456
transform 1 0 83352 0 -1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_865
timestamp 1636986456
transform 1 0 84456 0 -1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_151_877
timestamp 1636986456
transform 1 0 85560 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_151_889
timestamp 18001
transform 1 0 86664 0 -1 87584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_151_895
timestamp 18001
transform 1 0 87216 0 -1 87584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_151_897
timestamp 1636986456
transform 1 0 87400 0 -1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_151_909
timestamp 18001
transform 1 0 88504 0 -1 87584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_152_3
timestamp 1636986456
transform 1 0 5152 0 1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_15
timestamp 1636986456
transform 1 0 6256 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_152_27
timestamp 18001
transform 1 0 7360 0 1 87584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_152_29
timestamp 1636986456
transform 1 0 7544 0 1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_41
timestamp 1636986456
transform 1 0 8648 0 1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_53
timestamp 1636986456
transform 1 0 9752 0 1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_65
timestamp 1636986456
transform 1 0 10856 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_77
timestamp 18001
transform 1 0 11960 0 1 87584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_152_83
timestamp 18001
transform 1 0 12512 0 1 87584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_152_85
timestamp 1636986456
transform 1 0 12696 0 1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_97
timestamp 1636986456
transform 1 0 13800 0 1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_109
timestamp 1636986456
transform 1 0 14904 0 1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_121
timestamp 1636986456
transform 1 0 16008 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_133
timestamp 18001
transform 1 0 17112 0 1 87584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_152_139
timestamp 18001
transform 1 0 17664 0 1 87584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_152_141
timestamp 1636986456
transform 1 0 17848 0 1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_153
timestamp 1636986456
transform 1 0 18952 0 1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_165
timestamp 1636986456
transform 1 0 20056 0 1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_177
timestamp 1636986456
transform 1 0 21160 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_189
timestamp 18001
transform 1 0 22264 0 1 87584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_152_195
timestamp 18001
transform 1 0 22816 0 1 87584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_152_197
timestamp 1636986456
transform 1 0 23000 0 1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_209
timestamp 1636986456
transform 1 0 24104 0 1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_221
timestamp 1636986456
transform 1 0 25208 0 1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_233
timestamp 1636986456
transform 1 0 26312 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_245
timestamp 18001
transform 1 0 27416 0 1 87584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_152_251
timestamp 18001
transform 1 0 27968 0 1 87584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_152_253
timestamp 1636986456
transform 1 0 28152 0 1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_265
timestamp 1636986456
transform 1 0 29256 0 1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_277
timestamp 1636986456
transform 1 0 30360 0 1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_289
timestamp 1636986456
transform 1 0 31464 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_301
timestamp 18001
transform 1 0 32568 0 1 87584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_152_307
timestamp 18001
transform 1 0 33120 0 1 87584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_152_309
timestamp 1636986456
transform 1 0 33304 0 1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_321
timestamp 1636986456
transform 1 0 34408 0 1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_333
timestamp 1636986456
transform 1 0 35512 0 1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_345
timestamp 1636986456
transform 1 0 36616 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_357
timestamp 18001
transform 1 0 37720 0 1 87584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_152_363
timestamp 18001
transform 1 0 38272 0 1 87584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_152_365
timestamp 1636986456
transform 1 0 38456 0 1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_377
timestamp 1636986456
transform 1 0 39560 0 1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_389
timestamp 1636986456
transform 1 0 40664 0 1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_401
timestamp 1636986456
transform 1 0 41768 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_413
timestamp 18001
transform 1 0 42872 0 1 87584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_152_419
timestamp 18001
transform 1 0 43424 0 1 87584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_152_421
timestamp 1636986456
transform 1 0 43608 0 1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_433
timestamp 1636986456
transform 1 0 44712 0 1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_445
timestamp 1636986456
transform 1 0 45816 0 1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_457
timestamp 1636986456
transform 1 0 46920 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_469
timestamp 18001
transform 1 0 48024 0 1 87584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_152_475
timestamp 18001
transform 1 0 48576 0 1 87584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_152_477
timestamp 1636986456
transform 1 0 48760 0 1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_489
timestamp 1636986456
transform 1 0 49864 0 1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_501
timestamp 1636986456
transform 1 0 50968 0 1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_513
timestamp 1636986456
transform 1 0 52072 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_525
timestamp 18001
transform 1 0 53176 0 1 87584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_152_531
timestamp 18001
transform 1 0 53728 0 1 87584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_152_533
timestamp 1636986456
transform 1 0 53912 0 1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_545
timestamp 1636986456
transform 1 0 55016 0 1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_557
timestamp 1636986456
transform 1 0 56120 0 1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_569
timestamp 1636986456
transform 1 0 57224 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_581
timestamp 18001
transform 1 0 58328 0 1 87584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_152_587
timestamp 18001
transform 1 0 58880 0 1 87584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_152_589
timestamp 1636986456
transform 1 0 59064 0 1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_601
timestamp 1636986456
transform 1 0 60168 0 1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_613
timestamp 1636986456
transform 1 0 61272 0 1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_625
timestamp 1636986456
transform 1 0 62376 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_637
timestamp 18001
transform 1 0 63480 0 1 87584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_152_643
timestamp 18001
transform 1 0 64032 0 1 87584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_152_645
timestamp 1636986456
transform 1 0 64216 0 1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_657
timestamp 1636986456
transform 1 0 65320 0 1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_669
timestamp 1636986456
transform 1 0 66424 0 1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_681
timestamp 1636986456
transform 1 0 67528 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_693
timestamp 18001
transform 1 0 68632 0 1 87584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_152_699
timestamp 18001
transform 1 0 69184 0 1 87584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_152_701
timestamp 1636986456
transform 1 0 69368 0 1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_713
timestamp 1636986456
transform 1 0 70472 0 1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_725
timestamp 1636986456
transform 1 0 71576 0 1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_737
timestamp 1636986456
transform 1 0 72680 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_749
timestamp 18001
transform 1 0 73784 0 1 87584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_152_755
timestamp 18001
transform 1 0 74336 0 1 87584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_152_757
timestamp 1636986456
transform 1 0 74520 0 1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_769
timestamp 1636986456
transform 1 0 75624 0 1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_781
timestamp 1636986456
transform 1 0 76728 0 1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_793
timestamp 1636986456
transform 1 0 77832 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_805
timestamp 18001
transform 1 0 78936 0 1 87584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_152_811
timestamp 18001
transform 1 0 79488 0 1 87584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_152_813
timestamp 1636986456
transform 1 0 79672 0 1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_825
timestamp 1636986456
transform 1 0 80776 0 1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_837
timestamp 1636986456
transform 1 0 81880 0 1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_849
timestamp 1636986456
transform 1 0 82984 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_861
timestamp 18001
transform 1 0 84088 0 1 87584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_152_867
timestamp 18001
transform 1 0 84640 0 1 87584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_152_869
timestamp 1636986456
transform 1 0 84824 0 1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_881
timestamp 1636986456
transform 1 0 85928 0 1 87584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_152_893
timestamp 1636986456
transform 1 0 87032 0 1 87584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_152_905
timestamp 18001
transform 1 0 88136 0 1 87584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_153_3
timestamp 1636986456
transform 1 0 5152 0 -1 88672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_15
timestamp 1636986456
transform 1 0 6256 0 -1 88672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_27
timestamp 1636986456
transform 1 0 7360 0 -1 88672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_39
timestamp 1636986456
transform 1 0 8464 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_153_51
timestamp 18001
transform 1 0 9568 0 -1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_153_55
timestamp 18001
transform 1 0 9936 0 -1 88672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_153_57
timestamp 1636986456
transform 1 0 10120 0 -1 88672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_69
timestamp 1636986456
transform 1 0 11224 0 -1 88672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_81
timestamp 1636986456
transform 1 0 12328 0 -1 88672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_93
timestamp 1636986456
transform 1 0 13432 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_153_105
timestamp 18001
transform 1 0 14536 0 -1 88672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_153_111
timestamp 18001
transform 1 0 15088 0 -1 88672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_153_113
timestamp 1636986456
transform 1 0 15272 0 -1 88672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_125
timestamp 1636986456
transform 1 0 16376 0 -1 88672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_137
timestamp 1636986456
transform 1 0 17480 0 -1 88672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_149
timestamp 1636986456
transform 1 0 18584 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_153_161
timestamp 18001
transform 1 0 19688 0 -1 88672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_153_167
timestamp 18001
transform 1 0 20240 0 -1 88672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_153_169
timestamp 1636986456
transform 1 0 20424 0 -1 88672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_181
timestamp 1636986456
transform 1 0 21528 0 -1 88672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_193
timestamp 1636986456
transform 1 0 22632 0 -1 88672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_205
timestamp 1636986456
transform 1 0 23736 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_153_217
timestamp 18001
transform 1 0 24840 0 -1 88672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_153_223
timestamp 18001
transform 1 0 25392 0 -1 88672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_153_225
timestamp 1636986456
transform 1 0 25576 0 -1 88672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_237
timestamp 1636986456
transform 1 0 26680 0 -1 88672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_249
timestamp 1636986456
transform 1 0 27784 0 -1 88672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_261
timestamp 1636986456
transform 1 0 28888 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_153_273
timestamp 18001
transform 1 0 29992 0 -1 88672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_153_279
timestamp 18001
transform 1 0 30544 0 -1 88672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_153_281
timestamp 1636986456
transform 1 0 30728 0 -1 88672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_293
timestamp 1636986456
transform 1 0 31832 0 -1 88672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_305
timestamp 1636986456
transform 1 0 32936 0 -1 88672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_317
timestamp 1636986456
transform 1 0 34040 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_153_329
timestamp 18001
transform 1 0 35144 0 -1 88672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_153_335
timestamp 18001
transform 1 0 35696 0 -1 88672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_153_337
timestamp 1636986456
transform 1 0 35880 0 -1 88672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_349
timestamp 1636986456
transform 1 0 36984 0 -1 88672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_361
timestamp 1636986456
transform 1 0 38088 0 -1 88672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_373
timestamp 1636986456
transform 1 0 39192 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_153_385
timestamp 18001
transform 1 0 40296 0 -1 88672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_153_391
timestamp 18001
transform 1 0 40848 0 -1 88672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_153_393
timestamp 1636986456
transform 1 0 41032 0 -1 88672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_405
timestamp 1636986456
transform 1 0 42136 0 -1 88672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_417
timestamp 1636986456
transform 1 0 43240 0 -1 88672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_429
timestamp 1636986456
transform 1 0 44344 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_153_441
timestamp 18001
transform 1 0 45448 0 -1 88672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_153_447
timestamp 18001
transform 1 0 46000 0 -1 88672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_153_449
timestamp 1636986456
transform 1 0 46184 0 -1 88672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_461
timestamp 1636986456
transform 1 0 47288 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_153_473
timestamp 18001
transform 1 0 48392 0 -1 88672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_153_492
timestamp 1636986456
transform 1 0 50140 0 -1 88672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_505
timestamp 1636986456
transform 1 0 51336 0 -1 88672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_517
timestamp 1636986456
transform 1 0 52440 0 -1 88672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_529
timestamp 1636986456
transform 1 0 53544 0 -1 88672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_541
timestamp 1636986456
transform 1 0 54648 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_153_553
timestamp 18001
transform 1 0 55752 0 -1 88672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_153_559
timestamp 18001
transform 1 0 56304 0 -1 88672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_153_561
timestamp 1636986456
transform 1 0 56488 0 -1 88672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_573
timestamp 1636986456
transform 1 0 57592 0 -1 88672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_585
timestamp 1636986456
transform 1 0 58696 0 -1 88672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_597
timestamp 1636986456
transform 1 0 59800 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_153_609
timestamp 18001
transform 1 0 60904 0 -1 88672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_153_615
timestamp 18001
transform 1 0 61456 0 -1 88672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_153_617
timestamp 1636986456
transform 1 0 61640 0 -1 88672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_629
timestamp 1636986456
transform 1 0 62744 0 -1 88672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_641
timestamp 1636986456
transform 1 0 63848 0 -1 88672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_653
timestamp 1636986456
transform 1 0 64952 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_153_665
timestamp 18001
transform 1 0 66056 0 -1 88672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_153_671
timestamp 18001
transform 1 0 66608 0 -1 88672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_153_673
timestamp 1636986456
transform 1 0 66792 0 -1 88672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_685
timestamp 1636986456
transform 1 0 67896 0 -1 88672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_697
timestamp 1636986456
transform 1 0 69000 0 -1 88672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_709
timestamp 1636986456
transform 1 0 70104 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_153_721
timestamp 18001
transform 1 0 71208 0 -1 88672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_153_727
timestamp 18001
transform 1 0 71760 0 -1 88672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_153_729
timestamp 1636986456
transform 1 0 71944 0 -1 88672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_741
timestamp 1636986456
transform 1 0 73048 0 -1 88672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_753
timestamp 1636986456
transform 1 0 74152 0 -1 88672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_765
timestamp 1636986456
transform 1 0 75256 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_153_777
timestamp 18001
transform 1 0 76360 0 -1 88672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_153_783
timestamp 18001
transform 1 0 76912 0 -1 88672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_153_785
timestamp 1636986456
transform 1 0 77096 0 -1 88672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_797
timestamp 1636986456
transform 1 0 78200 0 -1 88672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_809
timestamp 1636986456
transform 1 0 79304 0 -1 88672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_821
timestamp 1636986456
transform 1 0 80408 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_153_833
timestamp 18001
transform 1 0 81512 0 -1 88672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_153_839
timestamp 18001
transform 1 0 82064 0 -1 88672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_153_841
timestamp 1636986456
transform 1 0 82248 0 -1 88672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_853
timestamp 1636986456
transform 1 0 83352 0 -1 88672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_865
timestamp 1636986456
transform 1 0 84456 0 -1 88672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_153_877
timestamp 1636986456
transform 1 0 85560 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_153_889
timestamp 18001
transform 1 0 86664 0 -1 88672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_153_895
timestamp 18001
transform 1 0 87216 0 -1 88672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_153_897
timestamp 1636986456
transform 1 0 87400 0 -1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_153_909
timestamp 18001
transform 1 0 88504 0 -1 88672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_154_3
timestamp 1636986456
transform 1 0 5152 0 1 88672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_15
timestamp 1636986456
transform 1 0 6256 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_154_27
timestamp 18001
transform 1 0 7360 0 1 88672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_154_29
timestamp 1636986456
transform 1 0 7544 0 1 88672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_41
timestamp 1636986456
transform 1 0 8648 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_154_53
timestamp 18001
transform 1 0 9752 0 1 88672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_154_57
timestamp 1636986456
transform 1 0 10120 0 1 88672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_69
timestamp 1636986456
transform 1 0 11224 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_154_81
timestamp 18001
transform 1 0 12328 0 1 88672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_154_85
timestamp 1636986456
transform 1 0 12696 0 1 88672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_97
timestamp 1636986456
transform 1 0 13800 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_154_109
timestamp 18001
transform 1 0 14904 0 1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_154_113
timestamp 18001
transform 1 0 15272 0 1 88672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_154_123
timestamp 18001
transform 1 0 16192 0 1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_154_130
timestamp 18001
transform 1 0 16836 0 1 88672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_154_138
timestamp 18001
transform 1 0 17572 0 1 88672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_154_147
timestamp 18001
transform 1 0 18400 0 1 88672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_154_153
timestamp 18001
transform 1 0 18952 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_154_158
timestamp 18001
transform 1 0 19412 0 1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_154_165
timestamp 18001
transform 1 0 20056 0 1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_154_169
timestamp 18001
transform 1 0 20424 0 1 88672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_154_179
timestamp 18001
transform 1 0 21344 0 1 88672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_154_187
timestamp 18001
transform 1 0 22080 0 1 88672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_154_193
timestamp 18001
transform 1 0 22632 0 1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_154_197
timestamp 18001
transform 1 0 23000 0 1 88672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_154_207
timestamp 18001
transform 1 0 23920 0 1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_154_216
timestamp 18001
transform 1 0 24748 0 1 88672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_154_235
timestamp 18001
transform 1 0 26496 0 1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_154_244
timestamp 18001
transform 1 0 27324 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_154_251
timestamp 18001
transform 1 0 27968 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_154_253
timestamp 18001
transform 1 0 28152 0 1 88672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_154_263
timestamp 18001
transform 1 0 29072 0 1 88672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_154_271
timestamp 18001
transform 1 0 29808 0 1 88672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_154_276
timestamp 18001
transform 1 0 30268 0 1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_154_281
timestamp 18001
transform 1 0 30728 0 1 88672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_154_291
timestamp 18001
transform 1 0 31648 0 1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_154_298
timestamp 18001
transform 1 0 32292 0 1 88672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_154_306
timestamp 18001
transform 1 0 33028 0 1 88672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_154_313
timestamp 18001
transform 1 0 33672 0 1 88672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_154_321
timestamp 18001
transform 1 0 34408 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_154_326
timestamp 18001
transform 1 0 34868 0 1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_154_333
timestamp 18001
transform 1 0 35512 0 1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_154_337
timestamp 18001
transform 1 0 35880 0 1 88672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_154_347
timestamp 18001
transform 1 0 36800 0 1 88672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_154_355
timestamp 18001
transform 1 0 37536 0 1 88672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_154_361
timestamp 18001
transform 1 0 38088 0 1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_154_365
timestamp 18001
transform 1 0 38456 0 1 88672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_154_375
timestamp 18001
transform 1 0 39376 0 1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_154_382
timestamp 18001
transform 1 0 40020 0 1 88672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_154_390
timestamp 18001
transform 1 0 40756 0 1 88672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_154_397
timestamp 18001
transform 1 0 41400 0 1 88672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_154_405
timestamp 18001
transform 1 0 42136 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_154_410
timestamp 18001
transform 1 0 42596 0 1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_154_417
timestamp 18001
transform 1 0 43240 0 1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_154_421
timestamp 18001
transform 1 0 43608 0 1 88672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_154_431
timestamp 18001
transform 1 0 44528 0 1 88672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_154_439
timestamp 18001
transform 1 0 45264 0 1 88672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_154_445
timestamp 18001
transform 1 0 45816 0 1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_154_449
timestamp 18001
transform 1 0 46184 0 1 88672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_154_458
timestamp 1636986456
transform 1 0 47012 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_154_470
timestamp 18001
transform 1 0 48116 0 1 88672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_154_477
timestamp 18001
transform 1 0 48760 0 1 88672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_154_485
timestamp 18001
transform 1 0 49496 0 1 88672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_154_505
timestamp 1636986456
transform 1 0 51336 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_154_517
timestamp 18001
transform 1 0 52440 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_154_522
timestamp 18001
transform 1 0 52900 0 1 88672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_154_530
timestamp 18001
transform 1 0 53636 0 1 88672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_154_537
timestamp 18001
transform 1 0 54280 0 1 88672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_154_545
timestamp 18001
transform 1 0 55016 0 1 88672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_154_557
timestamp 18001
transform 1 0 56120 0 1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_154_564
timestamp 18001
transform 1 0 56764 0 1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_154_571
timestamp 18001
transform 1 0 57408 0 1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_154_577
timestamp 18001
transform 1 0 57960 0 1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_154_585
timestamp 18001
transform 1 0 58696 0 1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_154_593
timestamp 18001
transform 1 0 59432 0 1 88672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_154_601
timestamp 18001
transform 1 0 60168 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_154_606
timestamp 18001
transform 1 0 60628 0 1 88672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_154_614
timestamp 18001
transform 1 0 61364 0 1 88672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_154_633
timestamp 18001
transform 1 0 63112 0 1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_154_643
timestamp 18001
transform 1 0 64032 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_154_645
timestamp 18001
transform 1 0 64216 0 1 88672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_154_657
timestamp 18001
transform 1 0 65320 0 1 88672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_154_669
timestamp 18001
transform 1 0 66424 0 1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_154_676
timestamp 18001
transform 1 0 67068 0 1 88672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_154_684
timestamp 18001
transform 1 0 67804 0 1 88672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_154_690
timestamp 18001
transform 1 0 68356 0 1 88672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_154_698
timestamp 18001
transform 1 0 69092 0 1 88672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_154_705
timestamp 18001
transform 1 0 69736 0 1 88672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_154_711
timestamp 18001
transform 1 0 70288 0 1 88672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_154_719
timestamp 18001
transform 1 0 71024 0 1 88672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_154_725
timestamp 18001
transform 1 0 71576 0 1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_154_729
timestamp 18001
transform 1 0 71944 0 1 88672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_154_739
timestamp 18001
transform 1 0 72864 0 1 88672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_154_747
timestamp 18001
transform 1 0 73600 0 1 88672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_154_753
timestamp 18001
transform 1 0 74152 0 1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_154_761
timestamp 18001
transform 1 0 74888 0 1 88672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_154_769
timestamp 18001
transform 1 0 75624 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_154_774
timestamp 18001
transform 1 0 76084 0 1 88672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_154_782
timestamp 18001
transform 1 0 76820 0 1 88672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_154_789
timestamp 18001
transform 1 0 77464 0 1 88672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_154_795
timestamp 18001
transform 1 0 78016 0 1 88672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_154_803
timestamp 18001
transform 1 0 78752 0 1 88672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_154_809
timestamp 18001
transform 1 0 79304 0 1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_154_813
timestamp 18001
transform 1 0 79672 0 1 88672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_154_823
timestamp 18001
transform 1 0 80592 0 1 88672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_154_831
timestamp 18001
transform 1 0 81328 0 1 88672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_154_837
timestamp 18001
transform 1 0 81880 0 1 88672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_154_845
timestamp 1636986456
transform 1 0 82616 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_154_857
timestamp 18001
transform 1 0 83720 0 1 88672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_154_865
timestamp 18001
transform 1 0 84456 0 1 88672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_154_869
timestamp 1636986456
transform 1 0 84824 0 1 88672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_154_881
timestamp 1636986456
transform 1 0 85928 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_154_893
timestamp 18001
transform 1 0 87032 0 1 88672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_154_897
timestamp 1636986456
transform 1 0 87400 0 1 88672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_154_909
timestamp 18001
transform 1 0 88504 0 1 88672
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  fpga_234
timestamp 18001
transform -1 0 5428 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_235
timestamp 18001
transform -1 0 5428 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_236
timestamp 18001
transform -1 0 5428 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_237
timestamp 18001
transform -1 0 5428 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_238
timestamp 18001
transform -1 0 56764 0 1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_239
timestamp 18001
transform 1 0 88320 0 1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_240
timestamp 18001
transform 1 0 88412 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_241
timestamp 18001
transform -1 0 57960 0 1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_242
timestamp 18001
transform 1 0 88320 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_243
timestamp 18001
transform -1 0 5428 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_244
timestamp 18001
transform 1 0 88320 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_245
timestamp 18001
transform 1 0 88320 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_246
timestamp 18001
transform -1 0 47012 0 1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_247
timestamp 18001
transform -1 0 5428 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_248
timestamp 18001
transform -1 0 5428 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  fpga_249
timestamp 18001
transform -1 0 5428 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input1
timestamp 18001
transform 1 0 5152 0 -1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__buf_12  input2
timestamp 18001
transform 1 0 49772 0 1 88672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 18001
transform -1 0 88596 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input4
timestamp 18001
transform -1 0 88596 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input5
timestamp 18001
transform -1 0 88688 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input6
timestamp 18001
transform -1 0 88596 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input7
timestamp 18001
transform -1 0 88596 0 1 42976
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 18001
transform -1 0 88688 0 -1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 18001
transform -1 0 88688 0 -1 68000
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 18001
transform -1 0 88688 0 -1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp 18001
transform -1 0 88688 0 -1 70176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 18001
transform -1 0 88688 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 18001
transform -1 0 88596 0 1 70176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 18001
transform -1 0 88688 0 -1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 18001
transform -1 0 88688 0 -1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 18001
transform -1 0 88688 0 -1 74528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 18001
transform -1 0 88688 0 -1 75616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input18
timestamp 18001
transform -1 0 88596 0 1 75616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input19
timestamp 18001
transform -1 0 88688 0 -1 77792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input20
timestamp 18001
transform -1 0 88688 0 -1 78880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input21
timestamp 18001
transform -1 0 88688 0 -1 79968
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input22
timestamp 18001
transform -1 0 88688 0 -1 81056
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input23
timestamp 18001
transform -1 0 88596 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 18001
transform -1 0 88596 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input25
timestamp 18001
transform -1 0 88596 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input26
timestamp 18001
transform -1 0 88596 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input27
timestamp 18001
transform -1 0 88688 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input28
timestamp 18001
transform -1 0 88596 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input29
timestamp 18001
transform -1 0 88596 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input30
timestamp 18001
transform -1 0 88596 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input31
timestamp 18001
transform 1 0 15824 0 1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input32
timestamp 18001
transform 1 0 26772 0 1 88672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input33
timestamp 18001
transform 1 0 27416 0 1 88672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input34
timestamp 18001
transform 1 0 28704 0 1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input35
timestamp 18001
transform -1 0 30268 0 1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input36
timestamp 18001
transform 1 0 52532 0 1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input37
timestamp 18001
transform 1 0 53912 0 1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input38
timestamp 18001
transform 1 0 54464 0 1 88672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input39
timestamp 18001
transform 1 0 55752 0 1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input40
timestamp 18001
transform 1 0 16468 0 1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input41
timestamp 18001
transform 1 0 57040 0 1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input42
timestamp 18001
transform -1 0 58696 0 1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input43
timestamp 18001
transform 1 0 59064 0 1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input44
timestamp 18001
transform 1 0 60260 0 1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input45
timestamp 18001
transform 1 0 61640 0 1 88672
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input46
timestamp 18001
transform 1 0 62192 0 1 88672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  input47
timestamp 18001
transform 1 0 63480 0 1 88672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input48
timestamp 18001
transform 1 0 64768 0 1 88672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input49
timestamp 18001
transform 1 0 66056 0 1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input50
timestamp 18001
transform 1 0 66792 0 1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input51
timestamp 18001
transform 1 0 17848 0 1 88672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input52
timestamp 18001
transform 1 0 19044 0 1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input53
timestamp 18001
transform 1 0 19688 0 1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input54
timestamp 18001
transform -1 0 21344 0 1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input55
timestamp 18001
transform 1 0 22264 0 1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input56
timestamp 18001
transform 1 0 23552 0 1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input57
timestamp 18001
transform 1 0 24196 0 1 88672
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input58
timestamp 18001
transform 1 0 25576 0 1 88672
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input59
timestamp 18001
transform -1 0 31556 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input60
timestamp 18001
transform -1 0 42596 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input61
timestamp 18001
transform 1 0 42872 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input62
timestamp 18001
transform 1 0 44160 0 1 4896
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input63
timestamp 18001
transform 1 0 46184 0 1 4896
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input64
timestamp 18001
transform -1 0 68264 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input65
timestamp 18001
transform -1 0 69644 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input66
timestamp 18001
transform 1 0 69920 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input67
timestamp 18001
transform 1 0 71208 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input68
timestamp 18001
transform 1 0 31924 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input69
timestamp 18001
transform -1 0 72772 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input70
timestamp 18001
transform -1 0 74060 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input71
timestamp 18001
transform 1 0 74520 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input72
timestamp 18001
transform -1 0 75992 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input73
timestamp 18001
transform -1 0 77372 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input74
timestamp 18001
transform 1 0 77648 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input75
timestamp 18001
transform 1 0 78936 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input76
timestamp 18001
transform -1 0 80592 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input77
timestamp 18001
transform 1 0 82248 0 1 4896
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input78
timestamp 18001
transform 1 0 82248 0 -1 5984
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input79
timestamp 18001
transform -1 0 33580 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input80
timestamp 18001
transform -1 0 34776 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input81
timestamp 18001
transform 1 0 35144 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input82
timestamp 18001
transform 1 0 36432 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input83
timestamp 18001
transform -1 0 37996 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input84
timestamp 18001
transform -1 0 39284 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input85
timestamp 18001
transform 1 0 39652 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input86
timestamp 18001
transform -1 0 41308 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input87
timestamp 18001
transform 1 0 5152 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input88
timestamp 18001
transform 1 0 5152 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input89
timestamp 18001
transform 1 0 5152 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input90
timestamp 18001
transform 1 0 5152 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input91
timestamp 18001
transform 1 0 5152 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input92
timestamp 18001
transform 1 0 5152 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input93
timestamp 18001
transform -1 0 5428 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input94
timestamp 18001
transform -1 0 5428 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input95
timestamp 18001
transform 1 0 5152 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input96
timestamp 18001
transform -1 0 5428 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input97
timestamp 18001
transform 1 0 5152 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input98
timestamp 18001
transform 1 0 5152 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input99
timestamp 18001
transform 1 0 5152 0 -1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input100
timestamp 18001
transform 1 0 5152 0 -1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input101
timestamp 18001
transform 1 0 5152 0 1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input102
timestamp 18001
transform 1 0 5152 0 -1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input103
timestamp 18001
transform 1 0 5152 0 -1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input104
timestamp 18001
transform 1 0 5152 0 -1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input105
timestamp 18001
transform 1 0 5152 0 -1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input106
timestamp 18001
transform 1 0 5152 0 1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input107
timestamp 18001
transform -1 0 5428 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input108
timestamp 18001
transform 1 0 5152 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input109
timestamp 18001
transform 1 0 5152 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input110
timestamp 18001
transform 1 0 5152 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input111
timestamp 18001
transform 1 0 5152 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input112
timestamp 18001
transform 1 0 5152 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input113
timestamp 18001
transform 1 0 5152 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input114
timestamp 18001
transform 1 0 5152 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  input115
timestamp 18001
transform 1 0 12696 0 1 4896
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  input116
timestamp 18001
transform 1 0 13892 0 1 4896
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  input117
timestamp 18001
transform 1 0 15272 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__buf_12  input118
timestamp 18001
transform 1 0 48668 0 -1 88672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  max_cap232
timestamp 18001
transform 1 0 49772 0 1 86496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  max_cap233
timestamp 18001
transform 1 0 49220 0 -1 87584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  output119
timestamp 18001
transform 1 0 88320 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output120
timestamp 18001
transform 1 0 88320 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output121
timestamp 18001
transform 1 0 88320 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output122
timestamp 18001
transform 1 0 88228 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output123
timestamp 18001
transform 1 0 88228 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output124
timestamp 18001
transform 1 0 88228 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output125
timestamp 18001
transform 1 0 88320 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output126
timestamp 18001
transform 1 0 88320 0 -1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output127
timestamp 18001
transform 1 0 88320 0 -1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output128
timestamp 18001
transform 1 0 88228 0 1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output129
timestamp 18001
transform 1 0 88228 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output130
timestamp 18001
transform 1 0 88320 0 -1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output131
timestamp 18001
transform 1 0 88320 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output132
timestamp 18001
transform 1 0 88320 0 -1 58208
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output133
timestamp 18001
transform 1 0 88320 0 -1 59296
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output134
timestamp 18001
transform 1 0 88228 0 1 59296
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output135
timestamp 18001
transform 1 0 88320 0 -1 61472
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output136
timestamp 18001
transform 1 0 88320 0 -1 62560
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output137
timestamp 18001
transform 1 0 88320 0 -1 63648
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output138
timestamp 18001
transform 1 0 88320 0 -1 64736
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output139
timestamp 18001
transform 1 0 88228 0 1 64736
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output140
timestamp 18001
transform 1 0 88228 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output141
timestamp 18001
transform 1 0 88228 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output142
timestamp 18001
transform 1 0 88228 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output143
timestamp 18001
transform 1 0 88320 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output144
timestamp 18001
transform 1 0 88228 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output145
timestamp 18001
transform 1 0 88228 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output146
timestamp 18001
transform 1 0 88228 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output147
timestamp 18001
transform 1 0 88228 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output148
timestamp 18001
transform 1 0 31280 0 1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output149
timestamp 18001
transform 1 0 42228 0 1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output150
timestamp 18001
transform -1 0 43240 0 1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output151
timestamp 18001
transform 1 0 44160 0 1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output152
timestamp 18001
transform 1 0 45448 0 1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output153
timestamp 18001
transform 1 0 67988 0 1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output154
timestamp 18001
transform 1 0 69368 0 1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output155
timestamp 18001
transform -1 0 70288 0 1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output156
timestamp 18001
transform 1 0 71208 0 1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output157
timestamp 18001
transform -1 0 32292 0 1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output158
timestamp 18001
transform 1 0 72496 0 1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output159
timestamp 18001
transform 1 0 73784 0 1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output160
timestamp 18001
transform 1 0 74520 0 1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output161
timestamp 18001
transform 1 0 75716 0 1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output162
timestamp 18001
transform 1 0 77096 0 1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output163
timestamp 18001
transform -1 0 78016 0 1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output164
timestamp 18001
transform 1 0 78936 0 1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output165
timestamp 18001
transform 1 0 80224 0 1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output166
timestamp 18001
transform 1 0 81512 0 1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output167
timestamp 18001
transform 1 0 82248 0 1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output168
timestamp 18001
transform 1 0 33304 0 1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output169
timestamp 18001
transform 1 0 34500 0 1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output170
timestamp 18001
transform -1 0 35512 0 1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output171
timestamp 18001
transform 1 0 36432 0 1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output172
timestamp 18001
transform 1 0 37720 0 1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output173
timestamp 18001
transform 1 0 39008 0 1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output174
timestamp 18001
transform -1 0 40020 0 1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output175
timestamp 18001
transform 1 0 41032 0 1 88672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output176
timestamp 18001
transform 1 0 15824 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output177
timestamp 18001
transform 1 0 26772 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output178
timestamp 18001
transform -1 0 27784 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output179
timestamp 18001
transform 1 0 28704 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output180
timestamp 18001
transform 1 0 29992 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output181
timestamp 18001
transform 1 0 52532 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output182
timestamp 18001
transform 1 0 53912 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output183
timestamp 18001
transform -1 0 54832 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output184
timestamp 18001
transform 1 0 55752 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output185
timestamp 18001
transform -1 0 16836 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output186
timestamp 18001
transform 1 0 57040 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output187
timestamp 18001
transform 1 0 58328 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output188
timestamp 18001
transform 1 0 59064 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output189
timestamp 18001
transform 1 0 60260 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output190
timestamp 18001
transform 1 0 61640 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output191
timestamp 18001
transform -1 0 62560 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output192
timestamp 18001
transform 1 0 63480 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output193
timestamp 18001
transform 1 0 64768 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output194
timestamp 18001
transform 1 0 66056 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output195
timestamp 18001
transform 1 0 66792 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output196
timestamp 18001
transform 1 0 17848 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output197
timestamp 18001
transform 1 0 19044 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output198
timestamp 18001
transform -1 0 20056 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output199
timestamp 18001
transform 1 0 20976 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output200
timestamp 18001
transform 1 0 22264 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output201
timestamp 18001
transform 1 0 23552 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output202
timestamp 18001
transform -1 0 24564 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output203
timestamp 18001
transform 1 0 25576 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output204
timestamp 18001
transform -1 0 5520 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output205
timestamp 18001
transform -1 0 5520 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output206
timestamp 18001
transform -1 0 5520 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output207
timestamp 18001
transform -1 0 5520 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output208
timestamp 18001
transform -1 0 5520 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output209
timestamp 18001
transform -1 0 5520 0 -1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output210
timestamp 18001
transform -1 0 5520 0 -1 68000
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output211
timestamp 18001
transform -1 0 5520 0 -1 69088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output212
timestamp 18001
transform -1 0 5520 0 -1 70176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output213
timestamp 18001
transform -1 0 5520 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output214
timestamp 18001
transform -1 0 5520 0 1 70176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output215
timestamp 18001
transform -1 0 5520 0 -1 72352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output216
timestamp 18001
transform -1 0 5520 0 -1 73440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output217
timestamp 18001
transform -1 0 5520 0 -1 74528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output218
timestamp 18001
transform -1 0 5520 0 -1 75616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output219
timestamp 18001
transform -1 0 5520 0 1 75616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output220
timestamp 18001
transform -1 0 5520 0 -1 77792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output221
timestamp 18001
transform -1 0 5520 0 -1 78880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output222
timestamp 18001
transform -1 0 5520 0 -1 79968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output223
timestamp 18001
transform -1 0 5520 0 -1 81056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output224
timestamp 18001
transform -1 0 5520 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output225
timestamp 18001
transform -1 0 5520 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output226
timestamp 18001
transform -1 0 5520 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output227
timestamp 18001
transform -1 0 5520 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output228
timestamp 18001
transform -1 0 5520 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output229
timestamp 18001
transform -1 0 5520 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output230
timestamp 18001
transform -1 0 5520 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output231
timestamp 18001
transform -1 0 5520 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_155
timestamp 18001
transform 1 0 4876 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 18001
transform -1 0 88964 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_156
timestamp 18001
transform 1 0 4876 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 18001
transform -1 0 88964 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_157
timestamp 18001
transform 1 0 4876 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 18001
transform -1 0 88964 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_158
timestamp 18001
transform 1 0 4876 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 18001
transform -1 0 88964 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_159
timestamp 18001
transform 1 0 4876 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 18001
transform -1 0 88964 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_1_Left_309
timestamp 18001
transform 1 0 4876 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_1_Right_599
timestamp 18001
transform -1 0 7912 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_3_Left_310
timestamp 18001
transform 1 0 86020 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_3_Right_10
timestamp 18001
transform -1 0 88964 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_1_Left_160
timestamp 18001
transform 1 0 4876 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_1_Right_455
timestamp 18001
transform -1 0 7912 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_3_Left_311
timestamp 18001
transform 1 0 86020 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_3_Right_11
timestamp 18001
transform -1 0 88964 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_1_Left_161
timestamp 18001
transform 1 0 4876 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_1_Right_456
timestamp 18001
transform -1 0 7912 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_3_Left_312
timestamp 18001
transform 1 0 86020 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_3_Right_12
timestamp 18001
transform -1 0 88964 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_1_Left_162
timestamp 18001
transform 1 0 4876 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_1_Right_457
timestamp 18001
transform -1 0 7912 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_3_Left_313
timestamp 18001
transform 1 0 86020 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_3_Right_13
timestamp 18001
transform -1 0 88964 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_1_Left_163
timestamp 18001
transform 1 0 4876 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_1_Right_458
timestamp 18001
transform -1 0 7912 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_3_Left_314
timestamp 18001
transform 1 0 86020 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_3_Right_14
timestamp 18001
transform -1 0 88964 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_1_Left_164
timestamp 18001
transform 1 0 4876 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_1_Right_459
timestamp 18001
transform -1 0 7912 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_3_Left_315
timestamp 18001
transform 1 0 86020 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_3_Right_15
timestamp 18001
transform -1 0 88964 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_1_Left_165
timestamp 18001
transform 1 0 4876 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_1_Right_460
timestamp 18001
transform -1 0 7912 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_3_Left_316
timestamp 18001
transform 1 0 86020 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_3_Right_16
timestamp 18001
transform -1 0 88964 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_1_Left_166
timestamp 18001
transform 1 0 4876 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_1_Right_461
timestamp 18001
transform -1 0 7912 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_3_Left_317
timestamp 18001
transform 1 0 86020 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_3_Right_17
timestamp 18001
transform -1 0 88964 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_1_Left_167
timestamp 18001
transform 1 0 4876 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_1_Right_462
timestamp 18001
transform -1 0 7912 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_3_Left_318
timestamp 18001
transform 1 0 86020 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_3_Right_18
timestamp 18001
transform -1 0 88964 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_1_Left_168
timestamp 18001
transform 1 0 4876 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_1_Right_463
timestamp 18001
transform -1 0 7912 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_3_Left_319
timestamp 18001
transform 1 0 86020 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_3_Right_19
timestamp 18001
transform -1 0 88964 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_1_Left_169
timestamp 18001
transform 1 0 4876 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_1_Right_464
timestamp 18001
transform -1 0 7912 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_3_Left_320
timestamp 18001
transform 1 0 86020 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_3_Right_20
timestamp 18001
transform -1 0 88964 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_1_Left_170
timestamp 18001
transform 1 0 4876 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_1_Right_465
timestamp 18001
transform -1 0 7912 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_3_Left_321
timestamp 18001
transform 1 0 86020 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_3_Right_21
timestamp 18001
transform -1 0 88964 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_1_Left_171
timestamp 18001
transform 1 0 4876 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_1_Right_466
timestamp 18001
transform -1 0 7912 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_3_Left_322
timestamp 18001
transform 1 0 86020 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_3_Right_22
timestamp 18001
transform -1 0 88964 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_1_Left_172
timestamp 18001
transform 1 0 4876 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_1_Right_467
timestamp 18001
transform -1 0 7912 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_3_Left_323
timestamp 18001
transform 1 0 86020 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_3_Right_23
timestamp 18001
transform -1 0 88964 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_1_Left_173
timestamp 18001
transform 1 0 4876 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_1_Right_468
timestamp 18001
transform -1 0 7912 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_3_Left_324
timestamp 18001
transform 1 0 86020 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_3_Right_24
timestamp 18001
transform -1 0 88964 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_1_Left_174
timestamp 18001
transform 1 0 4876 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_1_Right_469
timestamp 18001
transform -1 0 7912 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_3_Left_325
timestamp 18001
transform 1 0 86020 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_3_Right_25
timestamp 18001
transform -1 0 88964 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_1_Left_175
timestamp 18001
transform 1 0 4876 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_1_Right_470
timestamp 18001
transform -1 0 7912 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_3_Left_326
timestamp 18001
transform 1 0 86020 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_3_Right_26
timestamp 18001
transform -1 0 88964 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_1_Left_176
timestamp 18001
transform 1 0 4876 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_1_Right_471
timestamp 18001
transform -1 0 7912 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_3_Left_327
timestamp 18001
transform 1 0 86020 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_3_Right_27
timestamp 18001
transform -1 0 88964 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_1_Left_177
timestamp 18001
transform 1 0 4876 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_1_Right_472
timestamp 18001
transform -1 0 7912 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_3_Left_328
timestamp 18001
transform 1 0 86020 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_3_Right_28
timestamp 18001
transform -1 0 88964 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_1_Left_178
timestamp 18001
transform 1 0 4876 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_1_Right_473
timestamp 18001
transform -1 0 7912 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_3_Left_329
timestamp 18001
transform 1 0 86020 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_3_Right_29
timestamp 18001
transform -1 0 88964 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_1_Left_179
timestamp 18001
transform 1 0 4876 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_1_Right_474
timestamp 18001
transform -1 0 7912 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_3_Left_330
timestamp 18001
transform 1 0 86020 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_3_Right_30
timestamp 18001
transform -1 0 88964 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_1_Left_180
timestamp 18001
transform 1 0 4876 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_1_Right_475
timestamp 18001
transform -1 0 7912 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_3_Left_331
timestamp 18001
transform 1 0 86020 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_3_Right_31
timestamp 18001
transform -1 0 88964 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_1_Left_181
timestamp 18001
transform 1 0 4876 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_1_Right_476
timestamp 18001
transform -1 0 7912 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_3_Left_332
timestamp 18001
transform 1 0 86020 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_3_Right_32
timestamp 18001
transform -1 0 88964 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_1_Left_182
timestamp 18001
transform 1 0 4876 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_1_Right_477
timestamp 18001
transform -1 0 7912 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_3_Left_333
timestamp 18001
transform 1 0 86020 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_3_Right_33
timestamp 18001
transform -1 0 88964 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_1_Left_183
timestamp 18001
transform 1 0 4876 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_1_Right_478
timestamp 18001
transform -1 0 7912 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_3_Left_334
timestamp 18001
transform 1 0 86020 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_3_Right_34
timestamp 18001
transform -1 0 88964 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_1_Left_184
timestamp 18001
transform 1 0 4876 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_1_Right_479
timestamp 18001
transform -1 0 7912 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_3_Left_335
timestamp 18001
transform 1 0 86020 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_3_Right_35
timestamp 18001
transform -1 0 88964 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_1_Left_185
timestamp 18001
transform 1 0 4876 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_1_Right_480
timestamp 18001
transform -1 0 7912 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_3_Left_336
timestamp 18001
transform 1 0 86020 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_3_Right_36
timestamp 18001
transform -1 0 88964 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_1_Left_186
timestamp 18001
transform 1 0 4876 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_1_Right_481
timestamp 18001
transform -1 0 7912 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_3_Left_337
timestamp 18001
transform 1 0 86020 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_3_Right_37
timestamp 18001
transform -1 0 88964 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_1_Left_187
timestamp 18001
transform 1 0 4876 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_1_Right_482
timestamp 18001
transform -1 0 7912 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_3_Left_338
timestamp 18001
transform 1 0 86020 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_3_Right_38
timestamp 18001
transform -1 0 88964 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_1_Left_188
timestamp 18001
transform 1 0 4876 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_1_Right_483
timestamp 18001
transform -1 0 7912 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_3_Left_339
timestamp 18001
transform 1 0 86020 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_3_Right_39
timestamp 18001
transform -1 0 88964 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_1_Left_189
timestamp 18001
transform 1 0 4876 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_1_Right_484
timestamp 18001
transform -1 0 7912 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_3_Left_340
timestamp 18001
transform 1 0 86020 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_3_Right_40
timestamp 18001
transform -1 0 88964 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_1_Left_190
timestamp 18001
transform 1 0 4876 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_1_Right_485
timestamp 18001
transform -1 0 7912 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_3_Left_341
timestamp 18001
transform 1 0 86020 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_3_Right_41
timestamp 18001
transform -1 0 88964 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_1_Left_191
timestamp 18001
transform 1 0 4876 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_1_Right_486
timestamp 18001
transform -1 0 7912 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_3_Left_342
timestamp 18001
transform 1 0 86020 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_3_Right_42
timestamp 18001
transform -1 0 88964 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_1_Left_192
timestamp 18001
transform 1 0 4876 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_1_Right_487
timestamp 18001
transform -1 0 7912 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_3_Left_343
timestamp 18001
transform 1 0 86020 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_3_Right_43
timestamp 18001
transform -1 0 88964 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_1_Left_193
timestamp 18001
transform 1 0 4876 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_1_Right_488
timestamp 18001
transform -1 0 7912 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_3_Left_344
timestamp 18001
transform 1 0 86020 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_3_Right_44
timestamp 18001
transform -1 0 88964 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_1_Left_194
timestamp 18001
transform 1 0 4876 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_1_Right_489
timestamp 18001
transform -1 0 7912 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_3_Left_345
timestamp 18001
transform 1 0 86020 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_3_Right_45
timestamp 18001
transform -1 0 88964 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_1_Left_195
timestamp 18001
transform 1 0 4876 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_1_Right_490
timestamp 18001
transform -1 0 7912 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_3_Left_346
timestamp 18001
transform 1 0 86020 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_3_Right_46
timestamp 18001
transform -1 0 88964 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_1_Left_196
timestamp 18001
transform 1 0 4876 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_1_Right_491
timestamp 18001
transform -1 0 7912 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_3_Left_347
timestamp 18001
transform 1 0 86020 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_3_Right_47
timestamp 18001
transform -1 0 88964 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_1_Left_197
timestamp 18001
transform 1 0 4876 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_1_Right_492
timestamp 18001
transform -1 0 7912 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_3_Left_348
timestamp 18001
transform 1 0 86020 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_3_Right_48
timestamp 18001
transform -1 0 88964 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_1_Left_198
timestamp 18001
transform 1 0 4876 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_1_Right_493
timestamp 18001
transform -1 0 7912 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_3_Left_349
timestamp 18001
transform 1 0 86020 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_3_Right_49
timestamp 18001
transform -1 0 88964 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_1_Left_199
timestamp 18001
transform 1 0 4876 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_1_Right_494
timestamp 18001
transform -1 0 7912 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_3_Left_350
timestamp 18001
transform 1 0 86020 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_3_Right_50
timestamp 18001
transform -1 0 88964 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_1_Left_200
timestamp 18001
transform 1 0 4876 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_1_Right_495
timestamp 18001
transform -1 0 7912 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_3_Left_351
timestamp 18001
transform 1 0 86020 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_3_Right_51
timestamp 18001
transform -1 0 88964 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_1_Left_201
timestamp 18001
transform 1 0 4876 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_1_Right_496
timestamp 18001
transform -1 0 7912 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_3_Left_352
timestamp 18001
transform 1 0 86020 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_3_Right_52
timestamp 18001
transform -1 0 88964 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_1_Left_202
timestamp 18001
transform 1 0 4876 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_1_Right_497
timestamp 18001
transform -1 0 7912 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_3_Left_353
timestamp 18001
transform 1 0 86020 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_3_Right_53
timestamp 18001
transform -1 0 88964 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_1_Left_203
timestamp 18001
transform 1 0 4876 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_1_Right_498
timestamp 18001
transform -1 0 7912 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_3_Left_354
timestamp 18001
transform 1 0 86020 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_3_Right_54
timestamp 18001
transform -1 0 88964 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_1_Left_204
timestamp 18001
transform 1 0 4876 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_1_Right_499
timestamp 18001
transform -1 0 7912 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_3_Left_355
timestamp 18001
transform 1 0 86020 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_3_Right_55
timestamp 18001
transform -1 0 88964 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_1_Left_205
timestamp 18001
transform 1 0 4876 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_1_Right_500
timestamp 18001
transform -1 0 7912 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_3_Left_356
timestamp 18001
transform 1 0 86020 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_3_Right_56
timestamp 18001
transform -1 0 88964 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_1_Left_206
timestamp 18001
transform 1 0 4876 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_1_Right_501
timestamp 18001
transform -1 0 7912 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_3_Left_357
timestamp 18001
transform 1 0 86020 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_3_Right_57
timestamp 18001
transform -1 0 88964 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_1_Left_207
timestamp 18001
transform 1 0 4876 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_1_Right_502
timestamp 18001
transform -1 0 7912 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_3_Left_358
timestamp 18001
transform 1 0 86020 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_3_Right_58
timestamp 18001
transform -1 0 88964 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_1_Left_208
timestamp 18001
transform 1 0 4876 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_1_Right_503
timestamp 18001
transform -1 0 7912 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_3_Left_359
timestamp 18001
transform 1 0 86020 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_3_Right_59
timestamp 18001
transform -1 0 88964 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_1_Left_209
timestamp 18001
transform 1 0 4876 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_1_Right_504
timestamp 18001
transform -1 0 7912 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_3_Left_360
timestamp 18001
transform 1 0 86020 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_3_Right_60
timestamp 18001
transform -1 0 88964 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_1_Left_210
timestamp 18001
transform 1 0 4876 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_1_Right_505
timestamp 18001
transform -1 0 7912 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_3_Left_361
timestamp 18001
transform 1 0 86020 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_3_Right_61
timestamp 18001
transform -1 0 88964 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_1_Left_211
timestamp 18001
transform 1 0 4876 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_1_Right_506
timestamp 18001
transform -1 0 7912 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_3_Left_362
timestamp 18001
transform 1 0 86020 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_3_Right_62
timestamp 18001
transform -1 0 88964 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_1_Left_212
timestamp 18001
transform 1 0 4876 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_1_Right_507
timestamp 18001
transform -1 0 7912 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_3_Left_363
timestamp 18001
transform 1 0 86020 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_3_Right_63
timestamp 18001
transform -1 0 88964 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_1_Left_213
timestamp 18001
transform 1 0 4876 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_1_Right_508
timestamp 18001
transform -1 0 7912 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_3_Left_364
timestamp 18001
transform 1 0 86020 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_3_Right_64
timestamp 18001
transform -1 0 88964 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_1_Left_214
timestamp 18001
transform 1 0 4876 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_1_Right_509
timestamp 18001
transform -1 0 7912 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_3_Left_365
timestamp 18001
transform 1 0 86020 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_3_Right_65
timestamp 18001
transform -1 0 88964 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_1_Left_215
timestamp 18001
transform 1 0 4876 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_1_Right_510
timestamp 18001
transform -1 0 7912 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_3_Left_366
timestamp 18001
transform 1 0 86020 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_3_Right_66
timestamp 18001
transform -1 0 88964 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_1_Left_216
timestamp 18001
transform 1 0 4876 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_1_Right_511
timestamp 18001
transform -1 0 7912 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_3_Left_367
timestamp 18001
transform 1 0 86020 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_3_Right_67
timestamp 18001
transform -1 0 88964 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_1_Left_217
timestamp 18001
transform 1 0 4876 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_1_Right_512
timestamp 18001
transform -1 0 7912 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_3_Left_368
timestamp 18001
transform 1 0 86020 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_3_Right_68
timestamp 18001
transform -1 0 88964 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_1_Left_218
timestamp 18001
transform 1 0 4876 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_1_Right_513
timestamp 18001
transform -1 0 7912 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_3_Left_369
timestamp 18001
transform 1 0 86020 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_3_Right_69
timestamp 18001
transform -1 0 88964 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_1_Left_219
timestamp 18001
transform 1 0 4876 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_1_Right_514
timestamp 18001
transform -1 0 7912 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_3_Left_370
timestamp 18001
transform 1 0 86020 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_3_Right_70
timestamp 18001
transform -1 0 88964 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_1_Left_220
timestamp 18001
transform 1 0 4876 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_1_Right_515
timestamp 18001
transform -1 0 7912 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_3_Left_371
timestamp 18001
transform 1 0 86020 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_3_Right_71
timestamp 18001
transform -1 0 88964 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_1_Left_221
timestamp 18001
transform 1 0 4876 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_1_Right_516
timestamp 18001
transform -1 0 7912 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_3_Left_372
timestamp 18001
transform 1 0 86020 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_3_Right_72
timestamp 18001
transform -1 0 88964 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_1_Left_222
timestamp 18001
transform 1 0 4876 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_1_Right_517
timestamp 18001
transform -1 0 7912 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_3_Left_373
timestamp 18001
transform 1 0 86020 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_3_Right_73
timestamp 18001
transform -1 0 88964 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_1_Left_223
timestamp 18001
transform 1 0 4876 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_1_Right_518
timestamp 18001
transform -1 0 7912 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_3_Left_374
timestamp 18001
transform 1 0 86020 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_3_Right_74
timestamp 18001
transform -1 0 88964 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_1_Left_224
timestamp 18001
transform 1 0 4876 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_1_Right_519
timestamp 18001
transform -1 0 7912 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_3_Left_375
timestamp 18001
transform 1 0 86020 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_3_Right_75
timestamp 18001
transform -1 0 88964 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_1_Left_225
timestamp 18001
transform 1 0 4876 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_1_Right_520
timestamp 18001
transform -1 0 7912 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_3_Left_376
timestamp 18001
transform 1 0 86020 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_3_Right_76
timestamp 18001
transform -1 0 88964 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_1_Left_226
timestamp 18001
transform 1 0 4876 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_1_Right_521
timestamp 18001
transform -1 0 7912 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_3_Left_377
timestamp 18001
transform 1 0 86020 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_3_Right_77
timestamp 18001
transform -1 0 88964 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_1_Left_227
timestamp 18001
transform 1 0 4876 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_1_Right_522
timestamp 18001
transform -1 0 7912 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_3_Left_378
timestamp 18001
transform 1 0 86020 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_3_Right_78
timestamp 18001
transform -1 0 88964 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_1_Left_228
timestamp 18001
transform 1 0 4876 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_1_Right_523
timestamp 18001
transform -1 0 7912 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_5_Left_379
timestamp 18001
transform 1 0 86020 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_5_Right_79
timestamp 18001
transform -1 0 88964 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_1_Left_229
timestamp 18001
transform 1 0 4876 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_1_Right_524
timestamp 18001
transform -1 0 7912 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_5_Left_380
timestamp 18001
transform 1 0 86020 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_5_Right_80
timestamp 18001
transform -1 0 88964 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_1_Left_230
timestamp 18001
transform 1 0 4876 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_1_Right_525
timestamp 18001
transform -1 0 7912 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_5_Left_381
timestamp 18001
transform 1 0 86020 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_5_Right_81
timestamp 18001
transform -1 0 88964 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_1_Left_231
timestamp 18001
transform 1 0 4876 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_1_Right_526
timestamp 18001
transform -1 0 7912 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_5_Left_382
timestamp 18001
transform 1 0 86020 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_5_Right_82
timestamp 18001
transform -1 0 88964 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_1_Left_232
timestamp 18001
transform 1 0 4876 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_1_Right_527
timestamp 18001
transform -1 0 7912 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_5_Left_383
timestamp 18001
transform 1 0 86020 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_78_5_Right_83
timestamp 18001
transform -1 0 88964 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_1_Left_233
timestamp 18001
transform 1 0 4876 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_1_Right_528
timestamp 18001
transform -1 0 7912 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_5_Left_384
timestamp 18001
transform 1 0 86020 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_79_5_Right_84
timestamp 18001
transform -1 0 88964 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_1_Left_234
timestamp 18001
transform 1 0 4876 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_1_Right_529
timestamp 18001
transform -1 0 7912 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_5_Left_385
timestamp 18001
transform 1 0 86020 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_80_5_Right_85
timestamp 18001
transform -1 0 88964 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_1_Left_235
timestamp 18001
transform 1 0 4876 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_1_Right_530
timestamp 18001
transform -1 0 7912 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_5_Left_386
timestamp 18001
transform 1 0 86020 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_81_5_Right_86
timestamp 18001
transform -1 0 88964 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_1_Left_236
timestamp 18001
transform 1 0 4876 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_1_Right_531
timestamp 18001
transform -1 0 7912 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_3_Left_387
timestamp 18001
transform 1 0 86020 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_82_3_Right_87
timestamp 18001
transform -1 0 88964 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_1_Left_237
timestamp 18001
transform 1 0 4876 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_1_Right_532
timestamp 18001
transform -1 0 7912 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_3_Left_388
timestamp 18001
transform 1 0 86020 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_83_3_Right_88
timestamp 18001
transform -1 0 88964 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_1_Left_238
timestamp 18001
transform 1 0 4876 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_1_Right_533
timestamp 18001
transform -1 0 7912 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_3_Left_389
timestamp 18001
transform 1 0 86020 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_84_3_Right_89
timestamp 18001
transform -1 0 88964 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_1_Left_239
timestamp 18001
transform 1 0 4876 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_1_Right_534
timestamp 18001
transform -1 0 7912 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_3_Left_390
timestamp 18001
transform 1 0 86020 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_85_3_Right_90
timestamp 18001
transform -1 0 88964 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_1_Left_240
timestamp 18001
transform 1 0 4876 0 1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_1_Right_535
timestamp 18001
transform -1 0 7912 0 1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_3_Left_391
timestamp 18001
transform 1 0 86020 0 1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_86_3_Right_91
timestamp 18001
transform -1 0 88964 0 1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_1_Left_241
timestamp 18001
transform 1 0 4876 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_1_Right_536
timestamp 18001
transform -1 0 7912 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_3_Left_392
timestamp 18001
transform 1 0 86020 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_87_3_Right_92
timestamp 18001
transform -1 0 88964 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_1_Left_242
timestamp 18001
transform 1 0 4876 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_1_Right_537
timestamp 18001
transform -1 0 7912 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_3_Left_393
timestamp 18001
transform 1 0 86020 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_88_3_Right_93
timestamp 18001
transform -1 0 88964 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_1_Left_243
timestamp 18001
transform 1 0 4876 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_1_Right_538
timestamp 18001
transform -1 0 7912 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_3_Left_394
timestamp 18001
transform 1 0 86020 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_89_3_Right_94
timestamp 18001
transform -1 0 88964 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_1_Left_244
timestamp 18001
transform 1 0 4876 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_1_Right_539
timestamp 18001
transform -1 0 7912 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_3_Left_395
timestamp 18001
transform 1 0 86020 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_90_3_Right_95
timestamp 18001
transform -1 0 88964 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_1_Left_245
timestamp 18001
transform 1 0 4876 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_1_Right_540
timestamp 18001
transform -1 0 7912 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_3_Left_396
timestamp 18001
transform 1 0 86020 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_91_3_Right_96
timestamp 18001
transform -1 0 88964 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_1_Left_246
timestamp 18001
transform 1 0 4876 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_1_Right_541
timestamp 18001
transform -1 0 7912 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_3_Left_397
timestamp 18001
transform 1 0 86020 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_92_3_Right_97
timestamp 18001
transform -1 0 88964 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_1_Left_247
timestamp 18001
transform 1 0 4876 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_1_Right_542
timestamp 18001
transform -1 0 7912 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_3_Left_398
timestamp 18001
transform 1 0 86020 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_93_3_Right_98
timestamp 18001
transform -1 0 88964 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_1_Left_248
timestamp 18001
transform 1 0 4876 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_1_Right_543
timestamp 18001
transform -1 0 7912 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_3_Left_399
timestamp 18001
transform 1 0 86020 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_94_3_Right_99
timestamp 18001
transform -1 0 88964 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_1_Left_249
timestamp 18001
transform 1 0 4876 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_1_Right_544
timestamp 18001
transform -1 0 7912 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_3_Left_400
timestamp 18001
transform 1 0 86020 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_95_3_Right_100
timestamp 18001
transform -1 0 88964 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_1_Left_250
timestamp 18001
transform 1 0 4876 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_1_Right_545
timestamp 18001
transform -1 0 7912 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_3_Left_401
timestamp 18001
transform 1 0 86020 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_96_3_Right_101
timestamp 18001
transform -1 0 88964 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_1_Left_251
timestamp 18001
transform 1 0 4876 0 -1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_1_Right_546
timestamp 18001
transform -1 0 7912 0 -1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_3_Left_402
timestamp 18001
transform 1 0 86020 0 -1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_97_3_Right_102
timestamp 18001
transform -1 0 88964 0 -1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_1_Left_252
timestamp 18001
transform 1 0 4876 0 1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_1_Right_547
timestamp 18001
transform -1 0 7912 0 1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_3_Left_403
timestamp 18001
transform 1 0 86020 0 1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_98_3_Right_103
timestamp 18001
transform -1 0 88964 0 1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_1_Left_253
timestamp 18001
transform 1 0 4876 0 -1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_1_Right_548
timestamp 18001
transform -1 0 7912 0 -1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_3_Left_404
timestamp 18001
transform 1 0 86020 0 -1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_99_3_Right_104
timestamp 18001
transform -1 0 88964 0 -1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_1_Left_254
timestamp 18001
transform 1 0 4876 0 1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_1_Right_549
timestamp 18001
transform -1 0 7912 0 1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_3_Left_405
timestamp 18001
transform 1 0 86020 0 1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_100_3_Right_105
timestamp 18001
transform -1 0 88964 0 1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_1_Left_255
timestamp 18001
transform 1 0 4876 0 -1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_1_Right_550
timestamp 18001
transform -1 0 7912 0 -1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_3_Left_406
timestamp 18001
transform 1 0 86020 0 -1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_101_3_Right_106
timestamp 18001
transform -1 0 88964 0 -1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_1_Left_256
timestamp 18001
transform 1 0 4876 0 1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_1_Right_551
timestamp 18001
transform -1 0 7912 0 1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_3_Left_407
timestamp 18001
transform 1 0 86020 0 1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_102_3_Right_107
timestamp 18001
transform -1 0 88964 0 1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_1_Left_257
timestamp 18001
transform 1 0 4876 0 -1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_1_Right_552
timestamp 18001
transform -1 0 7912 0 -1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_3_Left_408
timestamp 18001
transform 1 0 86020 0 -1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_103_3_Right_108
timestamp 18001
transform -1 0 88964 0 -1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_1_Left_258
timestamp 18001
transform 1 0 4876 0 1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_1_Right_553
timestamp 18001
transform -1 0 7912 0 1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_3_Left_409
timestamp 18001
transform 1 0 86020 0 1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_104_3_Right_109
timestamp 18001
transform -1 0 88964 0 1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_1_Left_259
timestamp 18001
transform 1 0 4876 0 -1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_1_Right_554
timestamp 18001
transform -1 0 7912 0 -1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_3_Left_410
timestamp 18001
transform 1 0 86020 0 -1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_105_3_Right_110
timestamp 18001
transform -1 0 88964 0 -1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_1_Left_260
timestamp 18001
transform 1 0 4876 0 1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_1_Right_555
timestamp 18001
transform -1 0 7912 0 1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_3_Left_411
timestamp 18001
transform 1 0 86020 0 1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_106_3_Right_111
timestamp 18001
transform -1 0 88964 0 1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_1_Left_261
timestamp 18001
transform 1 0 4876 0 -1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_1_Right_556
timestamp 18001
transform -1 0 7912 0 -1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_3_Left_412
timestamp 18001
transform 1 0 86020 0 -1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_107_3_Right_112
timestamp 18001
transform -1 0 88964 0 -1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_1_Left_262
timestamp 18001
transform 1 0 4876 0 1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_1_Right_557
timestamp 18001
transform -1 0 7912 0 1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_3_Left_413
timestamp 18001
transform 1 0 86020 0 1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_108_3_Right_113
timestamp 18001
transform -1 0 88964 0 1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_1_Left_263
timestamp 18001
transform 1 0 4876 0 -1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_1_Right_558
timestamp 18001
transform -1 0 7912 0 -1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_3_Left_414
timestamp 18001
transform 1 0 86020 0 -1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_109_3_Right_114
timestamp 18001
transform -1 0 88964 0 -1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_1_Left_264
timestamp 18001
transform 1 0 4876 0 1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_1_Right_559
timestamp 18001
transform -1 0 7912 0 1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_3_Left_415
timestamp 18001
transform 1 0 86020 0 1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_110_3_Right_115
timestamp 18001
transform -1 0 88964 0 1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_1_Left_265
timestamp 18001
transform 1 0 4876 0 -1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_1_Right_560
timestamp 18001
transform -1 0 7912 0 -1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_3_Left_416
timestamp 18001
transform 1 0 86020 0 -1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_111_3_Right_116
timestamp 18001
transform -1 0 88964 0 -1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_1_Left_266
timestamp 18001
transform 1 0 4876 0 1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_1_Right_561
timestamp 18001
transform -1 0 7912 0 1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_3_Left_417
timestamp 18001
transform 1 0 86020 0 1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_112_3_Right_117
timestamp 18001
transform -1 0 88964 0 1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_1_Left_267
timestamp 18001
transform 1 0 4876 0 -1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_1_Right_562
timestamp 18001
transform -1 0 7912 0 -1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_3_Left_418
timestamp 18001
transform 1 0 86020 0 -1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_113_3_Right_118
timestamp 18001
transform -1 0 88964 0 -1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_1_Left_268
timestamp 18001
transform 1 0 4876 0 1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_1_Right_563
timestamp 18001
transform -1 0 7912 0 1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_3_Left_419
timestamp 18001
transform 1 0 86020 0 1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_114_3_Right_119
timestamp 18001
transform -1 0 88964 0 1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_1_Left_269
timestamp 18001
transform 1 0 4876 0 -1 68000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_1_Right_564
timestamp 18001
transform -1 0 7912 0 -1 68000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_3_Left_420
timestamp 18001
transform 1 0 86020 0 -1 68000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_115_3_Right_120
timestamp 18001
transform -1 0 88964 0 -1 68000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_1_Left_270
timestamp 18001
transform 1 0 4876 0 1 68000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_1_Right_565
timestamp 18001
transform -1 0 7912 0 1 68000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_3_Left_421
timestamp 18001
transform 1 0 86020 0 1 68000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_116_3_Right_121
timestamp 18001
transform -1 0 88964 0 1 68000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_117_1_Left_271
timestamp 18001
transform 1 0 4876 0 -1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_117_1_Right_566
timestamp 18001
transform -1 0 7912 0 -1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_117_3_Left_422
timestamp 18001
transform 1 0 86020 0 -1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_117_3_Right_122
timestamp 18001
transform -1 0 88964 0 -1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_118_1_Left_272
timestamp 18001
transform 1 0 4876 0 1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_118_1_Right_567
timestamp 18001
transform -1 0 7912 0 1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_118_3_Left_423
timestamp 18001
transform 1 0 86020 0 1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_118_3_Right_123
timestamp 18001
transform -1 0 88964 0 1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_119_1_Left_273
timestamp 18001
transform 1 0 4876 0 -1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_119_1_Right_568
timestamp 18001
transform -1 0 7912 0 -1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_119_3_Left_424
timestamp 18001
transform 1 0 86020 0 -1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_119_3_Right_124
timestamp 18001
transform -1 0 88964 0 -1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_120_1_Left_274
timestamp 18001
transform 1 0 4876 0 1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_120_1_Right_569
timestamp 18001
transform -1 0 7912 0 1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_120_3_Left_425
timestamp 18001
transform 1 0 86020 0 1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_120_3_Right_125
timestamp 18001
transform -1 0 88964 0 1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_121_1_Left_275
timestamp 18001
transform 1 0 4876 0 -1 71264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_121_1_Right_570
timestamp 18001
transform -1 0 7912 0 -1 71264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_121_3_Left_426
timestamp 18001
transform 1 0 86020 0 -1 71264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_121_3_Right_126
timestamp 18001
transform -1 0 88964 0 -1 71264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_122_1_Left_276
timestamp 18001
transform 1 0 4876 0 1 71264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_122_1_Right_571
timestamp 18001
transform -1 0 7912 0 1 71264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_122_3_Left_427
timestamp 18001
transform 1 0 86020 0 1 71264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_122_3_Right_127
timestamp 18001
transform -1 0 88964 0 1 71264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_123_1_Left_277
timestamp 18001
transform 1 0 4876 0 -1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_123_1_Right_572
timestamp 18001
transform -1 0 7912 0 -1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_123_3_Left_428
timestamp 18001
transform 1 0 86020 0 -1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_123_3_Right_128
timestamp 18001
transform -1 0 88964 0 -1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_124_1_Left_278
timestamp 18001
transform 1 0 4876 0 1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_124_1_Right_573
timestamp 18001
transform -1 0 7912 0 1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_124_3_Left_429
timestamp 18001
transform 1 0 86020 0 1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_124_3_Right_129
timestamp 18001
transform -1 0 88964 0 1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_125_1_Left_279
timestamp 18001
transform 1 0 4876 0 -1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_125_1_Right_574
timestamp 18001
transform -1 0 7912 0 -1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_125_3_Left_430
timestamp 18001
transform 1 0 86020 0 -1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_125_3_Right_130
timestamp 18001
transform -1 0 88964 0 -1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_126_1_Left_280
timestamp 18001
transform 1 0 4876 0 1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_126_1_Right_575
timestamp 18001
transform -1 0 7912 0 1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_126_3_Left_431
timestamp 18001
transform 1 0 86020 0 1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_126_3_Right_131
timestamp 18001
transform -1 0 88964 0 1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_127_1_Left_281
timestamp 18001
transform 1 0 4876 0 -1 74528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_127_1_Right_576
timestamp 18001
transform -1 0 7912 0 -1 74528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_127_3_Left_432
timestamp 18001
transform 1 0 86020 0 -1 74528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_127_3_Right_132
timestamp 18001
transform -1 0 88964 0 -1 74528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_128_1_Left_282
timestamp 18001
transform 1 0 4876 0 1 74528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_128_1_Right_577
timestamp 18001
transform -1 0 7912 0 1 74528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_128_3_Left_433
timestamp 18001
transform 1 0 86020 0 1 74528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_128_3_Right_133
timestamp 18001
transform -1 0 88964 0 1 74528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_129_1_Left_283
timestamp 18001
transform 1 0 4876 0 -1 75616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_129_1_Right_578
timestamp 18001
transform -1 0 7912 0 -1 75616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_129_3_Left_434
timestamp 18001
transform 1 0 86020 0 -1 75616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_129_3_Right_134
timestamp 18001
transform -1 0 88964 0 -1 75616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_130_1_Left_284
timestamp 18001
transform 1 0 4876 0 1 75616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_130_1_Right_579
timestamp 18001
transform -1 0 7912 0 1 75616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_130_3_Left_435
timestamp 18001
transform 1 0 86020 0 1 75616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_130_3_Right_135
timestamp 18001
transform -1 0 88964 0 1 75616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_131_1_Left_285
timestamp 18001
transform 1 0 4876 0 -1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_131_1_Right_580
timestamp 18001
transform -1 0 7912 0 -1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_131_3_Left_436
timestamp 18001
transform 1 0 86020 0 -1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_131_3_Right_136
timestamp 18001
transform -1 0 88964 0 -1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_132_1_Left_286
timestamp 18001
transform 1 0 4876 0 1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_132_1_Right_581
timestamp 18001
transform -1 0 7912 0 1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_132_3_Left_437
timestamp 18001
transform 1 0 86020 0 1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_132_3_Right_137
timestamp 18001
transform -1 0 88964 0 1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_133_1_Left_287
timestamp 18001
transform 1 0 4876 0 -1 77792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_133_1_Right_582
timestamp 18001
transform -1 0 7912 0 -1 77792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_133_3_Left_438
timestamp 18001
transform 1 0 86020 0 -1 77792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_133_3_Right_138
timestamp 18001
transform -1 0 88964 0 -1 77792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_134_1_Left_288
timestamp 18001
transform 1 0 4876 0 1 77792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_134_1_Right_583
timestamp 18001
transform -1 0 7912 0 1 77792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_134_3_Left_439
timestamp 18001
transform 1 0 86020 0 1 77792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_134_3_Right_139
timestamp 18001
transform -1 0 88964 0 1 77792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_135_1_Left_289
timestamp 18001
transform 1 0 4876 0 -1 78880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_135_1_Right_584
timestamp 18001
transform -1 0 7912 0 -1 78880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_135_3_Left_440
timestamp 18001
transform 1 0 86020 0 -1 78880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_135_3_Right_140
timestamp 18001
transform -1 0 88964 0 -1 78880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_136_1_Left_290
timestamp 18001
transform 1 0 4876 0 1 78880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_136_1_Right_585
timestamp 18001
transform -1 0 7912 0 1 78880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_136_3_Left_441
timestamp 18001
transform 1 0 86020 0 1 78880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_136_3_Right_141
timestamp 18001
transform -1 0 88964 0 1 78880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_137_1_Left_291
timestamp 18001
transform 1 0 4876 0 -1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_137_1_Right_586
timestamp 18001
transform -1 0 7912 0 -1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_137_3_Left_442
timestamp 18001
transform 1 0 86020 0 -1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_137_3_Right_142
timestamp 18001
transform -1 0 88964 0 -1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_138_1_Left_292
timestamp 18001
transform 1 0 4876 0 1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_138_1_Right_587
timestamp 18001
transform -1 0 7912 0 1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_138_3_Left_443
timestamp 18001
transform 1 0 86020 0 1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_138_3_Right_143
timestamp 18001
transform -1 0 88964 0 1 79968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_139_1_Left_293
timestamp 18001
transform 1 0 4876 0 -1 81056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_139_1_Right_588
timestamp 18001
transform -1 0 7912 0 -1 81056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_139_3_Left_444
timestamp 18001
transform 1 0 86020 0 -1 81056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_139_3_Right_144
timestamp 18001
transform -1 0 88964 0 -1 81056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_140_1_Left_294
timestamp 18001
transform 1 0 4876 0 1 81056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_140_1_Right_589
timestamp 18001
transform -1 0 7912 0 1 81056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_140_3_Left_445
timestamp 18001
transform 1 0 86020 0 1 81056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_140_3_Right_145
timestamp 18001
transform -1 0 88964 0 1 81056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_141_1_Left_295
timestamp 18001
transform 1 0 4876 0 -1 82144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_141_1_Right_590
timestamp 18001
transform -1 0 7912 0 -1 82144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_141_3_Left_446
timestamp 18001
transform 1 0 86020 0 -1 82144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_141_3_Right_146
timestamp 18001
transform -1 0 88964 0 -1 82144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_142_1_Left_296
timestamp 18001
transform 1 0 4876 0 1 82144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_142_1_Right_591
timestamp 18001
transform -1 0 7912 0 1 82144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_142_3_Left_447
timestamp 18001
transform 1 0 86020 0 1 82144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_142_3_Right_147
timestamp 18001
transform -1 0 88964 0 1 82144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_143_1_Left_297
timestamp 18001
transform 1 0 4876 0 -1 83232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_143_1_Right_592
timestamp 18001
transform -1 0 7912 0 -1 83232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_143_3_Left_448
timestamp 18001
transform 1 0 86020 0 -1 83232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_143_3_Right_148
timestamp 18001
transform -1 0 88964 0 -1 83232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_144_1_Left_298
timestamp 18001
transform 1 0 4876 0 1 83232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_144_1_Right_593
timestamp 18001
transform -1 0 7912 0 1 83232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_144_3_Left_449
timestamp 18001
transform 1 0 86020 0 1 83232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_144_3_Right_149
timestamp 18001
transform -1 0 88964 0 1 83232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_145_1_Left_299
timestamp 18001
transform 1 0 4876 0 -1 84320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_145_1_Right_594
timestamp 18001
transform -1 0 7912 0 -1 84320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_145_3_Left_450
timestamp 18001
transform 1 0 86020 0 -1 84320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_145_3_Right_150
timestamp 18001
transform -1 0 88964 0 -1 84320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_146_1_Left_300
timestamp 18001
transform 1 0 4876 0 1 84320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_146_1_Right_595
timestamp 18001
transform -1 0 7912 0 1 84320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_146_3_Left_451
timestamp 18001
transform 1 0 86020 0 1 84320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_146_3_Right_151
timestamp 18001
transform -1 0 88964 0 1 84320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_147_1_Left_301
timestamp 18001
transform 1 0 4876 0 -1 85408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_147_1_Right_596
timestamp 18001
transform -1 0 7912 0 -1 85408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_147_3_Left_452
timestamp 18001
transform 1 0 86020 0 -1 85408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_147_3_Right_152
timestamp 18001
transform -1 0 88964 0 -1 85408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_148_1_Left_302
timestamp 18001
transform 1 0 4876 0 1 85408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_148_1_Right_597
timestamp 18001
transform -1 0 7912 0 1 85408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_148_3_Left_453
timestamp 18001
transform 1 0 86020 0 1 85408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_148_3_Right_153
timestamp 18001
transform -1 0 88964 0 1 85408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_149_1_Left_303
timestamp 18001
transform 1 0 4876 0 -1 86496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_149_1_Right_598
timestamp 18001
transform -1 0 7912 0 -1 86496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_149_3_Left_454
timestamp 18001
transform 1 0 86020 0 -1 86496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_149_3_Right_154
timestamp 18001
transform -1 0 88964 0 -1 86496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_150_Left_304
timestamp 18001
transform 1 0 4876 0 1 86496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_150_Right_5
timestamp 18001
transform -1 0 88964 0 1 86496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_151_Left_305
timestamp 18001
transform 1 0 4876 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_151_Right_6
timestamp 18001
transform -1 0 88964 0 -1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_152_Left_306
timestamp 18001
transform 1 0 4876 0 1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_152_Right_7
timestamp 18001
transform -1 0 88964 0 1 87584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_153_Left_307
timestamp 18001
transform 1 0 4876 0 -1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_153_Right_8
timestamp 18001
transform -1 0 88964 0 -1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_154_Left_308
timestamp 18001
transform 1 0 4876 0 1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_154_Right_9
timestamp 18001
transform -1 0 88964 0 1 88672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_600
timestamp 18001
transform 1 0 7452 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_601
timestamp 18001
transform 1 0 10028 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_602
timestamp 18001
transform 1 0 12604 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_603
timestamp 18001
transform 1 0 15180 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_604
timestamp 18001
transform 1 0 17756 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_605
timestamp 18001
transform 1 0 20332 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_606
timestamp 18001
transform 1 0 22908 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_607
timestamp 18001
transform 1 0 25484 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_608
timestamp 18001
transform 1 0 28060 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_609
timestamp 18001
transform 1 0 30636 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_610
timestamp 18001
transform 1 0 33212 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_611
timestamp 18001
transform 1 0 35788 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_612
timestamp 18001
transform 1 0 38364 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_613
timestamp 18001
transform 1 0 40940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_614
timestamp 18001
transform 1 0 43516 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_615
timestamp 18001
transform 1 0 46092 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_616
timestamp 18001
transform 1 0 48668 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_617
timestamp 18001
transform 1 0 51244 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_618
timestamp 18001
transform 1 0 53820 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_619
timestamp 18001
transform 1 0 56396 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_620
timestamp 18001
transform 1 0 58972 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_621
timestamp 18001
transform 1 0 61548 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_622
timestamp 18001
transform 1 0 64124 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_623
timestamp 18001
transform 1 0 66700 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_624
timestamp 18001
transform 1 0 69276 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_625
timestamp 18001
transform 1 0 71852 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_626
timestamp 18001
transform 1 0 74428 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_627
timestamp 18001
transform 1 0 77004 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_628
timestamp 18001
transform 1 0 79580 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_629
timestamp 18001
transform 1 0 82156 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_630
timestamp 18001
transform 1 0 84732 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_631
timestamp 18001
transform 1 0 87308 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_632
timestamp 18001
transform 1 0 10028 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_633
timestamp 18001
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_634
timestamp 18001
transform 1 0 20332 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_635
timestamp 18001
transform 1 0 25484 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_636
timestamp 18001
transform 1 0 30636 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_637
timestamp 18001
transform 1 0 35788 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_638
timestamp 18001
transform 1 0 40940 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_639
timestamp 18001
transform 1 0 46092 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_640
timestamp 18001
transform 1 0 51244 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_641
timestamp 18001
transform 1 0 56396 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_642
timestamp 18001
transform 1 0 61548 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_643
timestamp 18001
transform 1 0 66700 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_644
timestamp 18001
transform 1 0 71852 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_645
timestamp 18001
transform 1 0 77004 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_646
timestamp 18001
transform 1 0 82156 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_647
timestamp 18001
transform 1 0 87308 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_648
timestamp 18001
transform 1 0 7452 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_649
timestamp 18001
transform 1 0 12604 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_650
timestamp 18001
transform 1 0 17756 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_651
timestamp 18001
transform 1 0 22908 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_652
timestamp 18001
transform 1 0 28060 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_653
timestamp 18001
transform 1 0 33212 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_654
timestamp 18001
transform 1 0 38364 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_655
timestamp 18001
transform 1 0 43516 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_656
timestamp 18001
transform 1 0 48668 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_657
timestamp 18001
transform 1 0 53820 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_658
timestamp 18001
transform 1 0 58972 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_659
timestamp 18001
transform 1 0 64124 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_660
timestamp 18001
transform 1 0 69276 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_661
timestamp 18001
transform 1 0 74428 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_662
timestamp 18001
transform 1 0 79580 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_663
timestamp 18001
transform 1 0 84732 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_664
timestamp 18001
transform 1 0 10028 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_665
timestamp 18001
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_666
timestamp 18001
transform 1 0 20332 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_667
timestamp 18001
transform 1 0 25484 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_668
timestamp 18001
transform 1 0 30636 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_669
timestamp 18001
transform 1 0 35788 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_670
timestamp 18001
transform 1 0 40940 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_671
timestamp 18001
transform 1 0 46092 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_672
timestamp 18001
transform 1 0 51244 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_673
timestamp 18001
transform 1 0 56396 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_674
timestamp 18001
transform 1 0 61548 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_675
timestamp 18001
transform 1 0 66700 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_676
timestamp 18001
transform 1 0 71852 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_677
timestamp 18001
transform 1 0 77004 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_678
timestamp 18001
transform 1 0 82156 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_679
timestamp 18001
transform 1 0 87308 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_680
timestamp 18001
transform 1 0 7452 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_681
timestamp 18001
transform 1 0 10028 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_682
timestamp 18001
transform 1 0 12604 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_683
timestamp 18001
transform 1 0 15180 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_684
timestamp 18001
transform 1 0 17756 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_685
timestamp 18001
transform 1 0 20332 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_686
timestamp 18001
transform 1 0 22908 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_687
timestamp 18001
transform 1 0 25484 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_688
timestamp 18001
transform 1 0 28060 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_689
timestamp 18001
transform 1 0 30636 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_690
timestamp 18001
transform 1 0 33212 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_691
timestamp 18001
transform 1 0 35788 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_692
timestamp 18001
transform 1 0 38364 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_693
timestamp 18001
transform 1 0 40940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_694
timestamp 18001
transform 1 0 43516 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_695
timestamp 18001
transform 1 0 46092 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_696
timestamp 18001
transform 1 0 48668 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_697
timestamp 18001
transform 1 0 51244 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_698
timestamp 18001
transform 1 0 53820 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_699
timestamp 18001
transform 1 0 56396 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_700
timestamp 18001
transform 1 0 58972 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_701
timestamp 18001
transform 1 0 61548 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_702
timestamp 18001
transform 1 0 64124 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_703
timestamp 18001
transform 1 0 66700 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_704
timestamp 18001
transform 1 0 69276 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_705
timestamp 18001
transform 1 0 71852 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_706
timestamp 18001
transform 1 0 74428 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_707
timestamp 18001
transform 1 0 77004 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_708
timestamp 18001
transform 1 0 79580 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_709
timestamp 18001
transform 1 0 82156 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_710
timestamp 18001
transform 1 0 84732 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_711
timestamp 18001
transform 1 0 87308 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1_712
timestamp 18001
transform 1 0 7452 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_3_896
timestamp 18001
transform 1 0 88596 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1_713
timestamp 18001
transform 1 0 7452 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_3_897
timestamp 18001
transform 1 0 88596 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_1_714
timestamp 18001
transform 1 0 7452 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_3_898
timestamp 18001
transform 1 0 88596 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_1_715
timestamp 18001
transform 1 0 7452 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_3_899
timestamp 18001
transform 1 0 88596 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_1_716
timestamp 18001
transform 1 0 7452 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_3_900
timestamp 18001
transform 1 0 88596 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_1_717
timestamp 18001
transform 1 0 7452 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_3_901
timestamp 18001
transform 1 0 88596 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_1_718
timestamp 18001
transform 1 0 7452 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_3_902
timestamp 18001
transform 1 0 88596 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_1_719
timestamp 18001
transform 1 0 7452 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_3_903
timestamp 18001
transform 1 0 88596 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_1_720
timestamp 18001
transform 1 0 7452 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_3_904
timestamp 18001
transform 1 0 88596 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_1_721
timestamp 18001
transform 1 0 7452 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_3_905
timestamp 18001
transform 1 0 88596 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_1_722
timestamp 18001
transform 1 0 7452 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_3_906
timestamp 18001
transform 1 0 88596 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_1_723
timestamp 18001
transform 1 0 7452 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_3_907
timestamp 18001
transform 1 0 88596 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_1_724
timestamp 18001
transform 1 0 7452 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_3_908
timestamp 18001
transform 1 0 88596 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_1_725
timestamp 18001
transform 1 0 7452 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_3_909
timestamp 18001
transform 1 0 88596 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_1_726
timestamp 18001
transform 1 0 7452 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_3_910
timestamp 18001
transform 1 0 88596 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_1_727
timestamp 18001
transform 1 0 7452 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_3_911
timestamp 18001
transform 1 0 88596 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_1_728
timestamp 18001
transform 1 0 7452 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_3_912
timestamp 18001
transform 1 0 88596 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_1_729
timestamp 18001
transform 1 0 7452 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_3_913
timestamp 18001
transform 1 0 88596 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_1_730
timestamp 18001
transform 1 0 7452 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_3_914
timestamp 18001
transform 1 0 88596 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_1_731
timestamp 18001
transform 1 0 7452 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_3_915
timestamp 18001
transform 1 0 88596 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_1_732
timestamp 18001
transform 1 0 7452 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_3_916
timestamp 18001
transform 1 0 88596 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_1_733
timestamp 18001
transform 1 0 7452 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_3_917
timestamp 18001
transform 1 0 88596 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_1_734
timestamp 18001
transform 1 0 7452 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_3_918
timestamp 18001
transform 1 0 88596 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_1_735
timestamp 18001
transform 1 0 7452 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_3_919
timestamp 18001
transform 1 0 88596 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_1_736
timestamp 18001
transform 1 0 7452 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_3_920
timestamp 18001
transform 1 0 88596 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_1_737
timestamp 18001
transform 1 0 7452 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_3_921
timestamp 18001
transform 1 0 88596 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_1_738
timestamp 18001
transform 1 0 7452 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_3_922
timestamp 18001
transform 1 0 88596 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_1_739
timestamp 18001
transform 1 0 7452 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_3_923
timestamp 18001
transform 1 0 88596 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_1_740
timestamp 18001
transform 1 0 7452 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_3_924
timestamp 18001
transform 1 0 88596 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_1_741
timestamp 18001
transform 1 0 7452 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_3_925
timestamp 18001
transform 1 0 88596 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_1_742
timestamp 18001
transform 1 0 7452 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_3_926
timestamp 18001
transform 1 0 88596 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_1_743
timestamp 18001
transform 1 0 7452 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_3_927
timestamp 18001
transform 1 0 88596 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_1_744
timestamp 18001
transform 1 0 7452 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_3_928
timestamp 18001
transform 1 0 88596 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_1_745
timestamp 18001
transform 1 0 7452 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_3_929
timestamp 18001
transform 1 0 88596 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_1_746
timestamp 18001
transform 1 0 7452 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_5_930
timestamp 18001
transform 1 0 88596 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_1_747
timestamp 18001
transform 1 0 7452 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_5_931
timestamp 18001
transform 1 0 88596 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_1_748
timestamp 18001
transform 1 0 7452 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_78_5_932
timestamp 18001
transform 1 0 88596 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_1_749
timestamp 18001
transform 1 0 7452 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_80_5_933
timestamp 18001
transform 1 0 88596 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_1_750
timestamp 18001
transform 1 0 7452 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_82_3_934
timestamp 18001
transform 1 0 88596 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_1_751
timestamp 18001
transform 1 0 7452 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_84_3_935
timestamp 18001
transform 1 0 88596 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_1_752
timestamp 18001
transform 1 0 7452 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_86_3_936
timestamp 18001
transform 1 0 88596 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_1_753
timestamp 18001
transform 1 0 7452 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_88_3_937
timestamp 18001
transform 1 0 88596 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_1_754
timestamp 18001
transform 1 0 7452 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_90_3_938
timestamp 18001
transform 1 0 88596 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_1_755
timestamp 18001
transform 1 0 7452 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_92_3_939
timestamp 18001
transform 1 0 88596 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_1_756
timestamp 18001
transform 1 0 7452 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_94_3_940
timestamp 18001
transform 1 0 88596 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_1_757
timestamp 18001
transform 1 0 7452 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_96_3_941
timestamp 18001
transform 1 0 88596 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_1_758
timestamp 18001
transform 1 0 7452 0 1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_98_3_942
timestamp 18001
transform 1 0 88596 0 1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_1_759
timestamp 18001
transform 1 0 7452 0 1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_100_3_943
timestamp 18001
transform 1 0 88596 0 1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_1_760
timestamp 18001
transform 1 0 7452 0 1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_102_3_944
timestamp 18001
transform 1 0 88596 0 1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_1_761
timestamp 18001
transform 1 0 7452 0 1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_104_3_945
timestamp 18001
transform 1 0 88596 0 1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_1_762
timestamp 18001
transform 1 0 7452 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_106_3_946
timestamp 18001
transform 1 0 88596 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_1_763
timestamp 18001
transform 1 0 7452 0 1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_108_3_947
timestamp 18001
transform 1 0 88596 0 1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_1_764
timestamp 18001
transform 1 0 7452 0 1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_110_3_948
timestamp 18001
transform 1 0 88596 0 1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_1_765
timestamp 18001
transform 1 0 7452 0 1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_112_3_949
timestamp 18001
transform 1 0 88596 0 1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_1_766
timestamp 18001
transform 1 0 7452 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_114_3_950
timestamp 18001
transform 1 0 88596 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_1_767
timestamp 18001
transform 1 0 7452 0 1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_116_3_951
timestamp 18001
transform 1 0 88596 0 1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_1_768
timestamp 18001
transform 1 0 7452 0 1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_118_3_952
timestamp 18001
transform 1 0 88596 0 1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_1_769
timestamp 18001
transform 1 0 7452 0 1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_120_3_953
timestamp 18001
transform 1 0 88596 0 1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_1_770
timestamp 18001
transform 1 0 7452 0 1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_122_3_954
timestamp 18001
transform 1 0 88596 0 1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_1_771
timestamp 18001
transform 1 0 7452 0 1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_124_3_955
timestamp 18001
transform 1 0 88596 0 1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_1_772
timestamp 18001
transform 1 0 7452 0 1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_126_3_956
timestamp 18001
transform 1 0 88596 0 1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_1_773
timestamp 18001
transform 1 0 7452 0 1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_128_3_957
timestamp 18001
transform 1 0 88596 0 1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_1_774
timestamp 18001
transform 1 0 7452 0 1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_130_3_958
timestamp 18001
transform 1 0 88596 0 1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_1_775
timestamp 18001
transform 1 0 7452 0 1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_132_3_959
timestamp 18001
transform 1 0 88596 0 1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_1_776
timestamp 18001
transform 1 0 7452 0 1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_134_3_960
timestamp 18001
transform 1 0 88596 0 1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_1_777
timestamp 18001
transform 1 0 7452 0 1 78880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_136_3_961
timestamp 18001
transform 1 0 88596 0 1 78880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_1_778
timestamp 18001
transform 1 0 7452 0 1 79968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_138_3_962
timestamp 18001
transform 1 0 88596 0 1 79968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_140_1_779
timestamp 18001
transform 1 0 7452 0 1 81056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_140_3_963
timestamp 18001
transform 1 0 88596 0 1 81056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_142_1_780
timestamp 18001
transform 1 0 7452 0 1 82144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_142_3_964
timestamp 18001
transform 1 0 88596 0 1 82144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_144_1_781
timestamp 18001
transform 1 0 7452 0 1 83232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_144_3_965
timestamp 18001
transform 1 0 88596 0 1 83232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_1_782
timestamp 18001
transform 1 0 7452 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_146_3_966
timestamp 18001
transform 1 0 88596 0 1 84320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_1_783
timestamp 18001
transform 1 0 7452 0 1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_148_3_967
timestamp 18001
transform 1 0 88596 0 1 85408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_784
timestamp 18001
transform 1 0 7452 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_785
timestamp 18001
transform 1 0 10028 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_786
timestamp 18001
transform 1 0 12604 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_787
timestamp 18001
transform 1 0 15180 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_788
timestamp 18001
transform 1 0 17756 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_789
timestamp 18001
transform 1 0 20332 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_790
timestamp 18001
transform 1 0 22908 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_791
timestamp 18001
transform 1 0 25484 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_792
timestamp 18001
transform 1 0 28060 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_793
timestamp 18001
transform 1 0 30636 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_794
timestamp 18001
transform 1 0 33212 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_795
timestamp 18001
transform 1 0 35788 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_796
timestamp 18001
transform 1 0 38364 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_797
timestamp 18001
transform 1 0 40940 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_798
timestamp 18001
transform 1 0 43516 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_799
timestamp 18001
transform 1 0 46092 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_800
timestamp 18001
transform 1 0 48668 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_801
timestamp 18001
transform 1 0 51244 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_802
timestamp 18001
transform 1 0 53820 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_803
timestamp 18001
transform 1 0 56396 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_804
timestamp 18001
transform 1 0 58972 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_805
timestamp 18001
transform 1 0 61548 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_806
timestamp 18001
transform 1 0 64124 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_807
timestamp 18001
transform 1 0 66700 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_808
timestamp 18001
transform 1 0 69276 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_809
timestamp 18001
transform 1 0 71852 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_810
timestamp 18001
transform 1 0 74428 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_811
timestamp 18001
transform 1 0 77004 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_812
timestamp 18001
transform 1 0 79580 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_813
timestamp 18001
transform 1 0 82156 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_814
timestamp 18001
transform 1 0 84732 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_150_815
timestamp 18001
transform 1 0 87308 0 1 86496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_816
timestamp 18001
transform 1 0 10028 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_817
timestamp 18001
transform 1 0 15180 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_818
timestamp 18001
transform 1 0 20332 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_819
timestamp 18001
transform 1 0 25484 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_820
timestamp 18001
transform 1 0 30636 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_821
timestamp 18001
transform 1 0 35788 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_822
timestamp 18001
transform 1 0 40940 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_823
timestamp 18001
transform 1 0 46092 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_824
timestamp 18001
transform 1 0 51244 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_825
timestamp 18001
transform 1 0 56396 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_826
timestamp 18001
transform 1 0 61548 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_827
timestamp 18001
transform 1 0 66700 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_828
timestamp 18001
transform 1 0 71852 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_829
timestamp 18001
transform 1 0 77004 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_830
timestamp 18001
transform 1 0 82156 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_151_831
timestamp 18001
transform 1 0 87308 0 -1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_152_832
timestamp 18001
transform 1 0 7452 0 1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_152_833
timestamp 18001
transform 1 0 12604 0 1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_152_834
timestamp 18001
transform 1 0 17756 0 1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_152_835
timestamp 18001
transform 1 0 22908 0 1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_152_836
timestamp 18001
transform 1 0 28060 0 1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_152_837
timestamp 18001
transform 1 0 33212 0 1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_152_838
timestamp 18001
transform 1 0 38364 0 1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_152_839
timestamp 18001
transform 1 0 43516 0 1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_152_840
timestamp 18001
transform 1 0 48668 0 1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_152_841
timestamp 18001
transform 1 0 53820 0 1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_152_842
timestamp 18001
transform 1 0 58972 0 1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_152_843
timestamp 18001
transform 1 0 64124 0 1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_152_844
timestamp 18001
transform 1 0 69276 0 1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_152_845
timestamp 18001
transform 1 0 74428 0 1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_152_846
timestamp 18001
transform 1 0 79580 0 1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_152_847
timestamp 18001
transform 1 0 84732 0 1 87584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_153_848
timestamp 18001
transform 1 0 10028 0 -1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_153_849
timestamp 18001
transform 1 0 15180 0 -1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_153_850
timestamp 18001
transform 1 0 20332 0 -1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_153_851
timestamp 18001
transform 1 0 25484 0 -1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_153_852
timestamp 18001
transform 1 0 30636 0 -1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_153_853
timestamp 18001
transform 1 0 35788 0 -1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_153_854
timestamp 18001
transform 1 0 40940 0 -1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_153_855
timestamp 18001
transform 1 0 46092 0 -1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_153_856
timestamp 18001
transform 1 0 51244 0 -1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_153_857
timestamp 18001
transform 1 0 56396 0 -1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_153_858
timestamp 18001
transform 1 0 61548 0 -1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_153_859
timestamp 18001
transform 1 0 66700 0 -1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_153_860
timestamp 18001
transform 1 0 71852 0 -1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_153_861
timestamp 18001
transform 1 0 77004 0 -1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_153_862
timestamp 18001
transform 1 0 82156 0 -1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_153_863
timestamp 18001
transform 1 0 87308 0 -1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_864
timestamp 18001
transform 1 0 7452 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_865
timestamp 18001
transform 1 0 10028 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_866
timestamp 18001
transform 1 0 12604 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_867
timestamp 18001
transform 1 0 15180 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_868
timestamp 18001
transform 1 0 17756 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_869
timestamp 18001
transform 1 0 20332 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_870
timestamp 18001
transform 1 0 22908 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_871
timestamp 18001
transform 1 0 25484 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_872
timestamp 18001
transform 1 0 28060 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_873
timestamp 18001
transform 1 0 30636 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_874
timestamp 18001
transform 1 0 33212 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_875
timestamp 18001
transform 1 0 35788 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_876
timestamp 18001
transform 1 0 38364 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_877
timestamp 18001
transform 1 0 40940 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_878
timestamp 18001
transform 1 0 43516 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_879
timestamp 18001
transform 1 0 46092 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_880
timestamp 18001
transform 1 0 48668 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_881
timestamp 18001
transform 1 0 51244 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_882
timestamp 18001
transform 1 0 53820 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_883
timestamp 18001
transform 1 0 56396 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_884
timestamp 18001
transform 1 0 58972 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_885
timestamp 18001
transform 1 0 61548 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_886
timestamp 18001
transform 1 0 64124 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_887
timestamp 18001
transform 1 0 66700 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_888
timestamp 18001
transform 1 0 69276 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_889
timestamp 18001
transform 1 0 71852 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_890
timestamp 18001
transform 1 0 74428 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_891
timestamp 18001
transform 1 0 77004 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_892
timestamp 18001
transform 1 0 79580 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_893
timestamp 18001
transform 1 0 82156 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_894
timestamp 18001
transform 1 0 84732 0 1 88672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_154_895
timestamp 18001
transform 1 0 87308 0 1 88672
box -38 -48 130 592
<< labels >>
flabel metal2 s 47986 91800 48042 92600 0 FreeSans 224 90 0 0 clk
port 0 nsew signal input
flabel metal3 s 1600 46488 2400 46608 0 FreeSans 480 0 0 0 config_data_in
port 1 nsew signal input
flabel metal3 s 91400 47848 92200 47968 0 FreeSans 480 0 0 0 config_data_out
port 2 nsew signal output
flabel metal2 s 49918 91800 49974 92600 0 FreeSans 224 90 0 0 config_en
port 3 nsew signal input
flabel metal3 s 91400 28808 92200 28928 0 FreeSans 480 0 0 0 io_east_in[0]
port 4 nsew signal input
flabel metal3 s 91400 39688 92200 39808 0 FreeSans 480 0 0 0 io_east_in[10]
port 5 nsew signal input
flabel metal3 s 91400 41048 92200 41168 0 FreeSans 480 0 0 0 io_east_in[11]
port 6 nsew signal input
flabel metal3 s 91400 41728 92200 41848 0 FreeSans 480 0 0 0 io_east_in[12]
port 7 nsew signal input
flabel metal3 s 91400 43088 92200 43208 0 FreeSans 480 0 0 0 io_east_in[13]
port 8 nsew signal input
flabel metal2 s 1618 1600 1674 2400 0 FreeSans 224 90 0 0 io_east_in[14]
port 9 nsew signal input
flabel metal2 s 2262 1600 2318 2400 0 FreeSans 224 90 0 0 io_east_in[15]
port 10 nsew signal input
flabel metal3 s 91400 66208 92200 66328 0 FreeSans 480 0 0 0 io_east_in[16]
port 11 nsew signal input
flabel metal3 s 91400 67568 92200 67688 0 FreeSans 480 0 0 0 io_east_in[17]
port 12 nsew signal input
flabel metal3 s 91400 68248 92200 68368 0 FreeSans 480 0 0 0 io_east_in[18]
port 13 nsew signal input
flabel metal3 s 91400 69608 92200 69728 0 FreeSans 480 0 0 0 io_east_in[19]
port 14 nsew signal input
flabel metal3 s 91400 30168 92200 30288 0 FreeSans 480 0 0 0 io_east_in[1]
port 15 nsew signal input
flabel metal3 s 91400 70288 92200 70408 0 FreeSans 480 0 0 0 io_east_in[20]
port 16 nsew signal input
flabel metal3 s 91400 71648 92200 71768 0 FreeSans 480 0 0 0 io_east_in[21]
port 17 nsew signal input
flabel metal3 s 91400 73008 92200 73128 0 FreeSans 480 0 0 0 io_east_in[22]
port 18 nsew signal input
flabel metal3 s 91400 73688 92200 73808 0 FreeSans 480 0 0 0 io_east_in[23]
port 19 nsew signal input
flabel metal3 s 91400 75048 92200 75168 0 FreeSans 480 0 0 0 io_east_in[24]
port 20 nsew signal input
flabel metal3 s 91400 75728 92200 75848 0 FreeSans 480 0 0 0 io_east_in[25]
port 21 nsew signal input
flabel metal3 s 91400 77088 92200 77208 0 FreeSans 480 0 0 0 io_east_in[26]
port 22 nsew signal input
flabel metal3 s 91400 78448 92200 78568 0 FreeSans 480 0 0 0 io_east_in[27]
port 23 nsew signal input
flabel metal3 s 91400 79128 92200 79248 0 FreeSans 480 0 0 0 io_east_in[28]
port 24 nsew signal input
flabel metal3 s 91400 80488 92200 80608 0 FreeSans 480 0 0 0 io_east_in[29]
port 25 nsew signal input
flabel metal3 s 91400 30848 92200 30968 0 FreeSans 480 0 0 0 io_east_in[2]
port 26 nsew signal input
flabel metal2 s 2906 1600 2962 2400 0 FreeSans 224 90 0 0 io_east_in[30]
port 27 nsew signal input
flabel metal2 s 3550 1600 3606 2400 0 FreeSans 224 90 0 0 io_east_in[31]
port 28 nsew signal input
flabel metal3 s 91400 32208 92200 32328 0 FreeSans 480 0 0 0 io_east_in[3]
port 29 nsew signal input
flabel metal3 s 91400 32888 92200 33008 0 FreeSans 480 0 0 0 io_east_in[4]
port 30 nsew signal input
flabel metal3 s 91400 34248 92200 34368 0 FreeSans 480 0 0 0 io_east_in[5]
port 31 nsew signal input
flabel metal3 s 91400 35608 92200 35728 0 FreeSans 480 0 0 0 io_east_in[6]
port 32 nsew signal input
flabel metal3 s 91400 36288 92200 36408 0 FreeSans 480 0 0 0 io_east_in[7]
port 33 nsew signal input
flabel metal3 s 91400 37648 92200 37768 0 FreeSans 480 0 0 0 io_east_in[8]
port 34 nsew signal input
flabel metal3 s 91400 38328 92200 38448 0 FreeSans 480 0 0 0 io_east_in[9]
port 35 nsew signal input
flabel metal3 s 91400 13848 92200 13968 0 FreeSans 480 0 0 0 io_east_out[0]
port 36 nsew signal output
flabel metal3 s 91400 24728 92200 24848 0 FreeSans 480 0 0 0 io_east_out[10]
port 37 nsew signal output
flabel metal3 s 91400 25408 92200 25528 0 FreeSans 480 0 0 0 io_east_out[11]
port 38 nsew signal output
flabel metal3 s 91400 26768 92200 26888 0 FreeSans 480 0 0 0 io_east_out[12]
port 39 nsew signal output
flabel metal3 s 91400 27448 92200 27568 0 FreeSans 480 0 0 0 io_east_out[13]
port 40 nsew signal output
flabel metal3 s 1600 44448 2400 44568 0 FreeSans 480 0 0 0 io_east_out[14]
port 41 nsew signal output
flabel metal3 s 1600 49208 2400 49328 0 FreeSans 480 0 0 0 io_east_out[15]
port 42 nsew signal output
flabel metal3 s 91400 51248 92200 51368 0 FreeSans 480 0 0 0 io_east_out[16]
port 43 nsew signal output
flabel metal3 s 91400 51928 92200 52048 0 FreeSans 480 0 0 0 io_east_out[17]
port 44 nsew signal output
flabel metal3 s 91400 53288 92200 53408 0 FreeSans 480 0 0 0 io_east_out[18]
port 45 nsew signal output
flabel metal3 s 91400 53968 92200 54088 0 FreeSans 480 0 0 0 io_east_out[19]
port 46 nsew signal output
flabel metal3 s 91400 14528 92200 14648 0 FreeSans 480 0 0 0 io_east_out[1]
port 47 nsew signal output
flabel metal3 s 91400 55328 92200 55448 0 FreeSans 480 0 0 0 io_east_out[20]
port 48 nsew signal output
flabel metal3 s 91400 56688 92200 56808 0 FreeSans 480 0 0 0 io_east_out[21]
port 49 nsew signal output
flabel metal3 s 91400 57368 92200 57488 0 FreeSans 480 0 0 0 io_east_out[22]
port 50 nsew signal output
flabel metal3 s 91400 58728 92200 58848 0 FreeSans 480 0 0 0 io_east_out[23]
port 51 nsew signal output
flabel metal3 s 91400 59408 92200 59528 0 FreeSans 480 0 0 0 io_east_out[24]
port 52 nsew signal output
flabel metal3 s 91400 60768 92200 60888 0 FreeSans 480 0 0 0 io_east_out[25]
port 53 nsew signal output
flabel metal3 s 91400 62128 92200 62248 0 FreeSans 480 0 0 0 io_east_out[26]
port 54 nsew signal output
flabel metal3 s 91400 62808 92200 62928 0 FreeSans 480 0 0 0 io_east_out[27]
port 55 nsew signal output
flabel metal3 s 91400 64168 92200 64288 0 FreeSans 480 0 0 0 io_east_out[28]
port 56 nsew signal output
flabel metal3 s 91400 64848 92200 64968 0 FreeSans 480 0 0 0 io_east_out[29]
port 57 nsew signal output
flabel metal3 s 91400 15888 92200 16008 0 FreeSans 480 0 0 0 io_east_out[2]
port 58 nsew signal output
flabel metal3 s 1600 33568 2400 33688 0 FreeSans 480 0 0 0 io_east_out[30]
port 59 nsew signal output
flabel metal3 s 1600 45808 2400 45928 0 FreeSans 480 0 0 0 io_east_out[31]
port 60 nsew signal output
flabel metal3 s 91400 16568 92200 16688 0 FreeSans 480 0 0 0 io_east_out[3]
port 61 nsew signal output
flabel metal3 s 91400 17928 92200 18048 0 FreeSans 480 0 0 0 io_east_out[4]
port 62 nsew signal output
flabel metal3 s 91400 19288 92200 19408 0 FreeSans 480 0 0 0 io_east_out[5]
port 63 nsew signal output
flabel metal3 s 91400 19968 92200 20088 0 FreeSans 480 0 0 0 io_east_out[6]
port 64 nsew signal output
flabel metal3 s 91400 21328 92200 21448 0 FreeSans 480 0 0 0 io_east_out[7]
port 65 nsew signal output
flabel metal3 s 91400 22008 92200 22128 0 FreeSans 480 0 0 0 io_east_out[8]
port 66 nsew signal output
flabel metal3 s 91400 23368 92200 23488 0 FreeSans 480 0 0 0 io_east_out[9]
port 67 nsew signal output
flabel metal2 s 15786 91800 15842 92600 0 FreeSans 224 90 0 0 io_north_in[0]
port 68 nsew signal input
flabel metal2 s 26734 91800 26790 92600 0 FreeSans 224 90 0 0 io_north_in[10]
port 69 nsew signal input
flabel metal2 s 27378 91800 27434 92600 0 FreeSans 224 90 0 0 io_north_in[11]
port 70 nsew signal input
flabel metal2 s 28666 91800 28722 92600 0 FreeSans 224 90 0 0 io_north_in[12]
port 71 nsew signal input
flabel metal2 s 29954 91800 30010 92600 0 FreeSans 224 90 0 0 io_north_in[13]
port 72 nsew signal input
flabel metal2 s 4194 1600 4250 2400 0 FreeSans 224 90 0 0 io_north_in[14]
port 73 nsew signal input
flabel metal2 s 4838 1600 4894 2400 0 FreeSans 224 90 0 0 io_north_in[15]
port 74 nsew signal input
flabel metal2 s 52494 91800 52550 92600 0 FreeSans 224 90 0 0 io_north_in[16]
port 75 nsew signal input
flabel metal2 s 53782 91800 53838 92600 0 FreeSans 224 90 0 0 io_north_in[17]
port 76 nsew signal input
flabel metal2 s 54426 91800 54482 92600 0 FreeSans 224 90 0 0 io_north_in[18]
port 77 nsew signal input
flabel metal2 s 55714 91800 55770 92600 0 FreeSans 224 90 0 0 io_north_in[19]
port 78 nsew signal input
flabel metal2 s 16430 91800 16486 92600 0 FreeSans 224 90 0 0 io_north_in[1]
port 79 nsew signal input
flabel metal2 s 57002 91800 57058 92600 0 FreeSans 224 90 0 0 io_north_in[20]
port 80 nsew signal input
flabel metal2 s 58290 91800 58346 92600 0 FreeSans 224 90 0 0 io_north_in[21]
port 81 nsew signal input
flabel metal2 s 58934 91800 58990 92600 0 FreeSans 224 90 0 0 io_north_in[22]
port 82 nsew signal input
flabel metal2 s 60222 91800 60278 92600 0 FreeSans 224 90 0 0 io_north_in[23]
port 83 nsew signal input
flabel metal2 s 61510 91800 61566 92600 0 FreeSans 224 90 0 0 io_north_in[24]
port 84 nsew signal input
flabel metal2 s 62154 91800 62210 92600 0 FreeSans 224 90 0 0 io_north_in[25]
port 85 nsew signal input
flabel metal2 s 63442 91800 63498 92600 0 FreeSans 224 90 0 0 io_north_in[26]
port 86 nsew signal input
flabel metal2 s 64730 91800 64786 92600 0 FreeSans 224 90 0 0 io_north_in[27]
port 87 nsew signal input
flabel metal2 s 66018 91800 66074 92600 0 FreeSans 224 90 0 0 io_north_in[28]
port 88 nsew signal input
flabel metal2 s 66662 91800 66718 92600 0 FreeSans 224 90 0 0 io_north_in[29]
port 89 nsew signal input
flabel metal2 s 17718 91800 17774 92600 0 FreeSans 224 90 0 0 io_north_in[2]
port 90 nsew signal input
flabel metal2 s 5482 1600 5538 2400 0 FreeSans 224 90 0 0 io_north_in[30]
port 91 nsew signal input
flabel metal2 s 6126 1600 6182 2400 0 FreeSans 224 90 0 0 io_north_in[31]
port 92 nsew signal input
flabel metal2 s 19006 91800 19062 92600 0 FreeSans 224 90 0 0 io_north_in[3]
port 93 nsew signal input
flabel metal2 s 19650 91800 19706 92600 0 FreeSans 224 90 0 0 io_north_in[4]
port 94 nsew signal input
flabel metal2 s 20938 91800 20994 92600 0 FreeSans 224 90 0 0 io_north_in[5]
port 95 nsew signal input
flabel metal2 s 22226 91800 22282 92600 0 FreeSans 224 90 0 0 io_north_in[6]
port 96 nsew signal input
flabel metal2 s 23514 91800 23570 92600 0 FreeSans 224 90 0 0 io_north_in[7]
port 97 nsew signal input
flabel metal2 s 24158 91800 24214 92600 0 FreeSans 224 90 0 0 io_north_in[8]
port 98 nsew signal input
flabel metal2 s 25446 91800 25502 92600 0 FreeSans 224 90 0 0 io_north_in[9]
port 99 nsew signal input
flabel metal2 s 31242 91800 31298 92600 0 FreeSans 224 90 0 0 io_north_out[0]
port 100 nsew signal output
flabel metal2 s 42190 91800 42246 92600 0 FreeSans 224 90 0 0 io_north_out[10]
port 101 nsew signal output
flabel metal2 s 42834 91800 42890 92600 0 FreeSans 224 90 0 0 io_north_out[11]
port 102 nsew signal output
flabel metal2 s 44122 91800 44178 92600 0 FreeSans 224 90 0 0 io_north_out[12]
port 103 nsew signal output
flabel metal2 s 45410 91800 45466 92600 0 FreeSans 224 90 0 0 io_north_out[13]
port 104 nsew signal output
flabel metal2 s 56358 91800 56414 92600 0 FreeSans 224 90 0 0 io_north_out[14]
port 105 nsew signal output
flabel metal3 s 91400 68928 92200 69048 0 FreeSans 480 0 0 0 io_north_out[15]
port 106 nsew signal output
flabel metal2 s 67950 91800 68006 92600 0 FreeSans 224 90 0 0 io_north_out[16]
port 107 nsew signal output
flabel metal2 s 69238 91800 69294 92600 0 FreeSans 224 90 0 0 io_north_out[17]
port 108 nsew signal output
flabel metal2 s 69882 91800 69938 92600 0 FreeSans 224 90 0 0 io_north_out[18]
port 109 nsew signal output
flabel metal2 s 71170 91800 71226 92600 0 FreeSans 224 90 0 0 io_north_out[19]
port 110 nsew signal output
flabel metal2 s 31886 91800 31942 92600 0 FreeSans 224 90 0 0 io_north_out[1]
port 111 nsew signal output
flabel metal2 s 72458 91800 72514 92600 0 FreeSans 224 90 0 0 io_north_out[20]
port 112 nsew signal output
flabel metal2 s 73746 91800 73802 92600 0 FreeSans 224 90 0 0 io_north_out[21]
port 113 nsew signal output
flabel metal2 s 74390 91800 74446 92600 0 FreeSans 224 90 0 0 io_north_out[22]
port 114 nsew signal output
flabel metal2 s 75678 91800 75734 92600 0 FreeSans 224 90 0 0 io_north_out[23]
port 115 nsew signal output
flabel metal2 s 76966 91800 77022 92600 0 FreeSans 224 90 0 0 io_north_out[24]
port 116 nsew signal output
flabel metal2 s 77610 91800 77666 92600 0 FreeSans 224 90 0 0 io_north_out[25]
port 117 nsew signal output
flabel metal2 s 78898 91800 78954 92600 0 FreeSans 224 90 0 0 io_north_out[26]
port 118 nsew signal output
flabel metal2 s 80186 91800 80242 92600 0 FreeSans 224 90 0 0 io_north_out[27]
port 119 nsew signal output
flabel metal2 s 81474 91800 81530 92600 0 FreeSans 224 90 0 0 io_north_out[28]
port 120 nsew signal output
flabel metal2 s 82118 91800 82174 92600 0 FreeSans 224 90 0 0 io_north_out[29]
port 121 nsew signal output
flabel metal2 s 33174 91800 33230 92600 0 FreeSans 224 90 0 0 io_north_out[2]
port 122 nsew signal output
flabel metal3 s 91400 46488 92200 46608 0 FreeSans 480 0 0 0 io_north_out[30]
port 123 nsew signal output
flabel metal2 s 57646 91800 57702 92600 0 FreeSans 224 90 0 0 io_north_out[31]
port 124 nsew signal output
flabel metal2 s 34462 91800 34518 92600 0 FreeSans 224 90 0 0 io_north_out[3]
port 125 nsew signal output
flabel metal2 s 35106 91800 35162 92600 0 FreeSans 224 90 0 0 io_north_out[4]
port 126 nsew signal output
flabel metal2 s 36394 91800 36450 92600 0 FreeSans 224 90 0 0 io_north_out[5]
port 127 nsew signal output
flabel metal2 s 37682 91800 37738 92600 0 FreeSans 224 90 0 0 io_north_out[6]
port 128 nsew signal output
flabel metal2 s 38970 91800 39026 92600 0 FreeSans 224 90 0 0 io_north_out[7]
port 129 nsew signal output
flabel metal2 s 39614 91800 39670 92600 0 FreeSans 224 90 0 0 io_north_out[8]
port 130 nsew signal output
flabel metal2 s 40902 91800 40958 92600 0 FreeSans 224 90 0 0 io_north_out[9]
port 131 nsew signal output
flabel metal2 s 31242 1600 31298 2400 0 FreeSans 224 90 0 0 io_south_in[0]
port 132 nsew signal input
flabel metal2 s 42190 1600 42246 2400 0 FreeSans 224 90 0 0 io_south_in[10]
port 133 nsew signal input
flabel metal2 s 42834 1600 42890 2400 0 FreeSans 224 90 0 0 io_south_in[11]
port 134 nsew signal input
flabel metal2 s 44122 1600 44178 2400 0 FreeSans 224 90 0 0 io_south_in[12]
port 135 nsew signal input
flabel metal2 s 45410 1600 45466 2400 0 FreeSans 224 90 0 0 io_south_in[13]
port 136 nsew signal input
flabel metal2 s 6770 1600 6826 2400 0 FreeSans 224 90 0 0 io_south_in[14]
port 137 nsew signal input
flabel metal2 s 7414 1600 7470 2400 0 FreeSans 224 90 0 0 io_south_in[15]
port 138 nsew signal input
flabel metal2 s 67950 1600 68006 2400 0 FreeSans 224 90 0 0 io_south_in[16]
port 139 nsew signal input
flabel metal2 s 69238 1600 69294 2400 0 FreeSans 224 90 0 0 io_south_in[17]
port 140 nsew signal input
flabel metal2 s 69882 1600 69938 2400 0 FreeSans 224 90 0 0 io_south_in[18]
port 141 nsew signal input
flabel metal2 s 71170 1600 71226 2400 0 FreeSans 224 90 0 0 io_south_in[19]
port 142 nsew signal input
flabel metal2 s 31886 1600 31942 2400 0 FreeSans 224 90 0 0 io_south_in[1]
port 143 nsew signal input
flabel metal2 s 72458 1600 72514 2400 0 FreeSans 224 90 0 0 io_south_in[20]
port 144 nsew signal input
flabel metal2 s 73746 1600 73802 2400 0 FreeSans 224 90 0 0 io_south_in[21]
port 145 nsew signal input
flabel metal2 s 74390 1600 74446 2400 0 FreeSans 224 90 0 0 io_south_in[22]
port 146 nsew signal input
flabel metal2 s 75678 1600 75734 2400 0 FreeSans 224 90 0 0 io_south_in[23]
port 147 nsew signal input
flabel metal2 s 76966 1600 77022 2400 0 FreeSans 224 90 0 0 io_south_in[24]
port 148 nsew signal input
flabel metal2 s 77610 1600 77666 2400 0 FreeSans 224 90 0 0 io_south_in[25]
port 149 nsew signal input
flabel metal2 s 78898 1600 78954 2400 0 FreeSans 224 90 0 0 io_south_in[26]
port 150 nsew signal input
flabel metal2 s 80186 1600 80242 2400 0 FreeSans 224 90 0 0 io_south_in[27]
port 151 nsew signal input
flabel metal2 s 81474 1600 81530 2400 0 FreeSans 224 90 0 0 io_south_in[28]
port 152 nsew signal input
flabel metal2 s 82118 1600 82174 2400 0 FreeSans 224 90 0 0 io_south_in[29]
port 153 nsew signal input
flabel metal2 s 33174 1600 33230 2400 0 FreeSans 224 90 0 0 io_south_in[2]
port 154 nsew signal input
flabel metal2 s 8058 1600 8114 2400 0 FreeSans 224 90 0 0 io_south_in[30]
port 155 nsew signal input
flabel metal2 s 8702 1600 8758 2400 0 FreeSans 224 90 0 0 io_south_in[31]
port 156 nsew signal input
flabel metal2 s 34462 1600 34518 2400 0 FreeSans 224 90 0 0 io_south_in[3]
port 157 nsew signal input
flabel metal2 s 35106 1600 35162 2400 0 FreeSans 224 90 0 0 io_south_in[4]
port 158 nsew signal input
flabel metal2 s 36394 1600 36450 2400 0 FreeSans 224 90 0 0 io_south_in[5]
port 159 nsew signal input
flabel metal2 s 37682 1600 37738 2400 0 FreeSans 224 90 0 0 io_south_in[6]
port 160 nsew signal input
flabel metal2 s 38970 1600 39026 2400 0 FreeSans 224 90 0 0 io_south_in[7]
port 161 nsew signal input
flabel metal2 s 39614 1600 39670 2400 0 FreeSans 224 90 0 0 io_south_in[8]
port 162 nsew signal input
flabel metal2 s 40902 1600 40958 2400 0 FreeSans 224 90 0 0 io_south_in[9]
port 163 nsew signal input
flabel metal2 s 15786 1600 15842 2400 0 FreeSans 224 90 0 0 io_south_out[0]
port 164 nsew signal output
flabel metal2 s 26734 1600 26790 2400 0 FreeSans 224 90 0 0 io_south_out[10]
port 165 nsew signal output
flabel metal2 s 27378 1600 27434 2400 0 FreeSans 224 90 0 0 io_south_out[11]
port 166 nsew signal output
flabel metal2 s 28666 1600 28722 2400 0 FreeSans 224 90 0 0 io_south_out[12]
port 167 nsew signal output
flabel metal2 s 29954 1600 30010 2400 0 FreeSans 224 90 0 0 io_south_out[13]
port 168 nsew signal output
flabel metal3 s 91400 48528 92200 48648 0 FreeSans 480 0 0 0 io_south_out[14]
port 169 nsew signal output
flabel metal3 s 1600 42408 2400 42528 0 FreeSans 480 0 0 0 io_south_out[15]
port 170 nsew signal output
flabel metal2 s 52494 1600 52550 2400 0 FreeSans 224 90 0 0 io_south_out[16]
port 171 nsew signal output
flabel metal2 s 53782 1600 53838 2400 0 FreeSans 224 90 0 0 io_south_out[17]
port 172 nsew signal output
flabel metal2 s 54426 1600 54482 2400 0 FreeSans 224 90 0 0 io_south_out[18]
port 173 nsew signal output
flabel metal2 s 55714 1600 55770 2400 0 FreeSans 224 90 0 0 io_south_out[19]
port 174 nsew signal output
flabel metal2 s 16430 1600 16486 2400 0 FreeSans 224 90 0 0 io_south_out[1]
port 175 nsew signal output
flabel metal2 s 57002 1600 57058 2400 0 FreeSans 224 90 0 0 io_south_out[20]
port 176 nsew signal output
flabel metal2 s 58290 1600 58346 2400 0 FreeSans 224 90 0 0 io_south_out[21]
port 177 nsew signal output
flabel metal2 s 58934 1600 58990 2400 0 FreeSans 224 90 0 0 io_south_out[22]
port 178 nsew signal output
flabel metal2 s 60222 1600 60278 2400 0 FreeSans 224 90 0 0 io_south_out[23]
port 179 nsew signal output
flabel metal2 s 61510 1600 61566 2400 0 FreeSans 224 90 0 0 io_south_out[24]
port 180 nsew signal output
flabel metal2 s 62154 1600 62210 2400 0 FreeSans 224 90 0 0 io_south_out[25]
port 181 nsew signal output
flabel metal2 s 63442 1600 63498 2400 0 FreeSans 224 90 0 0 io_south_out[26]
port 182 nsew signal output
flabel metal2 s 64730 1600 64786 2400 0 FreeSans 224 90 0 0 io_south_out[27]
port 183 nsew signal output
flabel metal2 s 66018 1600 66074 2400 0 FreeSans 224 90 0 0 io_south_out[28]
port 184 nsew signal output
flabel metal2 s 66662 1600 66718 2400 0 FreeSans 224 90 0 0 io_south_out[29]
port 185 nsew signal output
flabel metal2 s 17718 1600 17774 2400 0 FreeSans 224 90 0 0 io_south_out[2]
port 186 nsew signal output
flabel metal3 s 91400 49208 92200 49328 0 FreeSans 480 0 0 0 io_south_out[30]
port 187 nsew signal output
flabel metal3 s 91400 52608 92200 52728 0 FreeSans 480 0 0 0 io_south_out[31]
port 188 nsew signal output
flabel metal2 s 19006 1600 19062 2400 0 FreeSans 224 90 0 0 io_south_out[3]
port 189 nsew signal output
flabel metal2 s 19650 1600 19706 2400 0 FreeSans 224 90 0 0 io_south_out[4]
port 190 nsew signal output
flabel metal2 s 20938 1600 20994 2400 0 FreeSans 224 90 0 0 io_south_out[5]
port 191 nsew signal output
flabel metal2 s 22226 1600 22282 2400 0 FreeSans 224 90 0 0 io_south_out[6]
port 192 nsew signal output
flabel metal2 s 23514 1600 23570 2400 0 FreeSans 224 90 0 0 io_south_out[7]
port 193 nsew signal output
flabel metal2 s 24158 1600 24214 2400 0 FreeSans 224 90 0 0 io_south_out[8]
port 194 nsew signal output
flabel metal2 s 25446 1600 25502 2400 0 FreeSans 224 90 0 0 io_south_out[9]
port 195 nsew signal output
flabel metal3 s 1600 13848 2400 13968 0 FreeSans 480 0 0 0 io_west_in[0]
port 196 nsew signal input
flabel metal3 s 1600 24728 2400 24848 0 FreeSans 480 0 0 0 io_west_in[10]
port 197 nsew signal input
flabel metal3 s 1600 25408 2400 25528 0 FreeSans 480 0 0 0 io_west_in[11]
port 198 nsew signal input
flabel metal3 s 1600 26768 2400 26888 0 FreeSans 480 0 0 0 io_west_in[12]
port 199 nsew signal input
flabel metal3 s 1600 27448 2400 27568 0 FreeSans 480 0 0 0 io_west_in[13]
port 200 nsew signal input
flabel metal2 s 9346 1600 9402 2400 0 FreeSans 224 90 0 0 io_west_in[14]
port 201 nsew signal input
flabel metal2 s 9990 1600 10046 2400 0 FreeSans 224 90 0 0 io_west_in[15]
port 202 nsew signal input
flabel metal3 s 1600 51248 2400 51368 0 FreeSans 480 0 0 0 io_west_in[16]
port 203 nsew signal input
flabel metal3 s 1600 51928 2400 52048 0 FreeSans 480 0 0 0 io_west_in[17]
port 204 nsew signal input
flabel metal3 s 1600 52608 2400 52728 0 FreeSans 480 0 0 0 io_west_in[18]
port 205 nsew signal input
flabel metal3 s 1600 53288 2400 53408 0 FreeSans 480 0 0 0 io_west_in[19]
port 206 nsew signal input
flabel metal3 s 1600 14528 2400 14648 0 FreeSans 480 0 0 0 io_west_in[1]
port 207 nsew signal input
flabel metal3 s 1600 55328 2400 55448 0 FreeSans 480 0 0 0 io_west_in[20]
port 208 nsew signal input
flabel metal3 s 1600 56688 2400 56808 0 FreeSans 480 0 0 0 io_west_in[21]
port 209 nsew signal input
flabel metal3 s 1600 57368 2400 57488 0 FreeSans 480 0 0 0 io_west_in[22]
port 210 nsew signal input
flabel metal3 s 1600 58728 2400 58848 0 FreeSans 480 0 0 0 io_west_in[23]
port 211 nsew signal input
flabel metal3 s 1600 59408 2400 59528 0 FreeSans 480 0 0 0 io_west_in[24]
port 212 nsew signal input
flabel metal3 s 1600 60768 2400 60888 0 FreeSans 480 0 0 0 io_west_in[25]
port 213 nsew signal input
flabel metal3 s 1600 62128 2400 62248 0 FreeSans 480 0 0 0 io_west_in[26]
port 214 nsew signal input
flabel metal3 s 1600 62808 2400 62928 0 FreeSans 480 0 0 0 io_west_in[27]
port 215 nsew signal input
flabel metal3 s 1600 64168 2400 64288 0 FreeSans 480 0 0 0 io_west_in[28]
port 216 nsew signal input
flabel metal3 s 1600 64848 2400 64968 0 FreeSans 480 0 0 0 io_west_in[29]
port 217 nsew signal input
flabel metal3 s 1600 15888 2400 16008 0 FreeSans 480 0 0 0 io_west_in[2]
port 218 nsew signal input
flabel metal2 s 10634 1600 10690 2400 0 FreeSans 224 90 0 0 io_west_in[30]
port 219 nsew signal input
flabel metal2 s 11278 1600 11334 2400 0 FreeSans 224 90 0 0 io_west_in[31]
port 220 nsew signal input
flabel metal3 s 1600 16568 2400 16688 0 FreeSans 480 0 0 0 io_west_in[3]
port 221 nsew signal input
flabel metal3 s 1600 17928 2400 18048 0 FreeSans 480 0 0 0 io_west_in[4]
port 222 nsew signal input
flabel metal3 s 1600 19288 2400 19408 0 FreeSans 480 0 0 0 io_west_in[5]
port 223 nsew signal input
flabel metal3 s 1600 19968 2400 20088 0 FreeSans 480 0 0 0 io_west_in[6]
port 224 nsew signal input
flabel metal3 s 1600 21328 2400 21448 0 FreeSans 480 0 0 0 io_west_in[7]
port 225 nsew signal input
flabel metal3 s 1600 22008 2400 22128 0 FreeSans 480 0 0 0 io_west_in[8]
port 226 nsew signal input
flabel metal3 s 1600 23368 2400 23488 0 FreeSans 480 0 0 0 io_west_in[9]
port 227 nsew signal input
flabel metal3 s 1600 28808 2400 28928 0 FreeSans 480 0 0 0 io_west_out[0]
port 228 nsew signal output
flabel metal3 s 1600 39688 2400 39808 0 FreeSans 480 0 0 0 io_west_out[10]
port 229 nsew signal output
flabel metal3 s 1600 41048 2400 41168 0 FreeSans 480 0 0 0 io_west_out[11]
port 230 nsew signal output
flabel metal3 s 1600 41728 2400 41848 0 FreeSans 480 0 0 0 io_west_out[12]
port 231 nsew signal output
flabel metal3 s 1600 43088 2400 43208 0 FreeSans 480 0 0 0 io_west_out[13]
port 232 nsew signal output
flabel metal2 s 46698 91800 46754 92600 0 FreeSans 224 90 0 0 io_west_out[14]
port 233 nsew signal output
flabel metal3 s 1600 53968 2400 54088 0 FreeSans 480 0 0 0 io_west_out[15]
port 234 nsew signal output
flabel metal3 s 1600 66208 2400 66328 0 FreeSans 480 0 0 0 io_west_out[16]
port 235 nsew signal output
flabel metal3 s 1600 67568 2400 67688 0 FreeSans 480 0 0 0 io_west_out[17]
port 236 nsew signal output
flabel metal3 s 1600 68248 2400 68368 0 FreeSans 480 0 0 0 io_west_out[18]
port 237 nsew signal output
flabel metal3 s 1600 69608 2400 69728 0 FreeSans 480 0 0 0 io_west_out[19]
port 238 nsew signal output
flabel metal3 s 1600 30168 2400 30288 0 FreeSans 480 0 0 0 io_west_out[1]
port 239 nsew signal output
flabel metal3 s 1600 70288 2400 70408 0 FreeSans 480 0 0 0 io_west_out[20]
port 240 nsew signal output
flabel metal3 s 1600 71648 2400 71768 0 FreeSans 480 0 0 0 io_west_out[21]
port 241 nsew signal output
flabel metal3 s 1600 73008 2400 73128 0 FreeSans 480 0 0 0 io_west_out[22]
port 242 nsew signal output
flabel metal3 s 1600 73688 2400 73808 0 FreeSans 480 0 0 0 io_west_out[23]
port 243 nsew signal output
flabel metal3 s 1600 75048 2400 75168 0 FreeSans 480 0 0 0 io_west_out[24]
port 244 nsew signal output
flabel metal3 s 1600 75728 2400 75848 0 FreeSans 480 0 0 0 io_west_out[25]
port 245 nsew signal output
flabel metal3 s 1600 77088 2400 77208 0 FreeSans 480 0 0 0 io_west_out[26]
port 246 nsew signal output
flabel metal3 s 1600 78448 2400 78568 0 FreeSans 480 0 0 0 io_west_out[27]
port 247 nsew signal output
flabel metal3 s 1600 79128 2400 79248 0 FreeSans 480 0 0 0 io_west_out[28]
port 248 nsew signal output
flabel metal3 s 1600 80488 2400 80608 0 FreeSans 480 0 0 0 io_west_out[29]
port 249 nsew signal output
flabel metal3 s 1600 30848 2400 30968 0 FreeSans 480 0 0 0 io_west_out[2]
port 250 nsew signal output
flabel metal3 s 1600 54648 2400 54768 0 FreeSans 480 0 0 0 io_west_out[30]
port 251 nsew signal output
flabel metal3 s 1600 43768 2400 43888 0 FreeSans 480 0 0 0 io_west_out[31]
port 252 nsew signal output
flabel metal3 s 1600 32208 2400 32328 0 FreeSans 480 0 0 0 io_west_out[3]
port 253 nsew signal output
flabel metal3 s 1600 32888 2400 33008 0 FreeSans 480 0 0 0 io_west_out[4]
port 254 nsew signal output
flabel metal3 s 1600 34248 2400 34368 0 FreeSans 480 0 0 0 io_west_out[5]
port 255 nsew signal output
flabel metal3 s 1600 35608 2400 35728 0 FreeSans 480 0 0 0 io_west_out[6]
port 256 nsew signal output
flabel metal3 s 1600 36288 2400 36408 0 FreeSans 480 0 0 0 io_west_out[7]
port 257 nsew signal output
flabel metal3 s 1600 37648 2400 37768 0 FreeSans 480 0 0 0 io_west_out[8]
port 258 nsew signal output
flabel metal3 s 1600 38328 2400 38448 0 FreeSans 480 0 0 0 io_west_out[9]
port 259 nsew signal output
flabel metal2 s 12566 1600 12622 2400 0 FreeSans 224 90 0 0 le_clk
port 260 nsew signal input
flabel metal2 s 13854 1600 13910 2400 0 FreeSans 224 90 0 0 le_en
port 261 nsew signal input
flabel metal2 s 14498 1600 14554 2400 0 FreeSans 224 90 0 0 le_nrst
port 262 nsew signal input
flabel metal2 s 48630 91800 48686 92600 0 FreeSans 224 90 0 0 nrst
port 263 nsew signal input
flabel metal4 s 3356 3376 3676 90736 0 FreeSans 1920 90 0 0 vccd1
port 264 nsew power bidirectional
flabel metal5 s 3356 3376 90484 3696 0 FreeSans 2560 0 0 0 vccd1
port 264 nsew power bidirectional
flabel metal5 s 3356 90416 90484 90736 0 FreeSans 2560 0 0 0 vccd1
port 264 nsew power bidirectional
flabel metal4 s 90164 3376 90484 90736 0 FreeSans 1920 90 0 0 vccd1
port 264 nsew power bidirectional
flabel metal4 s 18716 2716 19036 8927 0 FreeSans 1920 90 0 0 vccd1
port 264 nsew power bidirectional
flabel metal4 s 18716 85601 19036 91396 0 FreeSans 1920 90 0 0 vccd1
port 264 nsew power bidirectional
flabel metal4 s 37716 2716 38036 8927 0 FreeSans 1920 90 0 0 vccd1
port 264 nsew power bidirectional
flabel metal4 s 37716 85601 38036 91396 0 FreeSans 1920 90 0 0 vccd1
port 264 nsew power bidirectional
flabel metal4 s 56716 2716 57036 8927 0 FreeSans 1920 90 0 0 vccd1
port 264 nsew power bidirectional
flabel metal4 s 56716 85601 57036 91396 0 FreeSans 1920 90 0 0 vccd1
port 264 nsew power bidirectional
flabel metal4 s 75716 2716 76036 8927 0 FreeSans 1920 90 0 0 vccd1
port 264 nsew power bidirectional
flabel metal4 s 75716 85601 76036 91396 0 FreeSans 1920 90 0 0 vccd1
port 264 nsew power bidirectional
flabel metal5 s 2696 18736 91144 19056 0 FreeSans 2560 0 0 0 vccd1
port 264 nsew power bidirectional
flabel metal5 s 2696 37736 91144 38056 0 FreeSans 2560 0 0 0 vccd1
port 264 nsew power bidirectional
flabel metal5 s 2696 56736 91144 57056 0 FreeSans 2560 0 0 0 vccd1
port 264 nsew power bidirectional
flabel metal5 s 2696 75736 91144 76056 0 FreeSans 2560 0 0 0 vccd1
port 264 nsew power bidirectional
flabel metal4 s 5948 7024 6268 87088 0 FreeSans 1920 90 0 0 vccd1
port 264 nsew power bidirectional
flabel metal4 s 87092 7024 87412 87088 0 FreeSans 1920 90 0 0 vccd1
port 264 nsew power bidirectional
flabel metal4 s 2696 2716 3016 91396 0 FreeSans 1920 90 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal5 s 2696 2716 91144 3036 0 FreeSans 2560 0 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal5 s 2696 91076 91144 91396 0 FreeSans 2560 0 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal4 s 90824 2716 91144 91396 0 FreeSans 1920 90 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal4 s 19376 2716 19696 8927 0 FreeSans 1920 90 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal4 s 19376 85601 19696 91396 0 FreeSans 1920 90 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal4 s 38376 2716 38696 8927 0 FreeSans 1920 90 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal4 s 38376 85601 38696 91396 0 FreeSans 1920 90 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal4 s 57376 2716 57696 8927 0 FreeSans 1920 90 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal4 s 57376 85601 57696 91396 0 FreeSans 1920 90 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal4 s 76376 2716 76696 8927 0 FreeSans 1920 90 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal4 s 76376 85601 76696 91396 0 FreeSans 1920 90 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal5 s 2696 19396 91144 19716 0 FreeSans 2560 0 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal5 s 2696 38396 91144 38716 0 FreeSans 2560 0 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal5 s 2696 57396 91144 57716 0 FreeSans 2560 0 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal5 s 2696 76396 91144 76716 0 FreeSans 2560 0 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal4 s 6684 7024 7004 87088 0 FreeSans 1920 90 0 0 vssd1
port 265 nsew ground bidirectional
flabel metal4 s 87828 7024 88148 87088 0 FreeSans 1920 90 0 0 vssd1
port 265 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 1600 1600 92200 92600
<< end >>
