VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO intro_2_stopwatch
  CLASS BLOCK ;
  FOREIGN intro_2_stopwatch ;
  ORIGIN 0.000 0.000 ;
  SIZE 145.100 BY 155.820 ;
  PIN BTN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 41.950 151.820 42.230 155.820 ;
    END
  END BTN[0]
  PIN BTN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END BTN[1]
  PIN BTN[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END BTN[2]
  PIN BTN[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END BTN[3]
  PIN CLK_10MHZ
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END CLK_10MHZ
  PIN D0_AN_0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END D0_AN_0
  PIN D0_AN_1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 45.170 151.820 45.450 155.820 ;
    END
  END D0_AN_1
  PIN D0_AN_2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END D0_AN_2
  PIN D0_AN_3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 151.820 16.470 155.820 ;
    END
  END D0_AN_3
  PIN D0_SEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END D0_SEG[0]
  PIN D0_SEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END D0_SEG[1]
  PIN D0_SEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 29.070 151.820 29.350 155.820 ;
    END
  END D0_SEG[2]
  PIN D0_SEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END D0_SEG[3]
  PIN D0_SEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END D0_SEG[4]
  PIN D0_SEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 32.290 151.820 32.570 155.820 ;
    END
  END D0_SEG[5]
  PIN D0_SEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 35.510 151.820 35.790 155.820 ;
    END
  END D0_SEG[6]
  PIN D0_SEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 141.100 13.640 145.100 14.240 ;
    END
  END D0_SEG[7]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 144.400 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 144.400 ;
    END
  END VPWR
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 139.570 144.350 ;
      LAYER li1 ;
        RECT 5.520 10.795 139.380 144.245 ;
      LAYER met1 ;
        RECT 4.210 10.640 139.380 144.400 ;
      LAYER met2 ;
        RECT 4.230 151.540 15.910 151.820 ;
        RECT 16.750 151.540 28.790 151.820 ;
        RECT 29.630 151.540 32.010 151.820 ;
        RECT 32.850 151.540 35.230 151.820 ;
        RECT 36.070 151.540 41.670 151.820 ;
        RECT 42.510 151.540 44.890 151.820 ;
        RECT 45.730 151.540 137.910 151.820 ;
        RECT 4.230 10.695 137.910 151.540 ;
      LAYER met3 ;
        RECT 3.990 140.440 141.100 144.325 ;
        RECT 4.400 139.040 141.100 140.440 ;
        RECT 3.990 133.640 141.100 139.040 ;
        RECT 4.400 132.240 141.100 133.640 ;
        RECT 3.990 130.240 141.100 132.240 ;
        RECT 4.400 128.840 141.100 130.240 ;
        RECT 3.990 126.840 141.100 128.840 ;
        RECT 4.400 125.440 141.100 126.840 ;
        RECT 3.990 123.440 141.100 125.440 ;
        RECT 4.400 122.040 141.100 123.440 ;
        RECT 3.990 120.040 141.100 122.040 ;
        RECT 4.400 118.640 141.100 120.040 ;
        RECT 3.990 116.640 141.100 118.640 ;
        RECT 4.400 115.240 141.100 116.640 ;
        RECT 3.990 106.440 141.100 115.240 ;
        RECT 4.400 105.040 141.100 106.440 ;
        RECT 3.990 99.640 141.100 105.040 ;
        RECT 4.400 98.240 141.100 99.640 ;
        RECT 3.990 14.640 141.100 98.240 ;
        RECT 4.400 13.240 140.700 14.640 ;
        RECT 3.990 10.715 141.100 13.240 ;
      LAYER met4 ;
        RECT 118.975 19.895 128.505 76.665 ;
  END
END intro_2_stopwatch
END LIBRARY

