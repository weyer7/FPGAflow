magic
tech sky130A
magscale 1 2
timestamp 1746144263
<< viali >>
rect 9229 25925 9263 25959
rect 9873 25925 9907 25959
rect 10517 25925 10551 25959
rect 12449 25925 12483 25959
rect 13737 25925 13771 25959
rect 14381 25925 14415 25959
rect 15025 25925 15059 25959
rect 17601 25925 17635 25959
rect 18245 25925 18279 25959
rect 3985 25857 4019 25891
rect 11253 25857 11287 25891
rect 11713 25857 11747 25891
rect 13001 25857 13035 25891
rect 15577 25857 15611 25891
rect 16221 25857 16255 25891
rect 4261 25789 4295 25823
rect 10057 25789 10091 25823
rect 15209 25789 15243 25823
rect 12633 25721 12667 25755
rect 13921 25721 13955 25755
rect 14565 25721 14599 25755
rect 15761 25721 15795 25755
rect 18429 25721 18463 25755
rect 3801 25653 3835 25687
rect 4169 25653 4203 25687
rect 9321 25653 9355 25687
rect 10609 25653 10643 25687
rect 11069 25653 11103 25687
rect 11897 25653 11931 25687
rect 13185 25653 13219 25687
rect 16405 25653 16439 25687
rect 17693 25653 17727 25687
rect 4445 25449 4479 25483
rect 4721 25449 4755 25483
rect 2053 25313 2087 25347
rect 3525 25313 3559 25347
rect 3801 25313 3835 25347
rect 13369 25313 13403 25347
rect 19257 25313 19291 25347
rect 1777 25245 1811 25279
rect 4537 25245 4571 25279
rect 4721 25245 4755 25279
rect 4813 25245 4847 25279
rect 4997 25245 5031 25279
rect 6009 25245 6043 25279
rect 8217 25245 8251 25279
rect 8309 25245 8343 25279
rect 8953 25245 8987 25279
rect 11069 25245 11103 25279
rect 13001 25245 13035 25279
rect 13277 25245 13311 25279
rect 15577 25245 15611 25279
rect 24869 25245 24903 25279
rect 7665 25177 7699 25211
rect 7849 25177 7883 25211
rect 9229 25177 9263 25211
rect 12725 25177 12759 25211
rect 15853 25177 15887 25211
rect 19533 25177 19567 25211
rect 4905 25109 4939 25143
rect 5457 25109 5491 25143
rect 8033 25109 8067 25143
rect 8493 25109 8527 25143
rect 10701 25109 10735 25143
rect 10977 25109 11011 25143
rect 11253 25109 11287 25143
rect 13645 25109 13679 25143
rect 17325 25109 17359 25143
rect 21005 25109 21039 25143
rect 5917 24905 5951 24939
rect 9137 24905 9171 24939
rect 14841 24905 14875 24939
rect 15669 24905 15703 24939
rect 18245 24905 18279 24939
rect 8953 24837 8987 24871
rect 17049 24837 17083 24871
rect 8493 24769 8527 24803
rect 9229 24769 9263 24803
rect 9413 24769 9447 24803
rect 9689 24769 9723 24803
rect 12633 24769 12667 24803
rect 15117 24769 15151 24803
rect 15209 24769 15243 24803
rect 15761 24769 15795 24803
rect 16037 24769 16071 24803
rect 16865 24769 16899 24803
rect 17141 24769 17175 24803
rect 17233 24769 17267 24803
rect 17417 24769 17451 24803
rect 17785 24769 17819 24803
rect 18061 24769 18095 24803
rect 18245 24769 18279 24803
rect 19165 24769 19199 24803
rect 19257 24769 19291 24803
rect 22201 24769 22235 24803
rect 22477 24769 22511 24803
rect 22661 24769 22695 24803
rect 1501 24701 1535 24735
rect 1777 24701 1811 24735
rect 3249 24701 3283 24735
rect 3893 24701 3927 24735
rect 4169 24701 4203 24735
rect 4445 24701 4479 24735
rect 8217 24701 8251 24735
rect 9597 24701 9631 24735
rect 12725 24701 12759 24735
rect 13093 24701 13127 24735
rect 13369 24701 13403 24735
rect 14933 24701 14967 24735
rect 16129 24701 16163 24735
rect 17509 24701 17543 24735
rect 17601 24701 17635 24735
rect 19533 24701 19567 24735
rect 19809 24701 19843 24735
rect 22293 24701 22327 24735
rect 8585 24633 8619 24667
rect 16405 24633 16439 24667
rect 21833 24633 21867 24667
rect 3341 24565 3375 24599
rect 6745 24565 6779 24599
rect 8953 24565 8987 24599
rect 9229 24565 9263 24599
rect 10057 24565 10091 24599
rect 12909 24565 12943 24599
rect 15025 24565 15059 24599
rect 16681 24565 16715 24599
rect 17969 24565 18003 24599
rect 21281 24565 21315 24599
rect 22661 24565 22695 24599
rect 4261 24361 4295 24395
rect 7389 24361 7423 24395
rect 8217 24361 8251 24395
rect 8401 24361 8435 24395
rect 12633 24361 12667 24395
rect 13001 24361 13035 24395
rect 15656 24361 15690 24395
rect 17233 24361 17267 24395
rect 17785 24361 17819 24395
rect 18705 24361 18739 24395
rect 18889 24361 18923 24395
rect 19349 24361 19383 24395
rect 21097 24361 21131 24395
rect 21373 24361 21407 24395
rect 2053 24293 2087 24327
rect 4629 24293 4663 24327
rect 8493 24293 8527 24327
rect 10793 24293 10827 24327
rect 13093 24293 13127 24327
rect 17693 24293 17727 24327
rect 18613 24293 18647 24327
rect 2513 24225 2547 24259
rect 3525 24225 3559 24259
rect 6929 24225 6963 24259
rect 7941 24225 7975 24259
rect 8585 24225 8619 24259
rect 17877 24225 17911 24259
rect 19257 24225 19291 24259
rect 20453 24225 20487 24259
rect 20545 24225 20579 24259
rect 20729 24225 20763 24259
rect 21189 24225 21223 24259
rect 3065 24157 3099 24191
rect 3249 24157 3283 24191
rect 3341 24157 3375 24191
rect 3433 24157 3467 24191
rect 3617 24157 3651 24191
rect 3893 24157 3927 24191
rect 3985 24157 4019 24191
rect 4353 24157 4387 24191
rect 4721 24157 4755 24191
rect 4813 24157 4847 24191
rect 4997 24157 5031 24191
rect 7849 24157 7883 24191
rect 8309 24157 8343 24191
rect 10241 24157 10275 24191
rect 10425 24157 10459 24191
rect 10517 24157 10551 24191
rect 11069 24157 11103 24191
rect 11162 24157 11196 24191
rect 12449 24157 12483 24191
rect 12633 24157 12667 24191
rect 12725 24157 12759 24191
rect 13277 24157 13311 24191
rect 13369 24157 13403 24191
rect 13553 24157 13587 24191
rect 13645 24157 13679 24191
rect 15393 24157 15427 24191
rect 17233 24157 17267 24191
rect 17509 24157 17543 24191
rect 17601 24157 17635 24191
rect 18429 24157 18463 24191
rect 18613 24157 18647 24191
rect 19625 24157 19659 24191
rect 19717 24157 19751 24191
rect 19993 24157 20027 24191
rect 20269 24157 20303 24191
rect 20821 24157 20855 24191
rect 20913 24157 20947 24191
rect 21097 24157 21131 24191
rect 21465 24157 21499 24191
rect 23305 24157 23339 24191
rect 2053 24089 2087 24123
rect 2605 24089 2639 24123
rect 5089 24089 5123 24123
rect 6653 24089 6687 24123
rect 7573 24089 7607 24123
rect 13001 24089 13035 24123
rect 19073 24089 19107 24123
rect 21189 24089 21223 24123
rect 23029 24089 23063 24123
rect 2789 24021 2823 24055
rect 2881 24021 2915 24055
rect 4537 24021 4571 24055
rect 5181 24021 5215 24055
rect 7205 24021 7239 24055
rect 7373 24021 7407 24055
rect 10333 24021 10367 24055
rect 10977 24021 11011 24055
rect 11437 24021 11471 24055
rect 12817 24021 12851 24055
rect 17141 24021 17175 24055
rect 17417 24021 17451 24055
rect 18873 24021 18907 24055
rect 19533 24021 19567 24055
rect 20085 24021 20119 24055
rect 20545 24021 20579 24055
rect 21557 24021 21591 24055
rect 1961 23817 1995 23851
rect 4169 23817 4203 23851
rect 5825 23817 5859 23851
rect 7757 23817 7791 23851
rect 11253 23817 11287 23851
rect 12817 23817 12851 23851
rect 22293 23817 22327 23851
rect 23029 23817 23063 23851
rect 5549 23749 5583 23783
rect 6929 23749 6963 23783
rect 7665 23749 7699 23783
rect 11897 23749 11931 23783
rect 17877 23749 17911 23783
rect 19165 23749 19199 23783
rect 19625 23749 19659 23783
rect 19901 23749 19935 23783
rect 20085 23749 20119 23783
rect 21281 23749 21315 23783
rect 22001 23749 22035 23783
rect 22201 23749 22235 23783
rect 2145 23681 2179 23715
rect 2421 23681 2455 23715
rect 3065 23681 3099 23715
rect 3617 23681 3651 23715
rect 3709 23681 3743 23715
rect 3893 23681 3927 23715
rect 4077 23681 4111 23715
rect 4813 23681 4847 23715
rect 5089 23681 5123 23715
rect 5365 23681 5399 23715
rect 5641 23681 5675 23715
rect 5917 23681 5951 23715
rect 7113 23681 7147 23715
rect 7573 23681 7607 23715
rect 8401 23681 8435 23715
rect 11069 23681 11103 23715
rect 11161 23681 11195 23715
rect 11805 23681 11839 23715
rect 11989 23681 12023 23715
rect 12357 23681 12391 23715
rect 12571 23681 12605 23715
rect 12725 23681 12759 23715
rect 13093 23681 13127 23715
rect 16681 23681 16715 23715
rect 16957 23681 16991 23715
rect 19257 23681 19291 23715
rect 19441 23681 19475 23715
rect 19533 23681 19567 23715
rect 20361 23681 20395 23715
rect 20453 23681 20487 23715
rect 22477 23681 22511 23715
rect 22569 23681 22603 23715
rect 22753 23681 22787 23715
rect 2329 23613 2363 23647
rect 3433 23613 3467 23647
rect 3801 23613 3835 23647
rect 4905 23613 4939 23647
rect 7941 23613 7975 23647
rect 12265 23613 12299 23647
rect 12817 23613 12851 23647
rect 17049 23613 17083 23647
rect 20177 23613 20211 23647
rect 23029 23613 23063 23647
rect 5365 23545 5399 23579
rect 8769 23545 8803 23579
rect 10885 23545 10919 23579
rect 11529 23545 11563 23579
rect 12173 23545 12207 23579
rect 16773 23545 16807 23579
rect 18153 23545 18187 23579
rect 20269 23545 20303 23579
rect 21005 23545 21039 23579
rect 21833 23545 21867 23579
rect 22845 23545 22879 23579
rect 2513 23477 2547 23511
rect 5273 23477 5307 23511
rect 7297 23477 7331 23511
rect 7389 23477 7423 23511
rect 8861 23477 8895 23511
rect 10701 23477 10735 23511
rect 10977 23477 11011 23511
rect 13001 23477 13035 23511
rect 18337 23477 18371 23511
rect 19717 23477 19751 23511
rect 20821 23477 20855 23511
rect 22017 23477 22051 23511
rect 4537 23273 4571 23307
rect 4721 23273 4755 23307
rect 7757 23273 7791 23307
rect 11069 23273 11103 23307
rect 11253 23273 11287 23307
rect 16037 23273 16071 23307
rect 17325 23273 17359 23307
rect 8585 23205 8619 23239
rect 9137 23205 9171 23239
rect 10977 23205 11011 23239
rect 11437 23205 11471 23239
rect 13001 23205 13035 23239
rect 16773 23205 16807 23239
rect 17969 23205 18003 23239
rect 1685 23137 1719 23171
rect 8769 23137 8803 23171
rect 10425 23137 10459 23171
rect 14105 23137 14139 23171
rect 15853 23137 15887 23171
rect 16957 23137 16991 23171
rect 17509 23137 17543 23171
rect 18337 23137 18371 23171
rect 1409 23069 1443 23103
rect 4169 23069 4203 23103
rect 7389 23069 7423 23103
rect 10241 23069 10275 23103
rect 11713 23069 11747 23103
rect 13215 23069 13249 23103
rect 13369 23069 13403 23103
rect 15945 23069 15979 23103
rect 17417 23069 17451 23103
rect 17601 23069 17635 23103
rect 17785 23069 17819 23103
rect 3433 23001 3467 23035
rect 3801 23001 3835 23035
rect 4353 23001 4387 23035
rect 7757 23001 7791 23035
rect 8309 23001 8343 23035
rect 9505 23001 9539 23035
rect 10149 23001 10183 23035
rect 10609 23001 10643 23035
rect 15577 23001 15611 23035
rect 16497 23001 16531 23035
rect 4553 22933 4587 22967
rect 7941 22933 7975 22967
rect 9045 22933 9079 22967
rect 9873 22933 9907 22967
rect 10057 22933 10091 22967
rect 17049 22933 17083 22967
rect 17877 22933 17911 22967
rect 3617 22729 3651 22763
rect 6377 22729 6411 22763
rect 10149 22729 10183 22763
rect 14355 22729 14389 22763
rect 15577 22729 15611 22763
rect 17417 22729 17451 22763
rect 22461 22729 22495 22763
rect 2145 22661 2179 22695
rect 9321 22661 9355 22695
rect 13461 22661 13495 22695
rect 14565 22661 14599 22695
rect 16957 22661 16991 22695
rect 22661 22661 22695 22695
rect 8125 22593 8159 22627
rect 8769 22593 8803 22627
rect 8861 22593 8895 22627
rect 9045 22593 9079 22627
rect 9137 22593 9171 22627
rect 9413 22593 9447 22627
rect 9597 22593 9631 22627
rect 9781 22593 9815 22627
rect 9965 22593 9999 22627
rect 10425 22593 10459 22627
rect 12173 22593 12207 22627
rect 12265 22593 12299 22627
rect 12357 22593 12391 22627
rect 13185 22593 13219 22627
rect 13277 22593 13311 22627
rect 14105 22593 14139 22627
rect 15485 22593 15519 22627
rect 21097 22593 21131 22627
rect 21190 22593 21224 22627
rect 21833 22593 21867 22627
rect 21926 22593 21960 22627
rect 1869 22525 1903 22559
rect 7849 22525 7883 22559
rect 9689 22525 9723 22559
rect 13829 22525 13863 22559
rect 10333 22457 10367 22491
rect 12541 22457 12575 22491
rect 13461 22457 13495 22491
rect 17233 22457 17267 22491
rect 21465 22457 21499 22491
rect 22201 22457 22235 22491
rect 8953 22389 8987 22423
rect 11989 22389 12023 22423
rect 13553 22389 13587 22423
rect 14013 22389 14047 22423
rect 14197 22389 14231 22423
rect 14381 22389 14415 22423
rect 22293 22389 22327 22423
rect 22477 22389 22511 22423
rect 8309 22185 8343 22219
rect 13093 22185 13127 22219
rect 13277 22185 13311 22219
rect 15761 22185 15795 22219
rect 17141 22185 17175 22219
rect 17969 22185 18003 22219
rect 18153 22185 18187 22219
rect 19901 22185 19935 22219
rect 22385 22185 22419 22219
rect 6377 22117 6411 22151
rect 8217 22117 8251 22151
rect 15301 22117 15335 22151
rect 16221 22117 16255 22151
rect 16865 22117 16899 22151
rect 18061 22117 18095 22151
rect 19441 22117 19475 22151
rect 19993 22117 20027 22151
rect 21281 22117 21315 22151
rect 22569 22117 22603 22151
rect 5917 22049 5951 22083
rect 9229 22049 9263 22083
rect 11989 22049 12023 22083
rect 12357 22049 12391 22083
rect 12817 22049 12851 22083
rect 13737 22049 13771 22083
rect 15209 22049 15243 22083
rect 16129 22049 16163 22083
rect 16589 22049 16623 22083
rect 17325 22049 17359 22083
rect 17693 22049 17727 22083
rect 20453 22049 20487 22083
rect 20913 22049 20947 22083
rect 5641 21981 5675 22015
rect 6193 21981 6227 22015
rect 6469 21981 6503 22015
rect 6561 21981 6595 22015
rect 6745 21981 6779 22015
rect 9321 21981 9355 22015
rect 11437 21981 11471 22015
rect 11529 21981 11563 22015
rect 11797 21981 11831 22015
rect 11897 21981 11931 22015
rect 12081 21981 12115 22015
rect 12265 21981 12299 22015
rect 12449 21981 12483 22015
rect 12633 21981 12667 22015
rect 13829 21981 13863 22015
rect 15117 21981 15151 22015
rect 16037 21981 16071 22015
rect 16313 21981 16347 22015
rect 16497 21981 16531 22015
rect 17141 21981 17175 22015
rect 17417 21981 17451 22015
rect 18245 21981 18279 22015
rect 18429 21981 18463 22015
rect 20361 21981 20395 22015
rect 20821 21981 20855 22015
rect 22017 21981 22051 22015
rect 22845 21981 22879 22015
rect 23121 21981 23155 22015
rect 7849 21913 7883 21947
rect 11713 21913 11747 21947
rect 12909 21913 12943 21947
rect 15669 21913 15703 21947
rect 19717 21913 19751 21947
rect 21557 21913 21591 21947
rect 6561 21845 6595 21879
rect 9689 21845 9723 21879
rect 13109 21845 13143 21879
rect 15025 21845 15059 21879
rect 17049 21845 17083 21879
rect 17601 21845 17635 21879
rect 19257 21845 19291 21879
rect 21097 21845 21131 21879
rect 22385 21845 22419 21879
rect 22661 21845 22695 21879
rect 23029 21845 23063 21879
rect 4813 21641 4847 21675
rect 8309 21641 8343 21675
rect 12265 21641 12299 21675
rect 12357 21641 12391 21675
rect 12541 21641 12575 21675
rect 15577 21641 15611 21675
rect 17969 21641 18003 21675
rect 18613 21641 18647 21675
rect 22017 21641 22051 21675
rect 24409 21641 24443 21675
rect 4353 21573 4387 21607
rect 5089 21573 5123 21607
rect 5457 21573 5491 21607
rect 8769 21573 8803 21607
rect 22937 21573 22971 21607
rect 4905 21505 4939 21539
rect 5641 21505 5675 21539
rect 6009 21505 6043 21539
rect 6193 21505 6227 21539
rect 6929 21505 6963 21539
rect 7941 21505 7975 21539
rect 8401 21505 8435 21539
rect 8555 21505 8589 21539
rect 11529 21505 11563 21539
rect 11713 21505 11747 21539
rect 11805 21505 11839 21539
rect 12081 21505 12115 21539
rect 12538 21505 12572 21539
rect 13001 21505 13035 21539
rect 13369 21505 13403 21539
rect 13461 21505 13495 21539
rect 13645 21505 13679 21539
rect 13737 21505 13771 21539
rect 16129 21505 16163 21539
rect 16681 21505 16715 21539
rect 16773 21505 16807 21539
rect 16957 21505 16991 21539
rect 17049 21505 17083 21539
rect 17141 21505 17175 21539
rect 18245 21505 18279 21539
rect 18337 21505 18371 21539
rect 18705 21505 18739 21539
rect 20361 21505 20395 21539
rect 21005 21505 21039 21539
rect 21649 21505 21683 21539
rect 22109 21505 22143 21539
rect 22385 21505 22419 21539
rect 5825 21437 5859 21471
rect 5917 21437 5951 21471
rect 6837 21437 6871 21471
rect 8033 21437 8067 21471
rect 11897 21437 11931 21471
rect 15117 21437 15151 21471
rect 18429 21437 18463 21471
rect 20085 21437 20119 21471
rect 21925 21437 21959 21471
rect 22661 21437 22695 21471
rect 4353 21369 4387 21403
rect 5733 21369 5767 21403
rect 6009 21369 6043 21403
rect 15485 21369 15519 21403
rect 17417 21369 17451 21403
rect 21281 21369 21315 21403
rect 21833 21369 21867 21403
rect 7297 21301 7331 21335
rect 12909 21301 12943 21335
rect 13185 21301 13219 21335
rect 19809 21301 19843 21335
rect 20269 21301 20303 21335
rect 21189 21301 21223 21335
rect 22293 21301 22327 21335
rect 4997 21097 5031 21131
rect 8309 21097 8343 21131
rect 10149 21097 10183 21131
rect 10793 21097 10827 21131
rect 10977 21097 11011 21131
rect 13553 21097 13587 21131
rect 18245 21097 18279 21131
rect 9965 21029 9999 21063
rect 15577 21029 15611 21063
rect 18061 21029 18095 21063
rect 20361 21029 20395 21063
rect 1409 20961 1443 20995
rect 3157 20961 3191 20995
rect 6745 20961 6779 20995
rect 8401 20961 8435 20995
rect 9689 20961 9723 20995
rect 10333 20961 10367 20995
rect 11069 20961 11103 20995
rect 13369 20961 13403 20995
rect 23581 20961 23615 20995
rect 3479 20893 3513 20927
rect 3617 20893 3651 20927
rect 3801 20893 3835 20927
rect 4169 20893 4203 20927
rect 4629 20893 4663 20927
rect 8585 20893 8619 20927
rect 9597 20893 9631 20927
rect 10517 20893 10551 20927
rect 10977 20893 11011 20927
rect 11253 20893 11287 20927
rect 13277 20893 13311 20927
rect 15209 20893 15243 20927
rect 15363 20893 15397 20927
rect 17417 20893 17451 20927
rect 19257 20893 19291 20927
rect 19441 20893 19475 20927
rect 19717 20893 19751 20927
rect 19993 20893 20027 20927
rect 20147 20893 20181 20927
rect 23029 20893 23063 20927
rect 23121 20893 23155 20927
rect 23213 20893 23247 20927
rect 23397 20893 23431 20927
rect 23489 20893 23523 20927
rect 23673 20893 23707 20927
rect 1685 20825 1719 20859
rect 6469 20825 6503 20859
rect 8309 20825 8343 20859
rect 10057 20825 10091 20859
rect 17785 20825 17819 20859
rect 18889 20825 18923 20859
rect 19073 20825 19107 20859
rect 20545 20825 20579 20859
rect 3249 20757 3283 20791
rect 3893 20757 3927 20791
rect 8769 20757 8803 20791
rect 10701 20757 10735 20791
rect 16129 20757 16163 20791
rect 18705 20757 18739 20791
rect 19901 20757 19935 20791
rect 21833 20757 21867 20791
rect 22753 20757 22787 20791
rect 2329 20553 2363 20587
rect 5457 20553 5491 20587
rect 9873 20553 9907 20587
rect 13645 20553 13679 20587
rect 16681 20553 16715 20587
rect 17233 20553 17267 20587
rect 20545 20553 20579 20587
rect 21189 20553 21223 20587
rect 24777 20553 24811 20587
rect 3249 20485 3283 20519
rect 4997 20485 5031 20519
rect 6745 20485 6779 20519
rect 8185 20485 8219 20519
rect 8401 20485 8435 20519
rect 8677 20485 8711 20519
rect 13277 20485 13311 20519
rect 17141 20485 17175 20519
rect 18613 20485 18647 20519
rect 2513 20417 2547 20451
rect 2605 20417 2639 20451
rect 2789 20417 2823 20451
rect 2881 20417 2915 20451
rect 5641 20417 5675 20451
rect 6009 20417 6043 20451
rect 7021 20417 7055 20451
rect 7573 20417 7607 20451
rect 10241 20417 10275 20451
rect 12817 20417 12851 20451
rect 13461 20417 13495 20451
rect 13737 20417 13771 20451
rect 15577 20417 15611 20451
rect 16037 20417 16071 20451
rect 17508 20417 17542 20451
rect 17601 20417 17635 20451
rect 18061 20417 18095 20451
rect 18797 20417 18831 20451
rect 18889 20417 18923 20451
rect 19625 20417 19659 20451
rect 21005 20417 21039 20451
rect 21281 20417 21315 20451
rect 22477 20417 22511 20451
rect 23029 20417 23063 20451
rect 2973 20349 3007 20383
rect 4721 20349 4755 20383
rect 6745 20349 6779 20383
rect 7481 20349 7515 20383
rect 7941 20349 7975 20383
rect 10333 20349 10367 20383
rect 12909 20349 12943 20383
rect 13185 20349 13219 20383
rect 15669 20349 15703 20383
rect 16497 20349 16531 20383
rect 18153 20349 18187 20383
rect 19717 20349 19751 20383
rect 20821 20349 20855 20383
rect 22569 20349 22603 20383
rect 23305 20349 23339 20383
rect 5365 20281 5399 20315
rect 6929 20281 6963 20315
rect 16313 20281 16347 20315
rect 16773 20281 16807 20315
rect 18613 20281 18647 20315
rect 20913 20281 20947 20315
rect 4813 20213 4847 20247
rect 4997 20213 5031 20247
rect 5641 20213 5675 20247
rect 8033 20213 8067 20247
rect 8217 20213 8251 20247
rect 8585 20213 8619 20247
rect 13829 20213 13863 20247
rect 15945 20213 15979 20247
rect 18429 20213 18463 20247
rect 19993 20213 20027 20247
rect 22109 20213 22143 20247
rect 11897 20009 11931 20043
rect 19257 20009 19291 20043
rect 20085 20009 20119 20043
rect 8217 19941 8251 19975
rect 10149 19941 10183 19975
rect 12173 19941 12207 19975
rect 1409 19873 1443 19907
rect 4905 19873 4939 19907
rect 6377 19873 6411 19907
rect 6653 19873 6687 19907
rect 9321 19873 9355 19907
rect 9689 19873 9723 19907
rect 11805 19873 11839 19907
rect 13645 19873 13679 19907
rect 16497 19873 16531 19907
rect 20177 19873 20211 19907
rect 3433 19805 3467 19839
rect 3617 19805 3651 19839
rect 3801 19805 3835 19839
rect 5365 19805 5399 19839
rect 8953 19805 8987 19839
rect 9137 19805 9171 19839
rect 9781 19805 9815 19839
rect 11989 19805 12023 19839
rect 12081 19805 12115 19839
rect 13921 19805 13955 19839
rect 16129 19805 16163 19839
rect 16222 19805 16256 19839
rect 19809 19805 19843 19839
rect 20085 19805 20119 19839
rect 20361 19805 20395 19839
rect 1685 19737 1719 19771
rect 3249 19737 3283 19771
rect 4997 19737 5031 19771
rect 5457 19737 5491 19771
rect 8585 19737 8619 19771
rect 3157 19669 3191 19703
rect 8125 19669 8159 19703
rect 8401 19669 8435 19703
rect 8493 19669 8527 19703
rect 8769 19669 8803 19703
rect 20545 19669 20579 19703
rect 2789 19465 2823 19499
rect 2881 19465 2915 19499
rect 7113 19465 7147 19499
rect 7297 19465 7331 19499
rect 12281 19465 12315 19499
rect 12449 19465 12483 19499
rect 12741 19465 12775 19499
rect 12909 19465 12943 19499
rect 16221 19465 16255 19499
rect 19533 19465 19567 19499
rect 20729 19465 20763 19499
rect 21833 19465 21867 19499
rect 2605 19397 2639 19431
rect 3617 19397 3651 19431
rect 3801 19397 3835 19431
rect 12081 19397 12115 19431
rect 12541 19397 12575 19431
rect 16037 19397 16071 19431
rect 22017 19397 22051 19431
rect 3065 19329 3099 19363
rect 5641 19329 5675 19363
rect 5825 19329 5859 19363
rect 6009 19329 6043 19363
rect 6193 19329 6227 19363
rect 6745 19329 6779 19363
rect 7849 19329 7883 19363
rect 9873 19329 9907 19363
rect 15853 19329 15887 19363
rect 16129 19329 16163 19363
rect 16221 19329 16255 19363
rect 16405 19329 16439 19363
rect 19901 19329 19935 19363
rect 20637 19329 20671 19363
rect 20913 19329 20947 19363
rect 21281 19329 21315 19363
rect 21465 19329 21499 19363
rect 3157 19261 3191 19295
rect 5733 19261 5767 19295
rect 9965 19261 9999 19295
rect 10241 19261 10275 19295
rect 19809 19261 19843 19295
rect 2237 19193 2271 19227
rect 3617 19193 3651 19227
rect 5089 19193 5123 19227
rect 6193 19193 6227 19227
rect 7665 19193 7699 19227
rect 9137 19193 9171 19227
rect 21649 19193 21683 19227
rect 22385 19193 22419 19227
rect 2605 19125 2639 19159
rect 7297 19125 7331 19159
rect 12265 19125 12299 19159
rect 12725 19125 12759 19159
rect 15669 19125 15703 19159
rect 19717 19125 19751 19159
rect 21097 19125 21131 19159
rect 22017 19125 22051 19159
rect 3939 18921 3973 18955
rect 8493 18921 8527 18955
rect 12449 18921 12483 18955
rect 12725 18921 12759 18955
rect 15209 18921 15243 18955
rect 15853 18921 15887 18955
rect 17785 18921 17819 18955
rect 18898 18921 18932 18955
rect 19257 18921 19291 18955
rect 19717 18921 19751 18955
rect 20269 18921 20303 18955
rect 20913 18921 20947 18955
rect 21741 18921 21775 18955
rect 8953 18853 8987 18887
rect 9597 18853 9631 18887
rect 11897 18853 11931 18887
rect 12541 18853 12575 18887
rect 15393 18853 15427 18887
rect 15485 18853 15519 18887
rect 16037 18853 16071 18887
rect 16681 18853 16715 18887
rect 20453 18853 20487 18887
rect 20545 18853 20579 18887
rect 5733 18785 5767 18819
rect 6561 18785 6595 18819
rect 6837 18785 6871 18819
rect 8677 18785 8711 18819
rect 9229 18785 9263 18819
rect 16221 18785 16255 18819
rect 17417 18785 17451 18819
rect 18337 18785 18371 18819
rect 18613 18785 18647 18819
rect 19349 18785 19383 18819
rect 22293 18785 22327 18819
rect 2973 18717 3007 18751
rect 3157 18717 3191 18751
rect 3249 18717 3283 18751
rect 3341 18717 3375 18751
rect 5365 18717 5399 18751
rect 8401 18717 8435 18751
rect 9321 18717 9355 18751
rect 9597 18717 9631 18751
rect 9781 18717 9815 18751
rect 12081 18717 12115 18751
rect 12173 18717 12207 18751
rect 13093 18717 13127 18751
rect 13369 18717 13403 18751
rect 16313 18717 16347 18751
rect 17509 18717 17543 18751
rect 18245 18717 18279 18751
rect 19533 18717 19567 18751
rect 21373 18717 21407 18751
rect 21557 18717 21591 18751
rect 22017 18717 22051 18751
rect 8677 18649 8711 18683
rect 12725 18649 12759 18683
rect 13553 18649 13587 18683
rect 15025 18649 15059 18683
rect 15225 18649 15259 18683
rect 15853 18649 15887 18683
rect 16773 18649 16807 18683
rect 16957 18649 16991 18683
rect 19073 18649 19107 18683
rect 19257 18649 19291 18683
rect 20085 18649 20119 18683
rect 20301 18649 20335 18683
rect 21189 18649 21223 18683
rect 21465 18649 21499 18683
rect 3617 18581 3651 18615
rect 8309 18581 8343 18615
rect 12265 18581 12299 18615
rect 13185 18581 13219 18615
rect 17141 18581 17175 18615
rect 18705 18581 18739 18615
rect 18873 18581 18907 18615
rect 20913 18581 20947 18615
rect 21097 18581 21131 18615
rect 23765 18581 23799 18615
rect 2973 18377 3007 18411
rect 5365 18377 5399 18411
rect 7297 18377 7331 18411
rect 8125 18377 8159 18411
rect 10425 18377 10459 18411
rect 11713 18377 11747 18411
rect 11897 18377 11931 18411
rect 12909 18377 12943 18411
rect 13277 18377 13311 18411
rect 14473 18377 14507 18411
rect 16957 18377 16991 18411
rect 17049 18377 17083 18411
rect 19533 18377 19567 18411
rect 21833 18377 21867 18411
rect 3709 18309 3743 18343
rect 7481 18309 7515 18343
rect 7665 18309 7699 18343
rect 8953 18309 8987 18343
rect 10977 18309 11011 18343
rect 11161 18309 11195 18343
rect 12449 18309 12483 18343
rect 12665 18309 12699 18343
rect 13553 18309 13587 18343
rect 15945 18309 15979 18343
rect 16681 18309 16715 18343
rect 17509 18309 17543 18343
rect 18061 18309 18095 18343
rect 21373 18309 21407 18343
rect 2881 18241 2915 18275
rect 3065 18241 3099 18275
rect 7849 18241 7883 18275
rect 8677 18241 8711 18275
rect 11345 18241 11379 18275
rect 12265 18241 12299 18275
rect 12909 18241 12943 18275
rect 13093 18241 13127 18275
rect 13185 18239 13219 18273
rect 13461 18241 13495 18275
rect 13645 18241 13679 18275
rect 13737 18241 13771 18275
rect 13921 18241 13955 18275
rect 16865 18241 16899 18275
rect 17325 18241 17359 18275
rect 22201 18241 22235 18275
rect 3433 18173 3467 18207
rect 5917 18173 5951 18207
rect 16221 18173 16255 18207
rect 17785 18173 17819 18207
rect 19901 18173 19935 18207
rect 21649 18173 21683 18207
rect 22293 18173 22327 18207
rect 13737 18105 13771 18139
rect 5181 18037 5215 18071
rect 11897 18037 11931 18071
rect 12633 18037 12667 18071
rect 12817 18037 12851 18071
rect 17233 18037 17267 18071
rect 17693 18037 17727 18071
rect 12081 17833 12115 17867
rect 13921 17833 13955 17867
rect 16865 17833 16899 17867
rect 18797 17833 18831 17867
rect 18981 17833 19015 17867
rect 21005 17833 21039 17867
rect 16681 17765 16715 17799
rect 1409 17697 1443 17731
rect 10609 17697 10643 17731
rect 12173 17697 12207 17731
rect 16313 17697 16347 17731
rect 19257 17697 19291 17731
rect 1777 17629 1811 17663
rect 3203 17629 3237 17663
rect 3801 17629 3835 17663
rect 10333 17629 10367 17663
rect 17233 17629 17267 17663
rect 18613 17629 18647 17663
rect 18889 17629 18923 17663
rect 19073 17629 19107 17663
rect 12449 17561 12483 17595
rect 16037 17561 16071 17595
rect 18429 17561 18463 17595
rect 19533 17561 19567 17595
rect 4445 17493 4479 17527
rect 14565 17493 14599 17527
rect 16865 17493 16899 17527
rect 2237 17289 2271 17323
rect 11345 17289 11379 17323
rect 15837 17289 15871 17323
rect 18521 17289 18555 17323
rect 18705 17289 18739 17323
rect 2743 17221 2777 17255
rect 9873 17221 9907 17255
rect 16037 17221 16071 17255
rect 17049 17221 17083 17255
rect 4169 17153 4203 17187
rect 4537 17153 4571 17187
rect 9597 17153 9631 17187
rect 16773 17153 16807 17187
rect 18889 17153 18923 17187
rect 2329 17085 2363 17119
rect 2513 17085 2547 17119
rect 15669 17017 15703 17051
rect 1869 16949 1903 16983
rect 15853 16949 15887 16983
rect 3203 16745 3237 16779
rect 9229 16745 9263 16779
rect 22293 16677 22327 16711
rect 1409 16609 1443 16643
rect 1777 16609 1811 16643
rect 5365 16609 5399 16643
rect 7159 16609 7193 16643
rect 8125 16609 8159 16643
rect 8217 16609 8251 16643
rect 22201 16609 22235 16643
rect 22385 16609 22419 16643
rect 5733 16541 5767 16575
rect 22477 16541 22511 16575
rect 9321 16473 9355 16507
rect 7665 16405 7699 16439
rect 8033 16405 8067 16439
rect 6377 16201 6411 16235
rect 6745 16201 6779 16235
rect 13921 16201 13955 16235
rect 14289 16201 14323 16235
rect 2789 16133 2823 16167
rect 9275 16133 9309 16167
rect 10517 16133 10551 16167
rect 5825 16065 5859 16099
rect 6837 16065 6871 16099
rect 7481 16065 7515 16099
rect 7849 16065 7883 16099
rect 10425 16065 10459 16099
rect 13553 16065 13587 16099
rect 14013 16065 14047 16099
rect 15025 16065 15059 16099
rect 15669 16065 15703 16099
rect 18429 16065 18463 16099
rect 20729 16065 20763 16099
rect 20913 16065 20947 16099
rect 21005 16065 21039 16099
rect 21189 16065 21223 16099
rect 21373 16065 21407 16099
rect 22845 16065 22879 16099
rect 2881 15997 2915 16031
rect 2973 15997 3007 16031
rect 5917 15997 5951 16031
rect 6009 15997 6043 16031
rect 6929 15997 6963 16031
rect 10609 15997 10643 16031
rect 13645 15997 13679 16031
rect 14289 15997 14323 16031
rect 14749 15997 14783 16031
rect 14841 15997 14875 16031
rect 14933 15997 14967 16031
rect 15577 15997 15611 16031
rect 18705 15997 18739 16031
rect 20177 15997 20211 16031
rect 21649 15997 21683 16031
rect 21833 15997 21867 16031
rect 22385 15997 22419 16031
rect 23121 15997 23155 16031
rect 15209 15929 15243 15963
rect 21005 15929 21039 15963
rect 21465 15929 21499 15963
rect 2421 15861 2455 15895
rect 5457 15861 5491 15895
rect 10057 15861 10091 15895
rect 13553 15861 13587 15895
rect 14105 15861 14139 15895
rect 15945 15861 15979 15895
rect 20913 15861 20947 15895
rect 21373 15861 21407 15895
rect 24593 15861 24627 15895
rect 7113 15657 7147 15691
rect 13185 15657 13219 15691
rect 19809 15657 19843 15691
rect 22937 15657 22971 15691
rect 24593 15657 24627 15691
rect 15393 15589 15427 15623
rect 15761 15589 15795 15623
rect 19717 15589 19751 15623
rect 22661 15589 22695 15623
rect 24041 15589 24075 15623
rect 1685 15521 1719 15555
rect 4445 15521 4479 15555
rect 4997 15521 5031 15555
rect 5365 15521 5399 15555
rect 6791 15521 6825 15555
rect 8125 15521 8159 15555
rect 8309 15521 8343 15555
rect 9137 15521 9171 15555
rect 9781 15521 9815 15555
rect 10149 15521 10183 15555
rect 13277 15521 13311 15555
rect 13553 15521 13587 15555
rect 14749 15521 14783 15555
rect 14933 15521 14967 15555
rect 15945 15521 15979 15555
rect 20913 15521 20947 15555
rect 23489 15521 23523 15555
rect 1409 15453 1443 15487
rect 2053 15453 2087 15487
rect 3479 15453 3513 15487
rect 4261 15453 4295 15487
rect 7021 15453 7055 15487
rect 11805 15453 11839 15487
rect 12909 15453 12943 15487
rect 13645 15453 13679 15487
rect 13742 15453 13776 15487
rect 14105 15453 14139 15487
rect 14289 15453 14323 15487
rect 14565 15453 14599 15487
rect 15025 15453 15059 15487
rect 15485 15453 15519 15487
rect 15577 15453 15611 15487
rect 15761 15453 15795 15487
rect 16313 15453 16347 15487
rect 18245 15453 18279 15487
rect 20177 15453 20211 15487
rect 20335 15453 20369 15487
rect 20637 15453 20671 15487
rect 23397 15453 23431 15487
rect 11989 15385 12023 15419
rect 13369 15385 13403 15419
rect 13553 15385 13587 15419
rect 17877 15385 17911 15419
rect 19349 15385 19383 15419
rect 20453 15385 20487 15419
rect 20545 15385 20579 15419
rect 21189 15385 21223 15419
rect 23765 15385 23799 15419
rect 24501 15385 24535 15419
rect 1593 15317 1627 15351
rect 3801 15317 3835 15351
rect 4169 15317 4203 15351
rect 7665 15317 7699 15351
rect 8033 15317 8067 15351
rect 9229 15317 9263 15351
rect 9321 15317 9355 15351
rect 9689 15317 9723 15351
rect 11575 15317 11609 15351
rect 13001 15317 13035 15351
rect 13093 15317 13127 15351
rect 17739 15317 17773 15351
rect 20821 15317 20855 15351
rect 23305 15317 23339 15351
rect 24225 15317 24259 15351
rect 15577 15113 15611 15147
rect 15761 15113 15795 15147
rect 22477 15113 22511 15147
rect 12541 15045 12575 15079
rect 12817 15045 12851 15079
rect 12909 15045 12943 15079
rect 14657 15045 14691 15079
rect 24593 15045 24627 15079
rect 2789 14977 2823 15011
rect 2881 14977 2915 15011
rect 3249 14977 3283 15011
rect 3617 14977 3651 15011
rect 6745 14977 6779 15011
rect 7481 14977 7515 15011
rect 9781 14977 9815 15011
rect 11207 14977 11241 15011
rect 12265 14977 12299 15011
rect 12449 14977 12483 15011
rect 12633 14977 12667 15011
rect 14933 14977 14967 15011
rect 15209 14977 15243 15011
rect 15393 14977 15427 15011
rect 15485 14977 15519 15011
rect 15669 14977 15703 15011
rect 15945 14977 15979 15011
rect 16037 14977 16071 15011
rect 16313 14977 16347 15011
rect 16405 14977 16439 15011
rect 21465 14977 21499 15011
rect 21649 14977 21683 15011
rect 22109 14977 22143 15011
rect 22293 14977 22327 15011
rect 22661 14977 22695 15011
rect 22937 14977 22971 15011
rect 3065 14909 3099 14943
rect 6837 14909 6871 14943
rect 6929 14909 6963 14943
rect 7849 14909 7883 14943
rect 9413 14909 9447 14943
rect 11713 14909 11747 14943
rect 16957 14909 16991 14943
rect 17325 14909 17359 14943
rect 19257 14909 19291 14943
rect 19533 14909 19567 14943
rect 21281 14909 21315 14943
rect 22753 14909 22787 14943
rect 24869 14909 24903 14943
rect 5043 14841 5077 14875
rect 12081 14841 12115 14875
rect 2421 14773 2455 14807
rect 6377 14773 6411 14807
rect 9275 14773 9309 14807
rect 12173 14773 12207 14807
rect 14749 14773 14783 14807
rect 18751 14773 18785 14807
rect 21649 14773 21683 14807
rect 21925 14773 21959 14807
rect 22661 14773 22695 14807
rect 23121 14773 23155 14807
rect 3203 14569 3237 14603
rect 5043 14569 5077 14603
rect 14289 14569 14323 14603
rect 14473 14569 14507 14603
rect 15485 14569 15519 14603
rect 17325 14569 17359 14603
rect 20453 14569 20487 14603
rect 21741 14569 21775 14603
rect 22753 14569 22787 14603
rect 22937 14569 22971 14603
rect 23305 14569 23339 14603
rect 7757 14501 7791 14535
rect 12081 14501 12115 14535
rect 14841 14501 14875 14535
rect 1777 14433 1811 14467
rect 4721 14433 4755 14467
rect 6469 14433 6503 14467
rect 7481 14433 7515 14467
rect 12449 14433 12483 14467
rect 12909 14433 12943 14467
rect 15209 14433 15243 14467
rect 17785 14433 17819 14467
rect 17877 14433 17911 14467
rect 20913 14433 20947 14467
rect 21005 14433 21039 14467
rect 1409 14365 1443 14399
rect 6837 14365 6871 14399
rect 9229 14365 9263 14399
rect 9597 14365 9631 14399
rect 11529 14365 11563 14399
rect 11897 14365 11931 14399
rect 12357 14365 12391 14399
rect 12817 14365 12851 14399
rect 13001 14365 13035 14399
rect 13093 14365 13127 14399
rect 13369 14365 13403 14399
rect 13461 14365 13495 14399
rect 15025 14365 15059 14399
rect 17693 14365 17727 14399
rect 20821 14365 20855 14399
rect 21741 14365 21775 14399
rect 21925 14365 21959 14399
rect 22201 14365 22235 14399
rect 22385 14365 22419 14399
rect 23213 14365 23247 14399
rect 23397 14365 23431 14399
rect 22891 14331 22925 14365
rect 7297 14297 7331 14331
rect 7941 14297 7975 14331
rect 11713 14297 11747 14331
rect 11805 14297 11839 14331
rect 13277 14297 13311 14331
rect 14105 14297 14139 14331
rect 15301 14297 15335 14331
rect 22017 14297 22051 14331
rect 23121 14297 23155 14331
rect 4169 14229 4203 14263
rect 4537 14229 4571 14263
rect 4629 14229 4663 14263
rect 6929 14229 6963 14263
rect 7389 14229 7423 14263
rect 11023 14229 11057 14263
rect 12725 14229 12759 14263
rect 13645 14229 13679 14263
rect 14305 14229 14339 14263
rect 15501 14229 15535 14263
rect 15669 14229 15703 14263
rect 1593 14025 1627 14059
rect 5871 14025 5905 14059
rect 6837 14025 6871 14059
rect 10057 14025 10091 14059
rect 10425 14025 10459 14059
rect 13730 14025 13764 14059
rect 17509 14025 17543 14059
rect 22845 14025 22879 14059
rect 7665 13957 7699 13991
rect 13829 13957 13863 13991
rect 1409 13889 1443 13923
rect 1961 13889 1995 13923
rect 3755 13889 3789 13923
rect 4445 13889 4479 13923
rect 6745 13889 6779 13923
rect 7573 13889 7607 13923
rect 8125 13889 8159 13923
rect 11897 13889 11931 13923
rect 12173 13889 12207 13923
rect 12633 13889 12667 13923
rect 13544 13879 13578 13913
rect 13645 13889 13679 13923
rect 17325 13889 17359 13923
rect 17509 13889 17543 13923
rect 22017 13889 22051 13923
rect 22201 13889 22235 13923
rect 22477 13889 22511 13923
rect 22569 13889 22603 13923
rect 23121 13889 23155 13923
rect 2329 13821 2363 13855
rect 4077 13821 4111 13855
rect 7021 13821 7055 13855
rect 7757 13821 7791 13855
rect 8493 13821 8527 13855
rect 10517 13821 10551 13855
rect 10701 13821 10735 13855
rect 11989 13821 12023 13855
rect 12081 13821 12115 13855
rect 12357 13821 12391 13855
rect 12725 13821 12759 13855
rect 17877 13821 17911 13855
rect 22753 13821 22787 13855
rect 22845 13821 22879 13855
rect 13001 13753 13035 13787
rect 18153 13753 18187 13787
rect 23029 13753 23063 13787
rect 6377 13685 6411 13719
rect 7205 13685 7239 13719
rect 9919 13685 9953 13719
rect 18337 13685 18371 13719
rect 22201 13685 22235 13719
rect 22385 13685 22419 13719
rect 22661 13685 22695 13719
rect 2789 13481 2823 13515
rect 8953 13481 8987 13515
rect 12081 13481 12115 13515
rect 14289 13481 14323 13515
rect 21833 13481 21867 13515
rect 22385 13481 22419 13515
rect 22569 13481 22603 13515
rect 22937 13481 22971 13515
rect 23121 13481 23155 13515
rect 23673 13481 23707 13515
rect 8631 13413 8665 13447
rect 11529 13413 11563 13447
rect 21281 13413 21315 13447
rect 22017 13413 22051 13447
rect 3249 13345 3283 13379
rect 3341 13345 3375 13379
rect 4905 13345 4939 13379
rect 5273 13345 5307 13379
rect 6837 13345 6871 13379
rect 7205 13345 7239 13379
rect 9413 13345 9447 13379
rect 9597 13345 9631 13379
rect 17969 13345 18003 13379
rect 18705 13345 18739 13379
rect 23397 13345 23431 13379
rect 3157 13277 3191 13311
rect 11805 13277 11839 13311
rect 15761 13277 15795 13311
rect 16037 13277 16071 13311
rect 16773 13277 16807 13311
rect 17141 13277 17175 13311
rect 17417 13277 17451 13311
rect 17693 13277 17727 13311
rect 17785 13277 17819 13311
rect 17877 13277 17911 13311
rect 18245 13277 18279 13311
rect 18521 13277 18555 13311
rect 21005 13277 21039 13311
rect 21097 13277 21131 13311
rect 21281 13277 21315 13311
rect 21557 13277 21591 13311
rect 21741 13277 21775 13311
rect 22293 13277 22327 13311
rect 22853 13287 22887 13321
rect 23029 13277 23063 13311
rect 23305 13277 23339 13311
rect 23489 13277 23523 13311
rect 23673 13277 23707 13311
rect 23857 13277 23891 13311
rect 23949 13277 23983 13311
rect 24133 13277 24167 13311
rect 24593 13277 24627 13311
rect 11897 13209 11931 13243
rect 14105 13209 14139 13243
rect 14310 13209 14344 13243
rect 22553 13209 22587 13243
rect 22707 13209 22741 13243
rect 6699 13141 6733 13175
rect 9321 13141 9355 13175
rect 11713 13141 11747 13175
rect 14473 13141 14507 13175
rect 15577 13141 15611 13175
rect 15945 13141 15979 13175
rect 16221 13141 16255 13175
rect 16957 13141 16991 13175
rect 17325 13141 17359 13175
rect 18153 13141 18187 13175
rect 18337 13141 18371 13175
rect 21373 13141 21407 13175
rect 24041 13141 24075 13175
rect 24777 13141 24811 13175
rect 3709 12937 3743 12971
rect 5181 12937 5215 12971
rect 8171 12937 8205 12971
rect 21373 12937 21407 12971
rect 21557 12937 21591 12971
rect 21833 12937 21867 12971
rect 22477 12937 22511 12971
rect 24133 12937 24167 12971
rect 17141 12869 17175 12903
rect 17601 12869 17635 12903
rect 19533 12869 19567 12903
rect 19625 12869 19659 12903
rect 22661 12869 22695 12903
rect 23581 12869 23615 12903
rect 24409 12869 24443 12903
rect 3801 12801 3835 12835
rect 6377 12801 6411 12835
rect 6745 12801 6779 12835
rect 9505 12801 9539 12835
rect 12081 12801 12115 12835
rect 12265 12801 12299 12835
rect 15025 12801 15059 12835
rect 16451 12801 16485 12835
rect 16681 12801 16715 12835
rect 16865 12801 16899 12835
rect 16957 12801 16991 12835
rect 17233 12801 17267 12835
rect 17325 12801 17359 12835
rect 17785 12801 17819 12835
rect 18245 12801 18279 12835
rect 18889 12801 18923 12835
rect 19349 12801 19383 12835
rect 19717 12801 19751 12835
rect 21189 12801 21223 12835
rect 21649 12801 21683 12835
rect 22569 12801 22603 12835
rect 23029 12801 23063 12835
rect 23121 12801 23155 12835
rect 23305 12801 23339 12835
rect 24225 12801 24259 12835
rect 24317 12801 24351 12835
rect 24501 12801 24535 12835
rect 3617 12733 3651 12767
rect 5273 12733 5307 12767
rect 5365 12733 5399 12767
rect 9597 12733 9631 12767
rect 9781 12733 9815 12767
rect 14657 12733 14691 12767
rect 18337 12733 18371 12767
rect 18613 12733 18647 12767
rect 18797 12733 18831 12767
rect 21281 12733 21315 12767
rect 22109 12733 22143 12767
rect 16773 12665 16807 12699
rect 19257 12665 19291 12699
rect 22201 12665 22235 12699
rect 22937 12665 22971 12699
rect 23949 12665 23983 12699
rect 4169 12597 4203 12631
rect 4813 12597 4847 12631
rect 9137 12597 9171 12631
rect 12173 12597 12207 12631
rect 17509 12597 17543 12631
rect 17969 12597 18003 12631
rect 19901 12597 19935 12631
rect 21005 12597 21039 12631
rect 22293 12597 22327 12631
rect 22845 12597 22879 12631
rect 23397 12597 23431 12631
rect 23581 12597 23615 12631
rect 10747 12393 10781 12427
rect 16635 12393 16669 12427
rect 17417 12393 17451 12427
rect 17601 12393 17635 12427
rect 18337 12393 18371 12427
rect 19441 12393 19475 12427
rect 22385 12393 22419 12427
rect 22734 12393 22768 12427
rect 24225 12393 24259 12427
rect 11713 12325 11747 12359
rect 13093 12325 13127 12359
rect 17785 12325 17819 12359
rect 18153 12325 18187 12359
rect 21557 12325 21591 12359
rect 1409 12257 1443 12291
rect 3801 12257 3835 12291
rect 9321 12257 9355 12291
rect 11161 12257 11195 12291
rect 12265 12257 12299 12291
rect 15209 12257 15243 12291
rect 19809 12257 19843 12291
rect 21005 12257 21039 12291
rect 22017 12257 22051 12291
rect 22109 12257 22143 12291
rect 22477 12257 22511 12291
rect 3433 12189 3467 12223
rect 4169 12189 4203 12223
rect 8953 12189 8987 12223
rect 11345 12189 11379 12223
rect 11437 12189 11471 12223
rect 11529 12189 11563 12223
rect 12173 12189 12207 12223
rect 12633 12189 12667 12223
rect 12817 12189 12851 12223
rect 13369 12189 13403 12223
rect 14841 12189 14875 12223
rect 17693 12189 17727 12223
rect 17969 12189 18003 12223
rect 18245 12189 18279 12223
rect 18429 12189 18463 12223
rect 18521 12189 18555 12223
rect 18705 12189 18739 12223
rect 18889 12189 18923 12223
rect 19625 12189 19659 12223
rect 19901 12189 19935 12223
rect 19993 12189 20027 12223
rect 20177 12189 20211 12223
rect 20637 12189 20671 12223
rect 20913 12189 20947 12223
rect 21189 12189 21223 12223
rect 21373 12189 21407 12223
rect 21465 12189 21499 12223
rect 21741 12189 21775 12223
rect 21925 12189 21959 12223
rect 22201 12189 22235 12223
rect 1685 12121 1719 12155
rect 13553 12121 13587 12155
rect 17233 12121 17267 12155
rect 17433 12121 17467 12155
rect 18613 12121 18647 12155
rect 3157 12053 3191 12087
rect 3341 12053 3375 12087
rect 5595 12053 5629 12087
rect 12541 12053 12575 12087
rect 12909 12053 12943 12087
rect 13737 12053 13771 12087
rect 20453 12053 20487 12087
rect 20821 12053 20855 12087
rect 2145 11849 2179 11883
rect 6837 11849 6871 11883
rect 12265 11849 12299 11883
rect 18245 11849 18279 11883
rect 18613 11849 18647 11883
rect 19073 11849 19107 11883
rect 19533 11849 19567 11883
rect 22385 11849 22419 11883
rect 1961 11781 1995 11815
rect 2513 11781 2547 11815
rect 2881 11781 2915 11815
rect 6147 11781 6181 11815
rect 11023 11781 11057 11815
rect 11805 11781 11839 11815
rect 11897 11781 11931 11815
rect 18705 11781 18739 11815
rect 18905 11781 18939 11815
rect 1685 11713 1719 11747
rect 1777 11713 1811 11747
rect 2053 11713 2087 11747
rect 2329 11713 2363 11747
rect 2605 11713 2639 11747
rect 4721 11713 4755 11747
rect 6745 11713 6779 11747
rect 8125 11713 8159 11747
rect 9229 11713 9263 11747
rect 11621 11713 11655 11747
rect 11994 11713 12028 11747
rect 12173 11713 12207 11747
rect 12357 11713 12391 11747
rect 12633 11713 12667 11747
rect 13185 11713 13219 11747
rect 13369 11713 13403 11747
rect 13921 11713 13955 11747
rect 18153 11713 18187 11747
rect 18429 11713 18463 11747
rect 19349 11713 19383 11747
rect 19993 11713 20027 11747
rect 20085 11713 20119 11747
rect 20269 11713 20303 11747
rect 20361 11713 20395 11747
rect 21925 11713 21959 11747
rect 22017 11713 22051 11747
rect 22201 11713 22235 11747
rect 3433 11645 3467 11679
rect 4169 11645 4203 11679
rect 4353 11645 4387 11679
rect 6929 11645 6963 11679
rect 8217 11645 8251 11679
rect 8309 11645 8343 11679
rect 9597 11645 9631 11679
rect 11805 11645 11839 11679
rect 12725 11645 12759 11679
rect 13277 11645 13311 11679
rect 13737 11645 13771 11679
rect 19165 11645 19199 11679
rect 3617 11577 3651 11611
rect 13001 11577 13035 11611
rect 1501 11509 1535 11543
rect 1777 11509 1811 11543
rect 6377 11509 6411 11543
rect 7757 11509 7791 11543
rect 14105 11509 14139 11543
rect 18889 11509 18923 11543
rect 20545 11509 20579 11543
rect 4261 11305 4295 11339
rect 6791 11305 6825 11339
rect 8677 11305 8711 11339
rect 9781 11305 9815 11339
rect 19993 11305 20027 11339
rect 20729 11305 20763 11339
rect 21925 11305 21959 11339
rect 10609 11237 10643 11271
rect 12725 11237 12759 11271
rect 20821 11237 20855 11271
rect 21833 11237 21867 11271
rect 1685 11169 1719 11203
rect 5365 11169 5399 11203
rect 6929 11169 6963 11203
rect 7297 11169 7331 11203
rect 10333 11169 10367 11203
rect 15209 11169 15243 11203
rect 17141 11169 17175 11203
rect 20637 11169 20671 11203
rect 21373 11169 21407 11203
rect 21649 11169 21683 11203
rect 1409 11101 1443 11135
rect 1593 11101 1627 11135
rect 4077 11101 4111 11135
rect 4997 11101 5031 11135
rect 10149 11101 10183 11135
rect 13001 11101 13035 11135
rect 13277 11101 13311 11135
rect 13553 11101 13587 11135
rect 13645 11101 13679 11135
rect 13921 11101 13955 11135
rect 15577 11101 15611 11135
rect 20177 11101 20211 11135
rect 20269 11101 20303 11135
rect 20361 11101 20395 11135
rect 20453 11101 20487 11135
rect 20913 11101 20947 11135
rect 21465 11101 21499 11135
rect 21557 11101 21591 11135
rect 22109 11101 22143 11135
rect 22201 11101 22235 11135
rect 22385 11101 22419 11135
rect 22477 11101 22511 11135
rect 1501 11033 1535 11067
rect 1961 11033 1995 11067
rect 4445 11033 4479 11067
rect 4629 11033 4663 11067
rect 10241 11033 10275 11067
rect 10793 11033 10827 11067
rect 13093 11033 13127 11067
rect 13737 11033 13771 11067
rect 17003 11033 17037 11067
rect 18889 11033 18923 11067
rect 3433 10965 3467 10999
rect 12909 10965 12943 10999
rect 13369 10965 13403 10999
rect 9183 10761 9217 10795
rect 14289 10761 14323 10795
rect 17141 10761 17175 10795
rect 17601 10761 17635 10795
rect 21557 10761 21591 10795
rect 22293 10761 22327 10795
rect 5457 10693 5491 10727
rect 13645 10693 13679 10727
rect 14197 10693 14231 10727
rect 2789 10625 2823 10659
rect 3065 10625 3099 10659
rect 7389 10625 7423 10659
rect 13276 10625 13310 10659
rect 13369 10625 13403 10659
rect 13461 10625 13495 10659
rect 13737 10625 13771 10659
rect 13829 10625 13863 10659
rect 14105 10625 14139 10659
rect 15945 10625 15979 10659
rect 17509 10625 17543 10659
rect 21097 10625 21131 10659
rect 21281 10625 21315 10659
rect 22477 10625 22511 10659
rect 22661 10625 22695 10659
rect 2973 10557 3007 10591
rect 7757 10557 7791 10591
rect 14473 10557 14507 10591
rect 17693 10557 17727 10591
rect 21557 10557 21591 10591
rect 3065 10421 3099 10455
rect 3249 10421 3283 10455
rect 4169 10421 4203 10455
rect 13185 10421 13219 10455
rect 14013 10421 14047 10455
rect 14381 10421 14415 10455
rect 21373 10421 21407 10455
rect 4537 10217 4571 10251
rect 17923 10217 17957 10251
rect 19901 10217 19935 10251
rect 21741 10217 21775 10251
rect 3157 10149 3191 10183
rect 3249 10149 3283 10183
rect 3985 10149 4019 10183
rect 6101 10149 6135 10183
rect 13921 10149 13955 10183
rect 20361 10149 20395 10183
rect 22293 10149 22327 10183
rect 2421 10081 2455 10115
rect 4353 10081 4387 10115
rect 7021 10081 7055 10115
rect 10057 10081 10091 10115
rect 10149 10081 10183 10115
rect 10885 10081 10919 10115
rect 10977 10081 11011 10115
rect 13461 10081 13495 10115
rect 16129 10081 16163 10115
rect 18521 10081 18555 10115
rect 18613 10081 18647 10115
rect 19349 10081 19383 10115
rect 22569 10081 22603 10115
rect 2329 10013 2363 10047
rect 3065 10013 3099 10047
rect 3341 10013 3375 10047
rect 4169 10013 4203 10047
rect 4610 10023 4644 10057
rect 4727 10013 4761 10047
rect 4905 10013 4939 10047
rect 6285 10013 6319 10047
rect 8769 10013 8803 10047
rect 13093 10013 13127 10047
rect 13277 10013 13311 10047
rect 13553 10013 13587 10047
rect 14105 10013 14139 10047
rect 14289 10013 14323 10047
rect 14381 10013 14415 10047
rect 14473 10013 14507 10047
rect 14749 10013 14783 10047
rect 15117 10013 15151 10047
rect 15761 10013 15795 10047
rect 16497 10013 16531 10047
rect 19257 10013 19291 10047
rect 19441 10013 19475 10047
rect 19533 10013 19567 10047
rect 19717 10013 19751 10047
rect 20085 10013 20119 10047
rect 20361 10013 20395 10047
rect 20453 10013 20487 10047
rect 22661 10013 22695 10047
rect 6469 9945 6503 9979
rect 13185 9945 13219 9979
rect 14611 9945 14645 9979
rect 18429 9945 18463 9979
rect 2145 9877 2179 9911
rect 2789 9877 2823 9911
rect 2881 9877 2915 9911
rect 4353 9877 4387 9911
rect 4813 9877 4847 9911
rect 9597 9877 9631 9911
rect 9965 9877 9999 9911
rect 10425 9877 10459 9911
rect 10793 9877 10827 9911
rect 18061 9877 18095 9911
rect 20177 9877 20211 9911
rect 4445 9673 4479 9707
rect 8401 9673 8435 9707
rect 15669 9673 15703 9707
rect 16681 9673 16715 9707
rect 17141 9673 17175 9707
rect 19717 9673 19751 9707
rect 2881 9605 2915 9639
rect 3617 9605 3651 9639
rect 4629 9605 4663 9639
rect 11989 9605 12023 9639
rect 19303 9605 19337 9639
rect 19993 9605 20027 9639
rect 20637 9605 20671 9639
rect 21373 9605 21407 9639
rect 3341 9537 3375 9571
rect 3801 9537 3835 9571
rect 4077 9537 4111 9571
rect 4261 9537 4295 9571
rect 4353 9537 4387 9571
rect 4537 9537 4571 9571
rect 4905 9537 4939 9571
rect 5181 9537 5215 9571
rect 5365 9537 5399 9571
rect 5917 9537 5951 9571
rect 6561 9537 6595 9571
rect 7021 9537 7055 9571
rect 7205 9537 7239 9571
rect 9505 9537 9539 9571
rect 11299 9537 11333 9571
rect 11897 9537 11931 9571
rect 13553 9537 13587 9571
rect 15610 9537 15644 9571
rect 17049 9537 17083 9571
rect 17509 9537 17543 9571
rect 19625 9537 19659 9571
rect 19809 9537 19843 9571
rect 19901 9537 19935 9571
rect 20085 9537 20119 9571
rect 20361 9537 20395 9571
rect 20729 9537 20763 9571
rect 20913 9537 20947 9571
rect 21189 9537 21223 9571
rect 21833 9537 21867 9571
rect 3249 9469 3283 9503
rect 4721 9469 4755 9503
rect 6469 9469 6503 9503
rect 7389 9469 7423 9503
rect 8493 9469 8527 9503
rect 8585 9469 8619 9503
rect 9873 9469 9907 9503
rect 12081 9469 12115 9503
rect 13921 9469 13955 9503
rect 15347 9469 15381 9503
rect 16129 9469 16163 9503
rect 17233 9469 17267 9503
rect 17877 9469 17911 9503
rect 20637 9469 20671 9503
rect 21925 9469 21959 9503
rect 8033 9401 8067 9435
rect 11529 9401 11563 9435
rect 20453 9401 20487 9435
rect 22201 9401 22235 9435
rect 3249 9333 3283 9367
rect 3525 9333 3559 9367
rect 4629 9333 4663 9367
rect 5089 9333 5123 9367
rect 6837 9333 6871 9367
rect 15485 9333 15519 9367
rect 16037 9333 16071 9367
rect 21833 9333 21867 9367
rect 6101 9129 6135 9163
rect 6285 9129 6319 9163
rect 12035 9129 12069 9163
rect 16819 9129 16853 9163
rect 20729 9129 20763 9163
rect 4997 9061 5031 9095
rect 12817 9061 12851 9095
rect 19809 9061 19843 9095
rect 21373 9061 21407 9095
rect 3525 8993 3559 9027
rect 3801 8993 3835 9027
rect 4629 8993 4663 9027
rect 6561 8993 6595 9027
rect 8309 8993 8343 9027
rect 9413 8993 9447 9027
rect 9505 8993 9539 9027
rect 10609 8993 10643 9027
rect 15025 8993 15059 9027
rect 19349 8993 19383 9027
rect 19901 8993 19935 9027
rect 21097 8993 21131 9027
rect 21833 8993 21867 9027
rect 2881 8925 2915 8959
rect 3157 8925 3191 8959
rect 3341 8925 3375 8959
rect 3433 8925 3467 8959
rect 3617 8925 3651 8959
rect 4169 8925 4203 8959
rect 4905 8925 4939 8959
rect 5089 8925 5123 8959
rect 5181 8925 5215 8959
rect 5365 8925 5399 8959
rect 5457 8925 5491 8959
rect 5549 8925 5583 8959
rect 10241 8925 10275 8959
rect 12265 8925 12299 8959
rect 12541 8925 12575 8959
rect 12633 8925 12667 8959
rect 13185 8925 13219 8959
rect 13277 8925 13311 8959
rect 13461 8925 13495 8959
rect 15393 8925 15427 8959
rect 16957 8925 16991 8959
rect 17325 8925 17359 8959
rect 19441 8925 19475 8959
rect 20085 8925 20119 8959
rect 20545 8925 20579 8959
rect 21005 8925 21039 8959
rect 21465 8925 21499 8959
rect 21558 8925 21592 8959
rect 4261 8857 4295 8891
rect 4445 8857 4479 8891
rect 5917 8857 5951 8891
rect 8033 8857 8067 8891
rect 12449 8857 12483 8891
rect 12909 8857 12943 8891
rect 13093 8857 13127 8891
rect 20361 8857 20395 8891
rect 2697 8789 2731 8823
rect 3801 8789 3835 8823
rect 3985 8789 4019 8823
rect 4077 8789 4111 8823
rect 5825 8789 5859 8823
rect 6117 8789 6151 8823
rect 8953 8789 8987 8823
rect 9321 8789 9355 8823
rect 13185 8789 13219 8823
rect 13645 8789 13679 8823
rect 18751 8789 18785 8823
rect 20269 8789 20303 8823
rect 3433 8585 3467 8619
rect 4445 8585 4479 8619
rect 5273 8585 5307 8619
rect 12725 8585 12759 8619
rect 17049 8585 17083 8619
rect 17417 8585 17451 8619
rect 20269 8585 20303 8619
rect 3893 8517 3927 8551
rect 8861 8517 8895 8551
rect 17509 8517 17543 8551
rect 2513 8449 2547 8483
rect 2789 8449 2823 8483
rect 2881 8449 2915 8483
rect 3065 8449 3099 8483
rect 3157 8449 3191 8483
rect 3249 8449 3283 8483
rect 3709 8449 3743 8483
rect 3805 8449 3839 8483
rect 4077 8449 4111 8483
rect 4353 8449 4387 8483
rect 4813 8449 4847 8483
rect 5181 8449 5215 8483
rect 5365 8449 5399 8483
rect 5641 8449 5675 8483
rect 7021 8449 7055 8483
rect 7389 8449 7423 8483
rect 8953 8449 8987 8483
rect 9321 8449 9355 8483
rect 10793 8449 10827 8483
rect 12541 8449 12575 8483
rect 13461 8449 13495 8483
rect 20453 8449 20487 8483
rect 20637 8449 20671 8483
rect 4721 8381 4755 8415
rect 12357 8381 12391 8415
rect 17601 8381 17635 8415
rect 2237 8313 2271 8347
rect 3525 8313 3559 8347
rect 2605 8245 2639 8279
rect 4261 8245 4295 8279
rect 4813 8245 4847 8279
rect 5733 8245 5767 8279
rect 13645 8245 13679 8279
rect 2697 8041 2731 8075
rect 2881 8041 2915 8075
rect 3341 8041 3375 8075
rect 3617 8041 3651 8075
rect 12357 8041 12391 8075
rect 16083 8041 16117 8075
rect 2973 7973 3007 8007
rect 6469 7973 6503 8007
rect 12725 7973 12759 8007
rect 13829 7973 13863 8007
rect 3249 7905 3283 7939
rect 6009 7905 6043 7939
rect 7481 7905 7515 7939
rect 13001 7905 13035 7939
rect 13185 7905 13219 7939
rect 14289 7905 14323 7939
rect 3341 7837 3375 7871
rect 3433 7837 3467 7871
rect 3617 7837 3651 7871
rect 3985 7837 4019 7871
rect 4077 7837 4111 7871
rect 4261 7837 4295 7871
rect 4353 7837 4387 7871
rect 6377 7837 6411 7871
rect 6561 7837 6595 7871
rect 6653 7837 6687 7871
rect 6837 7837 6871 7871
rect 6929 7837 6963 7871
rect 7113 7837 7147 7871
rect 7573 7837 7607 7871
rect 12357 7837 12391 7871
rect 12449 7837 12483 7871
rect 13093 7837 13127 7871
rect 13277 7837 13311 7871
rect 13553 7837 13587 7871
rect 13645 7837 13679 7871
rect 14657 7837 14691 7871
rect 18521 7837 18555 7871
rect 2513 7769 2547 7803
rect 3801 7769 3835 7803
rect 13829 7769 13863 7803
rect 2723 7701 2757 7735
rect 5457 7701 5491 7735
rect 6193 7701 6227 7735
rect 7297 7701 7331 7735
rect 13461 7701 13495 7735
rect 18797 7701 18831 7735
rect 2881 7497 2915 7531
rect 4169 7497 4203 7531
rect 4905 7497 4939 7531
rect 6929 7497 6963 7531
rect 9045 7497 9079 7531
rect 10241 7497 10275 7531
rect 11989 7497 12023 7531
rect 14289 7497 14323 7531
rect 19671 7497 19705 7531
rect 5089 7429 5123 7463
rect 6745 7429 6779 7463
rect 14933 7429 14967 7463
rect 17233 7429 17267 7463
rect 3156 7361 3190 7395
rect 3249 7361 3283 7395
rect 4077 7361 4111 7395
rect 4261 7361 4295 7395
rect 4353 7361 4387 7395
rect 4537 7361 4571 7395
rect 4629 7361 4663 7395
rect 4813 7361 4847 7395
rect 5273 7361 5307 7395
rect 5549 7361 5583 7395
rect 5825 7361 5859 7395
rect 5917 7361 5951 7395
rect 6561 7361 6595 7395
rect 8953 7361 8987 7395
rect 10149 7361 10183 7395
rect 10793 7361 10827 7395
rect 11713 7361 11747 7395
rect 11805 7361 11839 7395
rect 12081 7361 12115 7395
rect 12265 7361 12299 7395
rect 12541 7361 12575 7395
rect 13185 7361 13219 7395
rect 14565 7361 14599 7395
rect 16957 7361 16991 7395
rect 17141 7361 17175 7395
rect 17325 7361 17359 7395
rect 18245 7361 18279 7395
rect 9229 7293 9263 7327
rect 10333 7293 10367 7327
rect 11989 7293 12023 7327
rect 12725 7293 12759 7327
rect 13093 7293 13127 7327
rect 14473 7293 14507 7327
rect 14841 7293 14875 7327
rect 17877 7293 17911 7327
rect 4445 7225 4479 7259
rect 13553 7225 13587 7259
rect 17509 7225 17543 7259
rect 4813 7157 4847 7191
rect 5641 7157 5675 7191
rect 6009 7157 6043 7191
rect 8585 7157 8619 7191
rect 9781 7157 9815 7191
rect 10701 7157 10735 7191
rect 3617 6953 3651 6987
rect 4629 6953 4663 6987
rect 4905 6953 4939 6987
rect 5549 6953 5583 6987
rect 11023 6953 11057 6987
rect 12081 6953 12115 6987
rect 12725 6953 12759 6987
rect 16405 6953 16439 6987
rect 21051 6953 21085 6987
rect 3065 6885 3099 6919
rect 12633 6885 12667 6919
rect 2513 6817 2547 6851
rect 2973 6817 3007 6851
rect 4721 6817 4755 6851
rect 5273 6817 5307 6851
rect 7757 6817 7791 6851
rect 8493 6817 8527 6851
rect 8677 6817 8711 6851
rect 9597 6817 9631 6851
rect 16037 6817 16071 6851
rect 18061 6817 18095 6851
rect 19257 6817 19291 6851
rect 2329 6749 2363 6783
rect 3249 6749 3283 6783
rect 3433 6749 3467 6783
rect 3617 6749 3651 6783
rect 4077 6749 4111 6783
rect 4353 6749 4387 6783
rect 4445 6749 4479 6783
rect 4537 6749 4571 6783
rect 5089 6749 5123 6783
rect 5640 6749 5674 6783
rect 5733 6749 5767 6783
rect 5825 6749 5859 6783
rect 5918 6749 5952 6783
rect 7665 6749 7699 6783
rect 9229 6749 9263 6783
rect 12244 6743 12278 6777
rect 12360 6749 12394 6783
rect 12449 6749 12483 6783
rect 12633 6749 12667 6783
rect 12909 6749 12943 6783
rect 13001 6749 13035 6783
rect 16129 6749 16163 6783
rect 17417 6749 17451 6783
rect 19073 6749 19107 6783
rect 19625 6749 19659 6783
rect 2421 6681 2455 6715
rect 4261 6681 4295 6715
rect 11529 6681 11563 6715
rect 11713 6681 11747 6715
rect 11805 6681 11839 6715
rect 11897 6681 11931 6715
rect 15669 6681 15703 6715
rect 15853 6681 15887 6715
rect 16221 6681 16255 6715
rect 16405 6681 16439 6715
rect 18429 6681 18463 6715
rect 1961 6613 1995 6647
rect 3893 6613 3927 6647
rect 6193 6613 6227 6647
rect 7205 6613 7239 6647
rect 7573 6613 7607 6647
rect 8033 6613 8067 6647
rect 8401 6613 8435 6647
rect 17325 6613 17359 6647
rect 17509 6613 17543 6647
rect 3157 6409 3191 6443
rect 3617 6409 3651 6443
rect 6745 6409 6779 6443
rect 6837 6409 6871 6443
rect 10517 6409 10551 6443
rect 13185 6409 13219 6443
rect 14381 6409 14415 6443
rect 20545 6409 20579 6443
rect 21005 6409 21039 6443
rect 21557 6409 21591 6443
rect 1685 6341 1719 6375
rect 9597 6341 9631 6375
rect 12541 6341 12575 6375
rect 12817 6341 12851 6375
rect 13017 6341 13051 6375
rect 14197 6341 14231 6375
rect 15025 6341 15059 6375
rect 16359 6341 16393 6375
rect 7757 6273 7791 6307
rect 8125 6273 8159 6307
rect 10425 6273 10459 6307
rect 11529 6273 11563 6307
rect 11713 6273 11747 6307
rect 12440 6279 12474 6313
rect 12725 6273 12759 6307
rect 13461 6273 13495 6307
rect 13645 6273 13679 6307
rect 13737 6273 13771 6307
rect 14013 6273 14047 6307
rect 14841 6273 14875 6307
rect 14933 6273 14967 6307
rect 15209 6273 15243 6307
rect 15577 6273 15611 6307
rect 15761 6273 15795 6307
rect 16037 6273 16071 6307
rect 16129 6273 16163 6307
rect 16221 6273 16255 6307
rect 16497 6273 16531 6307
rect 16681 6273 16715 6307
rect 20913 6273 20947 6307
rect 21373 6273 21407 6307
rect 1409 6205 1443 6239
rect 3709 6205 3743 6239
rect 3893 6205 3927 6239
rect 6929 6205 6963 6239
rect 17049 6205 17083 6239
rect 20085 6205 20119 6239
rect 20453 6205 20487 6239
rect 21097 6205 21131 6239
rect 12725 6137 12759 6171
rect 14657 6137 14691 6171
rect 15577 6137 15611 6171
rect 15853 6137 15887 6171
rect 18475 6137 18509 6171
rect 18659 6137 18693 6171
rect 3249 6069 3283 6103
rect 6377 6069 6411 6103
rect 11621 6069 11655 6103
rect 13001 6069 13035 6103
rect 13277 6069 13311 6103
rect 1764 5865 1798 5899
rect 5089 5865 5123 5899
rect 8677 5865 8711 5899
rect 13277 5865 13311 5899
rect 16313 5865 16347 5899
rect 17141 5865 17175 5899
rect 12265 5797 12299 5831
rect 19073 5797 19107 5831
rect 1501 5729 1535 5763
rect 6561 5729 6595 5763
rect 6837 5729 6871 5763
rect 6929 5729 6963 5763
rect 10241 5729 10275 5763
rect 11805 5729 11839 5763
rect 12173 5729 12207 5763
rect 15669 5729 15703 5763
rect 16681 5729 16715 5763
rect 18521 5729 18555 5763
rect 20729 5729 20763 5763
rect 21097 5729 21131 5763
rect 7297 5661 7331 5695
rect 10609 5661 10643 5695
rect 10885 5661 10919 5695
rect 11161 5661 11195 5695
rect 11253 5661 11287 5695
rect 11713 5661 11747 5695
rect 13277 5661 13311 5695
rect 14565 5661 14599 5695
rect 14749 5661 14783 5695
rect 14933 5661 14967 5695
rect 15301 5661 15335 5695
rect 15761 5661 15795 5695
rect 15945 5661 15979 5695
rect 16037 5661 16071 5695
rect 16175 5661 16209 5695
rect 16589 5661 16623 5695
rect 17141 5661 17175 5695
rect 17417 5661 17451 5695
rect 17545 5661 17579 5695
rect 18613 5661 18647 5695
rect 19303 5661 19337 5695
rect 10425 5593 10459 5627
rect 10517 5593 10551 5627
rect 10793 5593 10827 5627
rect 11069 5593 11103 5627
rect 12633 5593 12667 5627
rect 13001 5593 13035 5627
rect 13185 5593 13219 5627
rect 14841 5593 14875 5627
rect 17325 5593 17359 5627
rect 3249 5525 3283 5559
rect 11437 5525 11471 5559
rect 12081 5525 12115 5559
rect 15117 5525 15151 5559
rect 15393 5525 15427 5559
rect 15485 5525 15519 5559
rect 15669 5525 15703 5559
rect 16957 5525 16991 5559
rect 18705 5525 18739 5559
rect 5457 5321 5491 5355
rect 13461 5321 13495 5355
rect 16037 5321 16071 5355
rect 19901 5321 19935 5355
rect 3985 5253 4019 5287
rect 6745 5253 6779 5287
rect 9735 5253 9769 5287
rect 13553 5253 13587 5287
rect 14013 5253 14047 5287
rect 3709 5185 3743 5219
rect 7941 5185 7975 5219
rect 8309 5185 8343 5219
rect 11621 5185 11655 5219
rect 11713 5185 11747 5219
rect 11805 5185 11839 5219
rect 12909 5185 12943 5219
rect 13093 5185 13127 5219
rect 13369 5185 13403 5219
rect 13829 5185 13863 5219
rect 14105 5185 14139 5219
rect 14202 5207 14236 5241
rect 15669 5185 15703 5219
rect 15762 5185 15796 5219
rect 20085 5185 20119 5219
rect 11897 5117 11931 5151
rect 13185 5049 13219 5083
rect 13737 5049 13771 5083
rect 6653 4981 6687 5015
rect 12081 4981 12115 5015
rect 13001 4981 13035 5015
rect 13829 4981 13863 5015
rect 13001 4641 13035 4675
rect 12909 4573 12943 4607
rect 13277 4437 13311 4471
rect 15301 4233 15335 4267
rect 15393 4165 15427 4199
rect 13369 4097 13403 4131
rect 13553 4097 13587 4131
rect 13829 4097 13863 4131
rect 14105 4097 14139 4131
rect 14933 4097 14967 4131
rect 15577 4097 15611 4131
rect 15761 4097 15795 4131
rect 16037 4097 16071 4131
rect 16221 4097 16255 4131
rect 14197 4029 14231 4063
rect 14841 4029 14875 4063
rect 15853 4029 15887 4063
rect 13553 3961 13587 3995
rect 14381 3893 14415 3927
rect 14105 3689 14139 3723
rect 14841 3689 14875 3723
rect 24685 3689 24719 3723
rect 14105 3485 14139 3519
rect 14289 3485 14323 3519
rect 14749 3485 14783 3519
rect 14933 3485 14967 3519
rect 24869 3485 24903 3519
<< metal1 >>
rect 1104 26138 25208 26160
rect 1104 26086 4874 26138
rect 4926 26086 4938 26138
rect 4990 26086 5002 26138
rect 5054 26086 5066 26138
rect 5118 26086 5130 26138
rect 5182 26086 25208 26138
rect 1104 26064 25208 26086
rect 9214 25916 9220 25968
rect 9272 25916 9278 25968
rect 9858 25916 9864 25968
rect 9916 25916 9922 25968
rect 10502 25916 10508 25968
rect 10560 25916 10566 25968
rect 12342 25916 12348 25968
rect 12400 25956 12406 25968
rect 12437 25959 12495 25965
rect 12437 25956 12449 25959
rect 12400 25928 12449 25956
rect 12400 25916 12406 25928
rect 12437 25925 12449 25928
rect 12483 25925 12495 25959
rect 12437 25919 12495 25925
rect 13722 25916 13728 25968
rect 13780 25916 13786 25968
rect 14366 25916 14372 25968
rect 14424 25916 14430 25968
rect 15010 25916 15016 25968
rect 15068 25916 15074 25968
rect 17586 25916 17592 25968
rect 17644 25916 17650 25968
rect 18230 25916 18236 25968
rect 18288 25916 18294 25968
rect 3973 25891 4031 25897
rect 3973 25857 3985 25891
rect 4019 25888 4031 25891
rect 4706 25888 4712 25900
rect 4019 25860 4712 25888
rect 4019 25857 4031 25860
rect 3973 25851 4031 25857
rect 4706 25848 4712 25860
rect 4764 25848 4770 25900
rect 10870 25848 10876 25900
rect 10928 25888 10934 25900
rect 11241 25891 11299 25897
rect 11241 25888 11253 25891
rect 10928 25860 11253 25888
rect 10928 25848 10934 25860
rect 11241 25857 11253 25860
rect 11287 25857 11299 25891
rect 11241 25851 11299 25857
rect 11698 25848 11704 25900
rect 11756 25848 11762 25900
rect 12986 25848 12992 25900
rect 13044 25848 13050 25900
rect 15562 25848 15568 25900
rect 15620 25848 15626 25900
rect 16206 25848 16212 25900
rect 16264 25848 16270 25900
rect 4249 25823 4307 25829
rect 4249 25789 4261 25823
rect 4295 25820 4307 25823
rect 4614 25820 4620 25832
rect 4295 25792 4620 25820
rect 4295 25789 4307 25792
rect 4249 25783 4307 25789
rect 4614 25780 4620 25792
rect 4672 25780 4678 25832
rect 10045 25823 10103 25829
rect 10045 25789 10057 25823
rect 10091 25820 10103 25823
rect 10594 25820 10600 25832
rect 10091 25792 10600 25820
rect 10091 25789 10103 25792
rect 10045 25783 10103 25789
rect 10594 25780 10600 25792
rect 10652 25780 10658 25832
rect 15197 25823 15255 25829
rect 15197 25789 15209 25823
rect 15243 25820 15255 25823
rect 17494 25820 17500 25832
rect 15243 25792 17500 25820
rect 15243 25789 15255 25792
rect 15197 25783 15255 25789
rect 17494 25780 17500 25792
rect 17552 25780 17558 25832
rect 12621 25755 12679 25761
rect 12621 25721 12633 25755
rect 12667 25752 12679 25755
rect 12802 25752 12808 25764
rect 12667 25724 12808 25752
rect 12667 25721 12679 25724
rect 12621 25715 12679 25721
rect 12802 25712 12808 25724
rect 12860 25712 12866 25764
rect 13906 25712 13912 25764
rect 13964 25712 13970 25764
rect 14553 25755 14611 25761
rect 14553 25721 14565 25755
rect 14599 25752 14611 25755
rect 14642 25752 14648 25764
rect 14599 25724 14648 25752
rect 14599 25721 14611 25724
rect 14553 25715 14611 25721
rect 14642 25712 14648 25724
rect 14700 25712 14706 25764
rect 15749 25755 15807 25761
rect 15749 25721 15761 25755
rect 15795 25752 15807 25755
rect 17770 25752 17776 25764
rect 15795 25724 17776 25752
rect 15795 25721 15807 25724
rect 15749 25715 15807 25721
rect 17770 25712 17776 25724
rect 17828 25712 17834 25764
rect 18414 25712 18420 25764
rect 18472 25712 18478 25764
rect 2038 25644 2044 25696
rect 2096 25684 2102 25696
rect 3789 25687 3847 25693
rect 3789 25684 3801 25687
rect 2096 25656 3801 25684
rect 2096 25644 2102 25656
rect 3789 25653 3801 25656
rect 3835 25653 3847 25687
rect 3789 25647 3847 25653
rect 4157 25687 4215 25693
rect 4157 25653 4169 25687
rect 4203 25684 4215 25687
rect 4798 25684 4804 25696
rect 4203 25656 4804 25684
rect 4203 25653 4215 25656
rect 4157 25647 4215 25653
rect 4798 25644 4804 25656
rect 4856 25644 4862 25696
rect 9306 25644 9312 25696
rect 9364 25644 9370 25696
rect 10134 25644 10140 25696
rect 10192 25684 10198 25696
rect 10597 25687 10655 25693
rect 10597 25684 10609 25687
rect 10192 25656 10609 25684
rect 10192 25644 10198 25656
rect 10597 25653 10609 25656
rect 10643 25653 10655 25687
rect 10597 25647 10655 25653
rect 11054 25644 11060 25696
rect 11112 25644 11118 25696
rect 11882 25644 11888 25696
rect 11940 25644 11946 25696
rect 13173 25687 13231 25693
rect 13173 25653 13185 25687
rect 13219 25684 13231 25687
rect 13814 25684 13820 25696
rect 13219 25656 13820 25684
rect 13219 25653 13231 25656
rect 13173 25647 13231 25653
rect 13814 25644 13820 25656
rect 13872 25644 13878 25696
rect 16393 25687 16451 25693
rect 16393 25653 16405 25687
rect 16439 25684 16451 25687
rect 16942 25684 16948 25696
rect 16439 25656 16948 25684
rect 16439 25653 16451 25656
rect 16393 25647 16451 25653
rect 16942 25644 16948 25656
rect 17000 25644 17006 25696
rect 17402 25644 17408 25696
rect 17460 25684 17466 25696
rect 17681 25687 17739 25693
rect 17681 25684 17693 25687
rect 17460 25656 17693 25684
rect 17460 25644 17466 25656
rect 17681 25653 17693 25656
rect 17727 25653 17739 25687
rect 17681 25647 17739 25653
rect 1104 25594 25208 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 25208 25594
rect 1104 25520 25208 25542
rect 4433 25483 4491 25489
rect 4433 25449 4445 25483
rect 4479 25480 4491 25483
rect 4614 25480 4620 25492
rect 4479 25452 4620 25480
rect 4479 25449 4491 25452
rect 4433 25443 4491 25449
rect 4614 25440 4620 25452
rect 4672 25440 4678 25492
rect 4706 25440 4712 25492
rect 4764 25440 4770 25492
rect 2038 25304 2044 25356
rect 2096 25304 2102 25356
rect 3513 25347 3571 25353
rect 3513 25313 3525 25347
rect 3559 25344 3571 25347
rect 3694 25344 3700 25356
rect 3559 25316 3700 25344
rect 3559 25313 3571 25316
rect 3513 25307 3571 25313
rect 3694 25304 3700 25316
rect 3752 25344 3758 25356
rect 3789 25347 3847 25353
rect 3789 25344 3801 25347
rect 3752 25316 3801 25344
rect 3752 25304 3758 25316
rect 3789 25313 3801 25316
rect 3835 25313 3847 25347
rect 3789 25307 3847 25313
rect 4540 25316 5028 25344
rect 1394 25236 1400 25288
rect 1452 25276 1458 25288
rect 1765 25279 1823 25285
rect 1765 25276 1777 25279
rect 1452 25248 1777 25276
rect 1452 25236 1458 25248
rect 1765 25245 1777 25248
rect 1811 25245 1823 25279
rect 1765 25239 1823 25245
rect 4154 25236 4160 25288
rect 4212 25276 4218 25288
rect 4540 25285 4568 25316
rect 4525 25279 4583 25285
rect 4525 25276 4537 25279
rect 4212 25248 4537 25276
rect 4212 25236 4218 25248
rect 4525 25245 4537 25248
rect 4571 25245 4583 25279
rect 4525 25239 4583 25245
rect 4706 25236 4712 25288
rect 4764 25236 4770 25288
rect 4798 25236 4804 25288
rect 4856 25236 4862 25288
rect 5000 25285 5028 25316
rect 7668 25316 8340 25344
rect 4985 25279 5043 25285
rect 4985 25245 4997 25279
rect 5031 25245 5043 25279
rect 4985 25239 5043 25245
rect 5994 25236 6000 25288
rect 6052 25236 6058 25288
rect 3050 25168 3056 25220
rect 3108 25168 3114 25220
rect 4816 25208 4844 25236
rect 5350 25208 5356 25220
rect 4816 25180 5356 25208
rect 5350 25168 5356 25180
rect 5408 25168 5414 25220
rect 7374 25168 7380 25220
rect 7432 25208 7438 25220
rect 7668 25217 7696 25316
rect 8312 25285 8340 25316
rect 12066 25304 12072 25356
rect 12124 25344 12130 25356
rect 12124 25316 13308 25344
rect 12124 25304 12130 25316
rect 8205 25279 8263 25285
rect 8205 25245 8217 25279
rect 8251 25245 8263 25279
rect 8205 25239 8263 25245
rect 8297 25279 8355 25285
rect 8297 25245 8309 25279
rect 8343 25245 8355 25279
rect 8297 25239 8355 25245
rect 7653 25211 7711 25217
rect 7653 25208 7665 25211
rect 7432 25180 7665 25208
rect 7432 25168 7438 25180
rect 7653 25177 7665 25180
rect 7699 25177 7711 25211
rect 7653 25171 7711 25177
rect 7837 25211 7895 25217
rect 7837 25177 7849 25211
rect 7883 25208 7895 25211
rect 8220 25208 8248 25239
rect 8478 25236 8484 25288
rect 8536 25276 8542 25288
rect 8941 25279 8999 25285
rect 8941 25276 8953 25279
rect 8536 25248 8953 25276
rect 8536 25236 8542 25248
rect 8941 25245 8953 25248
rect 8987 25245 8999 25279
rect 8941 25239 8999 25245
rect 11054 25236 11060 25288
rect 11112 25236 11118 25288
rect 12986 25236 12992 25288
rect 13044 25236 13050 25288
rect 13280 25285 13308 25316
rect 13354 25304 13360 25356
rect 13412 25304 13418 25356
rect 19245 25347 19303 25353
rect 19245 25313 19257 25347
rect 19291 25344 19303 25347
rect 19518 25344 19524 25356
rect 19291 25316 19524 25344
rect 19291 25313 19303 25316
rect 19245 25307 19303 25313
rect 19518 25304 19524 25316
rect 19576 25304 19582 25356
rect 13265 25279 13323 25285
rect 13265 25245 13277 25279
rect 13311 25276 13323 25279
rect 15286 25276 15292 25288
rect 13311 25248 15292 25276
rect 13311 25245 13323 25248
rect 13265 25239 13323 25245
rect 15286 25236 15292 25248
rect 15344 25236 15350 25288
rect 15470 25236 15476 25288
rect 15528 25276 15534 25288
rect 15565 25279 15623 25285
rect 15565 25276 15577 25279
rect 15528 25248 15577 25276
rect 15528 25236 15534 25248
rect 15565 25245 15577 25248
rect 15611 25245 15623 25279
rect 15565 25239 15623 25245
rect 24854 25236 24860 25288
rect 24912 25236 24918 25288
rect 7883 25180 8708 25208
rect 7883 25177 7895 25180
rect 7837 25171 7895 25177
rect 4798 25100 4804 25152
rect 4856 25140 4862 25152
rect 4893 25143 4951 25149
rect 4893 25140 4905 25143
rect 4856 25112 4905 25140
rect 4856 25100 4862 25112
rect 4893 25109 4905 25112
rect 4939 25109 4951 25143
rect 4893 25103 4951 25109
rect 5258 25100 5264 25152
rect 5316 25140 5322 25152
rect 5445 25143 5503 25149
rect 5445 25140 5457 25143
rect 5316 25112 5457 25140
rect 5316 25100 5322 25112
rect 5445 25109 5457 25112
rect 5491 25109 5503 25143
rect 5445 25103 5503 25109
rect 7558 25100 7564 25152
rect 7616 25140 7622 25152
rect 7852 25140 7880 25171
rect 7616 25112 7880 25140
rect 8021 25143 8079 25149
rect 7616 25100 7622 25112
rect 8021 25109 8033 25143
rect 8067 25140 8079 25143
rect 8386 25140 8392 25152
rect 8067 25112 8392 25140
rect 8067 25109 8079 25112
rect 8021 25103 8079 25109
rect 8386 25100 8392 25112
rect 8444 25100 8450 25152
rect 8481 25143 8539 25149
rect 8481 25109 8493 25143
rect 8527 25140 8539 25143
rect 8570 25140 8576 25152
rect 8527 25112 8576 25140
rect 8527 25109 8539 25112
rect 8481 25103 8539 25109
rect 8570 25100 8576 25112
rect 8628 25100 8634 25152
rect 8680 25140 8708 25180
rect 9214 25168 9220 25220
rect 9272 25168 9278 25220
rect 9950 25168 9956 25220
rect 10008 25168 10014 25220
rect 11330 25168 11336 25220
rect 11388 25208 11394 25220
rect 11388 25180 11546 25208
rect 11388 25168 11394 25180
rect 12710 25168 12716 25220
rect 12768 25168 12774 25220
rect 15838 25168 15844 25220
rect 15896 25168 15902 25220
rect 16850 25168 16856 25220
rect 16908 25168 16914 25220
rect 19426 25168 19432 25220
rect 19484 25208 19490 25220
rect 19521 25211 19579 25217
rect 19521 25208 19533 25211
rect 19484 25180 19533 25208
rect 19484 25168 19490 25180
rect 19521 25177 19533 25180
rect 19567 25177 19579 25211
rect 21082 25208 21088 25220
rect 20746 25180 21088 25208
rect 19521 25171 19579 25177
rect 21082 25168 21088 25180
rect 21140 25168 21146 25220
rect 10502 25140 10508 25152
rect 8680 25112 10508 25140
rect 10502 25100 10508 25112
rect 10560 25140 10566 25152
rect 10689 25143 10747 25149
rect 10689 25140 10701 25143
rect 10560 25112 10701 25140
rect 10560 25100 10566 25112
rect 10689 25109 10701 25112
rect 10735 25109 10747 25143
rect 10689 25103 10747 25109
rect 10962 25100 10968 25152
rect 11020 25100 11026 25152
rect 11238 25100 11244 25152
rect 11296 25100 11302 25152
rect 13538 25100 13544 25152
rect 13596 25140 13602 25152
rect 13633 25143 13691 25149
rect 13633 25140 13645 25143
rect 13596 25112 13645 25140
rect 13596 25100 13602 25112
rect 13633 25109 13645 25112
rect 13679 25109 13691 25143
rect 13633 25103 13691 25109
rect 17313 25143 17371 25149
rect 17313 25109 17325 25143
rect 17359 25140 17371 25143
rect 17586 25140 17592 25152
rect 17359 25112 17592 25140
rect 17359 25109 17371 25112
rect 17313 25103 17371 25109
rect 17586 25100 17592 25112
rect 17644 25100 17650 25152
rect 20990 25100 20996 25152
rect 21048 25100 21054 25152
rect 1104 25050 25208 25072
rect 1104 24998 4874 25050
rect 4926 24998 4938 25050
rect 4990 24998 5002 25050
rect 5054 24998 5066 25050
rect 5118 24998 5130 25050
rect 5182 24998 25208 25050
rect 1104 24976 25208 24998
rect 3050 24896 3056 24948
rect 3108 24936 3114 24948
rect 5905 24939 5963 24945
rect 3108 24908 5764 24936
rect 3108 24896 3114 24908
rect 3068 24868 3096 24896
rect 5736 24868 5764 24908
rect 5905 24905 5917 24939
rect 5951 24936 5963 24939
rect 5994 24936 6000 24948
rect 5951 24908 6000 24936
rect 5951 24905 5963 24908
rect 5905 24899 5963 24905
rect 5994 24896 6000 24908
rect 6052 24896 6058 24948
rect 9125 24939 9183 24945
rect 6104 24908 7880 24936
rect 6104 24868 6132 24908
rect 7852 24868 7880 24908
rect 9125 24905 9137 24939
rect 9171 24936 9183 24939
rect 9214 24936 9220 24948
rect 9171 24908 9220 24936
rect 9171 24905 9183 24908
rect 9125 24899 9183 24905
rect 9214 24896 9220 24908
rect 9272 24896 9278 24948
rect 14734 24896 14740 24948
rect 14792 24936 14798 24948
rect 14829 24939 14887 24945
rect 14829 24936 14841 24939
rect 14792 24908 14841 24936
rect 14792 24896 14798 24908
rect 14829 24905 14841 24908
rect 14875 24936 14887 24939
rect 15657 24939 15715 24945
rect 14875 24908 15240 24936
rect 14875 24905 14887 24908
rect 14829 24899 14887 24905
rect 8754 24868 8760 24880
rect 2990 24840 3096 24868
rect 5658 24840 6132 24868
rect 7774 24840 8760 24868
rect 8754 24828 8760 24840
rect 8812 24828 8818 24880
rect 8941 24871 8999 24877
rect 8941 24837 8953 24871
rect 8987 24837 8999 24871
rect 9232 24868 9260 24896
rect 9232 24840 9628 24868
rect 8941 24831 8999 24837
rect 8478 24760 8484 24812
rect 8536 24760 8542 24812
rect 8662 24760 8668 24812
rect 8720 24800 8726 24812
rect 8956 24800 8984 24831
rect 8720 24772 8984 24800
rect 8720 24760 8726 24772
rect 9214 24760 9220 24812
rect 9272 24760 9278 24812
rect 9398 24760 9404 24812
rect 9456 24760 9462 24812
rect 1394 24692 1400 24744
rect 1452 24732 1458 24744
rect 1489 24735 1547 24741
rect 1489 24732 1501 24735
rect 1452 24704 1501 24732
rect 1452 24692 1458 24704
rect 1489 24701 1501 24704
rect 1535 24701 1547 24735
rect 1489 24695 1547 24701
rect 1504 24596 1532 24695
rect 1762 24692 1768 24744
rect 1820 24692 1826 24744
rect 3237 24735 3295 24741
rect 3237 24701 3249 24735
rect 3283 24732 3295 24735
rect 3878 24732 3884 24744
rect 3283 24704 3884 24732
rect 3283 24701 3295 24704
rect 3237 24695 3295 24701
rect 3878 24692 3884 24704
rect 3936 24692 3942 24744
rect 4157 24735 4215 24741
rect 4157 24701 4169 24735
rect 4203 24701 4215 24735
rect 4157 24695 4215 24701
rect 4433 24735 4491 24741
rect 4433 24701 4445 24735
rect 4479 24732 4491 24735
rect 4522 24732 4528 24744
rect 4479 24704 4528 24732
rect 4479 24701 4491 24704
rect 4433 24695 4491 24701
rect 4172 24664 4200 24695
rect 4522 24692 4528 24704
rect 4580 24692 4586 24744
rect 8202 24692 8208 24744
rect 8260 24692 8266 24744
rect 9600 24741 9628 24840
rect 9677 24803 9735 24809
rect 9677 24769 9689 24803
rect 9723 24800 9735 24803
rect 10778 24800 10784 24812
rect 9723 24772 10784 24800
rect 9723 24769 9735 24772
rect 9677 24763 9735 24769
rect 10778 24760 10784 24772
rect 10836 24760 10842 24812
rect 12526 24760 12532 24812
rect 12584 24800 12590 24812
rect 12621 24803 12679 24809
rect 12621 24800 12633 24803
rect 12584 24772 12633 24800
rect 12584 24760 12590 24772
rect 12621 24769 12633 24772
rect 12667 24769 12679 24803
rect 12621 24763 12679 24769
rect 14458 24760 14464 24812
rect 14516 24760 14522 24812
rect 15212 24809 15240 24908
rect 15657 24905 15669 24939
rect 15703 24936 15715 24939
rect 15838 24936 15844 24948
rect 15703 24908 15844 24936
rect 15703 24905 15715 24908
rect 15657 24899 15715 24905
rect 15838 24896 15844 24908
rect 15896 24896 15902 24948
rect 18233 24939 18291 24945
rect 18233 24905 18245 24939
rect 18279 24936 18291 24939
rect 19886 24936 19892 24948
rect 18279 24908 19892 24936
rect 18279 24905 18291 24908
rect 18233 24899 18291 24905
rect 19886 24896 19892 24908
rect 19944 24896 19950 24948
rect 17037 24871 17095 24877
rect 17037 24837 17049 24871
rect 17083 24868 17095 24871
rect 17586 24868 17592 24880
rect 17083 24840 17592 24868
rect 17083 24837 17095 24840
rect 17037 24831 17095 24837
rect 17586 24828 17592 24840
rect 17644 24828 17650 24880
rect 17862 24868 17868 24880
rect 17696 24840 17868 24868
rect 15105 24803 15163 24809
rect 15105 24800 15117 24803
rect 14568 24772 15117 24800
rect 9585 24735 9643 24741
rect 9585 24701 9597 24735
rect 9631 24701 9643 24735
rect 9585 24695 9643 24701
rect 12710 24692 12716 24744
rect 12768 24692 12774 24744
rect 12986 24692 12992 24744
rect 13044 24732 13050 24744
rect 13081 24735 13139 24741
rect 13081 24732 13093 24735
rect 13044 24704 13093 24732
rect 13044 24692 13050 24704
rect 13081 24701 13093 24704
rect 13127 24701 13139 24735
rect 13081 24695 13139 24701
rect 8573 24667 8631 24673
rect 8573 24664 8585 24667
rect 3160 24636 4200 24664
rect 8404 24636 8585 24664
rect 3160 24596 3188 24636
rect 8404 24608 8432 24636
rect 8573 24633 8585 24636
rect 8619 24633 8631 24667
rect 8573 24627 8631 24633
rect 8754 24624 8760 24676
rect 8812 24664 8818 24676
rect 9950 24664 9956 24676
rect 8812 24636 9956 24664
rect 8812 24624 8818 24636
rect 9950 24624 9956 24636
rect 10008 24624 10014 24676
rect 1504 24568 3188 24596
rect 3326 24556 3332 24608
rect 3384 24556 3390 24608
rect 6733 24599 6791 24605
rect 6733 24565 6745 24599
rect 6779 24596 6791 24599
rect 7190 24596 7196 24608
rect 6779 24568 7196 24596
rect 6779 24565 6791 24568
rect 6733 24559 6791 24565
rect 7190 24556 7196 24568
rect 7248 24556 7254 24608
rect 8386 24556 8392 24608
rect 8444 24556 8450 24608
rect 8478 24556 8484 24608
rect 8536 24596 8542 24608
rect 8941 24599 8999 24605
rect 8941 24596 8953 24599
rect 8536 24568 8953 24596
rect 8536 24556 8542 24568
rect 8941 24565 8953 24568
rect 8987 24565 8999 24599
rect 8941 24559 8999 24565
rect 9030 24556 9036 24608
rect 9088 24596 9094 24608
rect 9217 24599 9275 24605
rect 9217 24596 9229 24599
rect 9088 24568 9229 24596
rect 9088 24556 9094 24568
rect 9217 24565 9229 24568
rect 9263 24565 9275 24599
rect 9217 24559 9275 24565
rect 10045 24599 10103 24605
rect 10045 24565 10057 24599
rect 10091 24596 10103 24599
rect 10226 24596 10232 24608
rect 10091 24568 10232 24596
rect 10091 24565 10103 24568
rect 10045 24559 10103 24565
rect 10226 24556 10232 24568
rect 10284 24556 10290 24608
rect 12894 24556 12900 24608
rect 12952 24556 12958 24608
rect 13096 24596 13124 24695
rect 13354 24692 13360 24744
rect 13412 24692 13418 24744
rect 13722 24692 13728 24744
rect 13780 24732 13786 24744
rect 14568 24732 14596 24772
rect 15105 24769 15117 24772
rect 15151 24769 15163 24803
rect 15105 24763 15163 24769
rect 15197 24803 15255 24809
rect 15197 24769 15209 24803
rect 15243 24769 15255 24803
rect 15197 24763 15255 24769
rect 15749 24803 15807 24809
rect 15749 24769 15761 24803
rect 15795 24769 15807 24803
rect 15749 24763 15807 24769
rect 13780 24704 14596 24732
rect 13780 24692 13786 24704
rect 14918 24692 14924 24744
rect 14976 24692 14982 24744
rect 15470 24664 15476 24676
rect 14384 24636 15476 24664
rect 14384 24596 14412 24636
rect 15470 24624 15476 24636
rect 15528 24624 15534 24676
rect 13096 24568 14412 24596
rect 15010 24556 15016 24608
rect 15068 24556 15074 24608
rect 15764 24596 15792 24763
rect 16022 24760 16028 24812
rect 16080 24760 16086 24812
rect 16853 24803 16911 24809
rect 16853 24769 16865 24803
rect 16899 24769 16911 24803
rect 16853 24763 16911 24769
rect 16114 24692 16120 24744
rect 16172 24692 16178 24744
rect 16868 24732 16896 24763
rect 17126 24760 17132 24812
rect 17184 24760 17190 24812
rect 17218 24760 17224 24812
rect 17276 24760 17282 24812
rect 17405 24803 17463 24809
rect 17405 24769 17417 24803
rect 17451 24769 17463 24803
rect 17696 24800 17724 24840
rect 17862 24828 17868 24840
rect 17920 24828 17926 24880
rect 21082 24868 21088 24880
rect 17972 24840 18368 24868
rect 21022 24840 21088 24868
rect 17405 24763 17463 24769
rect 17512 24772 17724 24800
rect 17310 24732 17316 24744
rect 16868 24704 17316 24732
rect 17310 24692 17316 24704
rect 17368 24692 17374 24744
rect 16393 24667 16451 24673
rect 16393 24633 16405 24667
rect 16439 24664 16451 24667
rect 17126 24664 17132 24676
rect 16439 24636 17132 24664
rect 16439 24633 16451 24636
rect 16393 24627 16451 24633
rect 17126 24624 17132 24636
rect 17184 24624 17190 24676
rect 17420 24664 17448 24763
rect 17512 24744 17540 24772
rect 17770 24760 17776 24812
rect 17828 24760 17834 24812
rect 17494 24692 17500 24744
rect 17552 24692 17558 24744
rect 17589 24735 17647 24741
rect 17589 24701 17601 24735
rect 17635 24732 17647 24735
rect 17678 24732 17684 24744
rect 17635 24704 17684 24732
rect 17635 24701 17647 24704
rect 17589 24695 17647 24701
rect 17678 24692 17684 24704
rect 17736 24732 17742 24744
rect 17972 24732 18000 24840
rect 18049 24803 18107 24809
rect 18049 24769 18061 24803
rect 18095 24769 18107 24803
rect 18049 24763 18107 24769
rect 17736 24704 18000 24732
rect 17736 24692 17742 24704
rect 18064 24664 18092 24763
rect 18138 24760 18144 24812
rect 18196 24800 18202 24812
rect 18233 24803 18291 24809
rect 18233 24800 18245 24803
rect 18196 24772 18245 24800
rect 18196 24760 18202 24772
rect 18233 24769 18245 24772
rect 18279 24769 18291 24803
rect 18340 24800 18368 24840
rect 21082 24828 21088 24840
rect 21140 24868 21146 24880
rect 21542 24868 21548 24880
rect 21140 24840 21548 24868
rect 21140 24828 21146 24840
rect 21542 24828 21548 24840
rect 21600 24828 21606 24880
rect 19153 24803 19211 24809
rect 19153 24800 19165 24803
rect 18340 24772 19165 24800
rect 18233 24763 18291 24769
rect 19153 24769 19165 24772
rect 19199 24769 19211 24803
rect 19153 24763 19211 24769
rect 19245 24803 19303 24809
rect 19245 24769 19257 24803
rect 19291 24800 19303 24803
rect 19426 24800 19432 24812
rect 19291 24772 19432 24800
rect 19291 24769 19303 24772
rect 19245 24763 19303 24769
rect 19168 24732 19196 24763
rect 19426 24760 19432 24772
rect 19484 24760 19490 24812
rect 21358 24760 21364 24812
rect 21416 24800 21422 24812
rect 22189 24803 22247 24809
rect 22189 24800 22201 24803
rect 21416 24772 22201 24800
rect 21416 24760 21422 24772
rect 22189 24769 22201 24772
rect 22235 24769 22247 24803
rect 22189 24763 22247 24769
rect 22370 24760 22376 24812
rect 22428 24800 22434 24812
rect 22465 24803 22523 24809
rect 22465 24800 22477 24803
rect 22428 24772 22477 24800
rect 22428 24760 22434 24772
rect 22465 24769 22477 24772
rect 22511 24769 22523 24803
rect 22465 24763 22523 24769
rect 22646 24760 22652 24812
rect 22704 24760 22710 24812
rect 19334 24732 19340 24744
rect 19168 24704 19340 24732
rect 19334 24692 19340 24704
rect 19392 24692 19398 24744
rect 19518 24692 19524 24744
rect 19576 24692 19582 24744
rect 19794 24692 19800 24744
rect 19852 24692 19858 24744
rect 22281 24735 22339 24741
rect 22281 24701 22293 24735
rect 22327 24732 22339 24735
rect 22327 24704 22692 24732
rect 22327 24701 22339 24704
rect 22281 24695 22339 24701
rect 17420 24636 18092 24664
rect 16669 24599 16727 24605
rect 16669 24596 16681 24599
rect 15764 24568 16681 24596
rect 16669 24565 16681 24568
rect 16715 24596 16727 24599
rect 17420 24596 17448 24636
rect 16715 24568 17448 24596
rect 17957 24599 18015 24605
rect 16715 24565 16727 24568
rect 16669 24559 16727 24565
rect 17957 24565 17969 24599
rect 18003 24596 18015 24599
rect 19426 24596 19432 24608
rect 18003 24568 19432 24596
rect 18003 24565 18015 24568
rect 17957 24559 18015 24565
rect 19426 24556 19432 24568
rect 19484 24556 19490 24608
rect 19536 24596 19564 24692
rect 20806 24624 20812 24676
rect 20864 24664 20870 24676
rect 21821 24667 21879 24673
rect 21821 24664 21833 24667
rect 20864 24636 21833 24664
rect 20864 24624 20870 24636
rect 21821 24633 21833 24636
rect 21867 24633 21879 24667
rect 21821 24627 21879 24633
rect 20530 24596 20536 24608
rect 19536 24568 20536 24596
rect 20530 24556 20536 24568
rect 20588 24556 20594 24608
rect 21174 24556 21180 24608
rect 21232 24596 21238 24608
rect 22664 24605 22692 24704
rect 21269 24599 21327 24605
rect 21269 24596 21281 24599
rect 21232 24568 21281 24596
rect 21232 24556 21238 24568
rect 21269 24565 21281 24568
rect 21315 24565 21327 24599
rect 21269 24559 21327 24565
rect 22649 24599 22707 24605
rect 22649 24565 22661 24599
rect 22695 24596 22707 24599
rect 23014 24596 23020 24608
rect 22695 24568 23020 24596
rect 22695 24565 22707 24568
rect 22649 24559 22707 24565
rect 23014 24556 23020 24568
rect 23072 24556 23078 24608
rect 1104 24506 25208 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 25208 24506
rect 1104 24432 25208 24454
rect 3878 24352 3884 24404
rect 3936 24392 3942 24404
rect 4246 24392 4252 24404
rect 3936 24364 4252 24392
rect 3936 24352 3942 24364
rect 4246 24352 4252 24364
rect 4304 24352 4310 24404
rect 4338 24352 4344 24404
rect 4396 24392 4402 24404
rect 4798 24392 4804 24404
rect 4396 24364 4804 24392
rect 4396 24352 4402 24364
rect 4798 24352 4804 24364
rect 4856 24352 4862 24404
rect 7190 24352 7196 24404
rect 7248 24392 7254 24404
rect 7377 24395 7435 24401
rect 7377 24392 7389 24395
rect 7248 24364 7389 24392
rect 7248 24352 7254 24364
rect 7377 24361 7389 24364
rect 7423 24361 7435 24395
rect 7377 24355 7435 24361
rect 8205 24395 8263 24401
rect 8205 24361 8217 24395
rect 8251 24392 8263 24395
rect 8294 24392 8300 24404
rect 8251 24364 8300 24392
rect 8251 24361 8263 24364
rect 8205 24355 8263 24361
rect 8294 24352 8300 24364
rect 8352 24352 8358 24404
rect 8386 24352 8392 24404
rect 8444 24392 8450 24404
rect 8570 24392 8576 24404
rect 8444 24364 8576 24392
rect 8444 24352 8450 24364
rect 8570 24352 8576 24364
rect 8628 24352 8634 24404
rect 10502 24352 10508 24404
rect 10560 24392 10566 24404
rect 11146 24392 11152 24404
rect 10560 24364 11152 24392
rect 10560 24352 10566 24364
rect 11146 24352 11152 24364
rect 11204 24352 11210 24404
rect 12621 24395 12679 24401
rect 12621 24361 12633 24395
rect 12667 24392 12679 24395
rect 12710 24392 12716 24404
rect 12667 24364 12716 24392
rect 12667 24361 12679 24364
rect 12621 24355 12679 24361
rect 12710 24352 12716 24364
rect 12768 24352 12774 24404
rect 12989 24395 13047 24401
rect 12989 24361 13001 24395
rect 13035 24392 13047 24395
rect 13354 24392 13360 24404
rect 13035 24364 13360 24392
rect 13035 24361 13047 24364
rect 12989 24355 13047 24361
rect 13354 24352 13360 24364
rect 13412 24352 13418 24404
rect 15644 24395 15702 24401
rect 15644 24361 15656 24395
rect 15690 24392 15702 24395
rect 16114 24392 16120 24404
rect 15690 24364 16120 24392
rect 15690 24361 15702 24364
rect 15644 24355 15702 24361
rect 16114 24352 16120 24364
rect 16172 24352 16178 24404
rect 17218 24352 17224 24404
rect 17276 24352 17282 24404
rect 17310 24352 17316 24404
rect 17368 24392 17374 24404
rect 17773 24395 17831 24401
rect 17773 24392 17785 24395
rect 17368 24364 17785 24392
rect 17368 24352 17374 24364
rect 17773 24361 17785 24364
rect 17819 24361 17831 24395
rect 18693 24395 18751 24401
rect 18693 24392 18705 24395
rect 17773 24355 17831 24361
rect 18432 24364 18705 24392
rect 1762 24284 1768 24336
rect 1820 24324 1826 24336
rect 2041 24327 2099 24333
rect 2041 24324 2053 24327
rect 1820 24296 2053 24324
rect 1820 24284 1826 24296
rect 2041 24293 2053 24296
rect 2087 24293 2099 24327
rect 4614 24324 4620 24336
rect 2041 24287 2099 24293
rect 2516 24296 4620 24324
rect 2516 24265 2544 24296
rect 4614 24284 4620 24296
rect 4672 24284 4678 24336
rect 8110 24324 8116 24336
rect 6932 24296 8116 24324
rect 2501 24259 2559 24265
rect 2501 24225 2513 24259
rect 2547 24225 2559 24259
rect 3513 24259 3571 24265
rect 3513 24256 3525 24259
rect 2501 24219 2559 24225
rect 3068 24228 3525 24256
rect 3068 24197 3096 24228
rect 3513 24225 3525 24228
rect 3559 24225 3571 24259
rect 3513 24219 3571 24225
rect 3694 24216 3700 24268
rect 3752 24256 3758 24268
rect 6932 24265 6960 24296
rect 8110 24284 8116 24296
rect 8168 24284 8174 24336
rect 8481 24327 8539 24333
rect 8481 24293 8493 24327
rect 8527 24324 8539 24327
rect 9214 24324 9220 24336
rect 8527 24296 9220 24324
rect 8527 24293 8539 24296
rect 8481 24287 8539 24293
rect 9214 24284 9220 24296
rect 9272 24284 9278 24336
rect 10778 24284 10784 24336
rect 10836 24284 10842 24336
rect 13081 24327 13139 24333
rect 13081 24324 13093 24327
rect 11072 24296 13093 24324
rect 6917 24259 6975 24265
rect 3752 24228 4384 24256
rect 3752 24216 3758 24228
rect 3053 24191 3111 24197
rect 3053 24157 3065 24191
rect 3099 24157 3111 24191
rect 3053 24151 3111 24157
rect 3234 24148 3240 24200
rect 3292 24148 3298 24200
rect 3329 24191 3387 24197
rect 3329 24157 3341 24191
rect 3375 24157 3387 24191
rect 3329 24151 3387 24157
rect 2038 24080 2044 24132
rect 2096 24080 2102 24132
rect 2593 24123 2651 24129
rect 2593 24089 2605 24123
rect 2639 24120 2651 24123
rect 3344 24120 3372 24151
rect 3418 24148 3424 24200
rect 3476 24148 3482 24200
rect 3602 24148 3608 24200
rect 3660 24148 3666 24200
rect 3878 24148 3884 24200
rect 3936 24148 3942 24200
rect 3973 24191 4031 24197
rect 3973 24157 3985 24191
rect 4019 24188 4031 24191
rect 4154 24188 4160 24200
rect 4019 24160 4160 24188
rect 4019 24157 4031 24160
rect 3973 24151 4031 24157
rect 4154 24148 4160 24160
rect 4212 24148 4218 24200
rect 4356 24197 4384 24228
rect 6917 24225 6929 24259
rect 6963 24225 6975 24259
rect 7929 24259 7987 24265
rect 6917 24219 6975 24225
rect 7116 24228 7788 24256
rect 4341 24191 4399 24197
rect 4341 24157 4353 24191
rect 4387 24157 4399 24191
rect 4709 24191 4767 24197
rect 4709 24188 4721 24191
rect 4341 24151 4399 24157
rect 4448 24160 4721 24188
rect 3896 24120 3924 24148
rect 2639 24092 2912 24120
rect 3344 24092 3924 24120
rect 2639 24089 2651 24092
rect 2593 24083 2651 24089
rect 2884 24064 2912 24092
rect 2774 24012 2780 24064
rect 2832 24012 2838 24064
rect 2866 24012 2872 24064
rect 2924 24012 2930 24064
rect 3602 24012 3608 24064
rect 3660 24052 3666 24064
rect 4062 24052 4068 24064
rect 3660 24024 4068 24052
rect 3660 24012 3666 24024
rect 4062 24012 4068 24024
rect 4120 24052 4126 24064
rect 4448 24052 4476 24160
rect 4709 24157 4721 24160
rect 4755 24157 4767 24191
rect 4709 24151 4767 24157
rect 4798 24148 4804 24200
rect 4856 24148 4862 24200
rect 4985 24191 5043 24197
rect 4985 24157 4997 24191
rect 5031 24188 5043 24191
rect 5258 24188 5264 24200
rect 5031 24160 5264 24188
rect 5031 24157 5043 24160
rect 4985 24151 5043 24157
rect 5258 24148 5264 24160
rect 5316 24148 5322 24200
rect 5077 24123 5135 24129
rect 5077 24120 5089 24123
rect 4724 24092 5089 24120
rect 4724 24064 4752 24092
rect 5077 24089 5089 24092
rect 5123 24089 5135 24123
rect 5077 24083 5135 24089
rect 6178 24080 6184 24132
rect 6236 24080 6242 24132
rect 6641 24123 6699 24129
rect 6641 24089 6653 24123
rect 6687 24120 6699 24123
rect 7116 24120 7144 24228
rect 7466 24120 7472 24132
rect 6687 24092 7144 24120
rect 7208 24092 7472 24120
rect 6687 24089 6699 24092
rect 6641 24083 6699 24089
rect 4120 24024 4476 24052
rect 4120 24012 4126 24024
rect 4522 24012 4528 24064
rect 4580 24012 4586 24064
rect 4706 24012 4712 24064
rect 4764 24012 4770 24064
rect 5169 24055 5227 24061
rect 5169 24021 5181 24055
rect 5215 24052 5227 24055
rect 5258 24052 5264 24064
rect 5215 24024 5264 24052
rect 5215 24021 5227 24024
rect 5169 24015 5227 24021
rect 5258 24012 5264 24024
rect 5316 24012 5322 24064
rect 6914 24012 6920 24064
rect 6972 24052 6978 24064
rect 7208 24061 7236 24092
rect 7466 24080 7472 24092
rect 7524 24080 7530 24132
rect 7558 24080 7564 24132
rect 7616 24080 7622 24132
rect 7374 24061 7380 24064
rect 7193 24055 7251 24061
rect 7193 24052 7205 24055
rect 6972 24024 7205 24052
rect 6972 24012 6978 24024
rect 7193 24021 7205 24024
rect 7239 24021 7251 24055
rect 7193 24015 7251 24021
rect 7361 24055 7380 24061
rect 7361 24021 7373 24055
rect 7361 24015 7380 24021
rect 7374 24012 7380 24015
rect 7432 24012 7438 24064
rect 7760 24052 7788 24228
rect 7929 24225 7941 24259
rect 7975 24256 7987 24259
rect 8202 24256 8208 24268
rect 7975 24228 8208 24256
rect 7975 24225 7987 24228
rect 7929 24219 7987 24225
rect 8202 24216 8208 24228
rect 8260 24216 8266 24268
rect 8573 24259 8631 24265
rect 8573 24225 8585 24259
rect 8619 24256 8631 24259
rect 8662 24256 8668 24268
rect 8619 24228 8668 24256
rect 8619 24225 8631 24228
rect 8573 24219 8631 24225
rect 8662 24216 8668 24228
rect 8720 24216 8726 24268
rect 11072 24256 11100 24296
rect 13081 24293 13093 24296
rect 13127 24293 13139 24327
rect 13081 24287 13139 24293
rect 17034 24284 17040 24336
rect 17092 24324 17098 24336
rect 17681 24327 17739 24333
rect 17681 24324 17693 24327
rect 17092 24296 17693 24324
rect 17092 24284 17098 24296
rect 17681 24293 17693 24296
rect 17727 24324 17739 24327
rect 18432 24324 18460 24364
rect 18693 24361 18705 24364
rect 18739 24361 18751 24395
rect 18693 24355 18751 24361
rect 18874 24352 18880 24404
rect 18932 24352 18938 24404
rect 19337 24395 19395 24401
rect 19337 24361 19349 24395
rect 19383 24392 19395 24395
rect 19794 24392 19800 24404
rect 19383 24364 19800 24392
rect 19383 24361 19395 24364
rect 19337 24355 19395 24361
rect 17727 24296 18460 24324
rect 17727 24293 17739 24296
rect 17681 24287 17739 24293
rect 12802 24256 12808 24268
rect 10244 24228 11100 24256
rect 12360 24228 12808 24256
rect 7834 24148 7840 24200
rect 7892 24148 7898 24200
rect 8297 24191 8355 24197
rect 8297 24157 8309 24191
rect 8343 24188 8355 24191
rect 8386 24188 8392 24200
rect 8343 24160 8392 24188
rect 8343 24157 8355 24160
rect 8297 24151 8355 24157
rect 8386 24148 8392 24160
rect 8444 24148 8450 24200
rect 10244 24197 10272 24228
rect 10229 24191 10287 24197
rect 10229 24157 10241 24191
rect 10275 24157 10287 24191
rect 10229 24151 10287 24157
rect 10410 24148 10416 24200
rect 10468 24148 10474 24200
rect 10502 24148 10508 24200
rect 10560 24148 10566 24200
rect 10778 24148 10784 24200
rect 10836 24188 10842 24200
rect 11057 24191 11115 24197
rect 11057 24188 11069 24191
rect 10836 24160 11069 24188
rect 10836 24148 10842 24160
rect 11057 24157 11069 24160
rect 11103 24157 11115 24191
rect 11057 24151 11115 24157
rect 11072 24120 11100 24151
rect 11146 24148 11152 24200
rect 11204 24188 11210 24200
rect 11204 24160 11249 24188
rect 11204 24148 11210 24160
rect 12360 24120 12388 24228
rect 12802 24216 12808 24228
rect 12860 24216 12866 24268
rect 12894 24216 12900 24268
rect 12952 24256 12958 24268
rect 12952 24228 13676 24256
rect 12952 24216 12958 24228
rect 12437 24191 12495 24197
rect 12437 24157 12449 24191
rect 12483 24157 12495 24191
rect 12437 24151 12495 24157
rect 11072 24092 12388 24120
rect 12452 24120 12480 24151
rect 12618 24148 12624 24200
rect 12676 24148 12682 24200
rect 12713 24191 12771 24197
rect 12713 24157 12725 24191
rect 12759 24188 12771 24191
rect 12759 24160 12940 24188
rect 12759 24157 12771 24160
rect 12713 24151 12771 24157
rect 12912 24120 12940 24160
rect 13262 24148 13268 24200
rect 13320 24148 13326 24200
rect 13354 24148 13360 24200
rect 13412 24148 13418 24200
rect 13538 24148 13544 24200
rect 13596 24148 13602 24200
rect 13648 24197 13676 24228
rect 14458 24216 14464 24268
rect 14516 24256 14522 24268
rect 16850 24256 16856 24268
rect 14516 24228 16856 24256
rect 14516 24216 14522 24228
rect 13633 24191 13691 24197
rect 13633 24157 13645 24191
rect 13679 24157 13691 24191
rect 13633 24151 13691 24157
rect 15378 24148 15384 24200
rect 15436 24148 15442 24200
rect 16776 24174 16804 24228
rect 16850 24216 16856 24228
rect 16908 24216 16914 24268
rect 17865 24259 17923 24265
rect 17865 24225 17877 24259
rect 17911 24225 17923 24259
rect 17865 24219 17923 24225
rect 17126 24148 17132 24200
rect 17184 24188 17190 24200
rect 17221 24191 17279 24197
rect 17221 24188 17233 24191
rect 17184 24160 17233 24188
rect 17184 24148 17190 24160
rect 17221 24157 17233 24160
rect 17267 24157 17279 24191
rect 17221 24151 17279 24157
rect 17497 24191 17555 24197
rect 17497 24157 17509 24191
rect 17543 24157 17555 24191
rect 17497 24151 17555 24157
rect 12452 24092 12940 24120
rect 10321 24055 10379 24061
rect 10321 24052 10333 24055
rect 7760 24024 10333 24052
rect 10321 24021 10333 24024
rect 10367 24021 10379 24055
rect 10321 24015 10379 24021
rect 10965 24055 11023 24061
rect 10965 24021 10977 24055
rect 11011 24052 11023 24055
rect 11054 24052 11060 24064
rect 11011 24024 11060 24052
rect 11011 24021 11023 24024
rect 10965 24015 11023 24021
rect 11054 24012 11060 24024
rect 11112 24012 11118 24064
rect 11425 24055 11483 24061
rect 11425 24021 11437 24055
rect 11471 24052 11483 24055
rect 11790 24052 11796 24064
rect 11471 24024 11796 24052
rect 11471 24021 11483 24024
rect 11425 24015 11483 24021
rect 11790 24012 11796 24024
rect 11848 24012 11854 24064
rect 12710 24012 12716 24064
rect 12768 24052 12774 24064
rect 12805 24055 12863 24061
rect 12805 24052 12817 24055
rect 12768 24024 12817 24052
rect 12768 24012 12774 24024
rect 12805 24021 12817 24024
rect 12851 24021 12863 24055
rect 12912 24052 12940 24092
rect 12989 24123 13047 24129
rect 12989 24089 13001 24123
rect 13035 24120 13047 24123
rect 15010 24120 15016 24132
rect 13035 24092 15016 24120
rect 13035 24089 13047 24092
rect 12989 24083 13047 24089
rect 15010 24080 15016 24092
rect 15068 24080 15074 24132
rect 17512 24120 17540 24151
rect 17586 24148 17592 24200
rect 17644 24148 17650 24200
rect 17678 24120 17684 24132
rect 17512 24092 17684 24120
rect 17678 24080 17684 24092
rect 17736 24080 17742 24132
rect 13722 24052 13728 24064
rect 12912 24024 13728 24052
rect 12805 24015 12863 24021
rect 13722 24012 13728 24024
rect 13780 24012 13786 24064
rect 16574 24012 16580 24064
rect 16632 24052 16638 24064
rect 17129 24055 17187 24061
rect 17129 24052 17141 24055
rect 16632 24024 17141 24052
rect 16632 24012 16638 24024
rect 17129 24021 17141 24024
rect 17175 24021 17187 24055
rect 17129 24015 17187 24021
rect 17405 24055 17463 24061
rect 17405 24021 17417 24055
rect 17451 24052 17463 24055
rect 17770 24052 17776 24064
rect 17451 24024 17776 24052
rect 17451 24021 17463 24024
rect 17405 24015 17463 24021
rect 17770 24012 17776 24024
rect 17828 24012 17834 24064
rect 17880 24052 17908 24219
rect 18432 24197 18460 24296
rect 18601 24327 18659 24333
rect 18601 24293 18613 24327
rect 18647 24324 18659 24327
rect 19150 24324 19156 24336
rect 18647 24296 19156 24324
rect 18647 24293 18659 24296
rect 18601 24287 18659 24293
rect 19150 24284 19156 24296
rect 19208 24324 19214 24336
rect 19352 24324 19380 24355
rect 19794 24352 19800 24364
rect 19852 24352 19858 24404
rect 21082 24352 21088 24404
rect 21140 24352 21146 24404
rect 21361 24395 21419 24401
rect 21361 24361 21373 24395
rect 21407 24392 21419 24395
rect 22370 24392 22376 24404
rect 21407 24364 22376 24392
rect 21407 24361 21419 24364
rect 21361 24355 21419 24361
rect 22370 24352 22376 24364
rect 22428 24352 22434 24404
rect 20990 24324 20996 24336
rect 19208 24296 19380 24324
rect 19444 24296 20996 24324
rect 19208 24284 19214 24296
rect 19242 24216 19248 24268
rect 19300 24216 19306 24268
rect 18417 24191 18475 24197
rect 18417 24157 18429 24191
rect 18463 24157 18475 24191
rect 18417 24151 18475 24157
rect 18601 24191 18659 24197
rect 18601 24157 18613 24191
rect 18647 24188 18659 24191
rect 18966 24188 18972 24200
rect 18647 24160 18972 24188
rect 18647 24157 18659 24160
rect 18601 24151 18659 24157
rect 18966 24148 18972 24160
rect 19024 24148 19030 24200
rect 19444 24182 19472 24296
rect 19886 24256 19892 24268
rect 19628 24228 19892 24256
rect 19628 24197 19656 24228
rect 19886 24216 19892 24228
rect 19944 24216 19950 24268
rect 20456 24265 20484 24296
rect 20990 24284 20996 24296
rect 21048 24284 21054 24336
rect 20441 24259 20499 24265
rect 20441 24225 20453 24259
rect 20487 24225 20499 24259
rect 20441 24219 20499 24225
rect 20533 24259 20591 24265
rect 20533 24225 20545 24259
rect 20579 24256 20591 24259
rect 20622 24256 20628 24268
rect 20579 24228 20628 24256
rect 20579 24225 20591 24228
rect 20533 24219 20591 24225
rect 19260 24154 19472 24182
rect 19613 24191 19671 24197
rect 19613 24157 19625 24191
rect 19659 24157 19671 24191
rect 17954 24080 17960 24132
rect 18012 24120 18018 24132
rect 19061 24123 19119 24129
rect 19061 24120 19073 24123
rect 18012 24092 19073 24120
rect 18012 24080 18018 24092
rect 19061 24089 19073 24092
rect 19107 24120 19119 24123
rect 19260 24120 19288 24154
rect 19613 24151 19671 24157
rect 19702 24148 19708 24200
rect 19760 24148 19766 24200
rect 19981 24191 20039 24197
rect 19981 24157 19993 24191
rect 20027 24188 20039 24191
rect 20070 24188 20076 24200
rect 20027 24160 20076 24188
rect 20027 24157 20039 24160
rect 19981 24151 20039 24157
rect 20070 24148 20076 24160
rect 20128 24148 20134 24200
rect 20257 24191 20315 24197
rect 20257 24157 20269 24191
rect 20303 24157 20315 24191
rect 20456 24188 20484 24219
rect 20622 24216 20628 24228
rect 20680 24216 20686 24268
rect 20717 24259 20775 24265
rect 20717 24225 20729 24259
rect 20763 24256 20775 24259
rect 21177 24259 21235 24265
rect 20763 24228 20944 24256
rect 20763 24225 20775 24228
rect 20717 24219 20775 24225
rect 20916 24200 20944 24228
rect 21177 24225 21189 24259
rect 21223 24256 21235 24259
rect 22922 24256 22928 24268
rect 21223 24228 22928 24256
rect 21223 24225 21235 24228
rect 21177 24219 21235 24225
rect 22922 24216 22928 24228
rect 22980 24216 22986 24268
rect 20809 24191 20867 24197
rect 20809 24188 20821 24191
rect 20456 24160 20821 24188
rect 20257 24151 20315 24157
rect 20809 24157 20821 24160
rect 20855 24157 20867 24191
rect 20809 24151 20867 24157
rect 20272 24120 20300 24151
rect 20898 24148 20904 24200
rect 20956 24148 20962 24200
rect 21085 24191 21143 24197
rect 21085 24157 21097 24191
rect 21131 24188 21143 24191
rect 21131 24160 21220 24188
rect 21131 24157 21143 24160
rect 21085 24151 21143 24157
rect 20916 24120 20944 24148
rect 21192 24129 21220 24160
rect 21266 24148 21272 24200
rect 21324 24188 21330 24200
rect 21453 24191 21511 24197
rect 21453 24188 21465 24191
rect 21324 24160 21465 24188
rect 21324 24148 21330 24160
rect 21453 24157 21465 24160
rect 21499 24157 21511 24191
rect 21453 24151 21511 24157
rect 21542 24148 21548 24200
rect 21600 24188 21606 24200
rect 23293 24191 23351 24197
rect 21600 24160 21942 24188
rect 21600 24148 21606 24160
rect 23293 24157 23305 24191
rect 23339 24157 23351 24191
rect 23293 24151 23351 24157
rect 19107 24092 19288 24120
rect 19444 24092 20944 24120
rect 21177 24123 21235 24129
rect 19107 24089 19119 24092
rect 19061 24083 19119 24089
rect 18598 24052 18604 24064
rect 17880 24024 18604 24052
rect 18598 24012 18604 24024
rect 18656 24012 18662 24064
rect 18861 24055 18919 24061
rect 18861 24021 18873 24055
rect 18907 24052 18919 24055
rect 19444 24052 19472 24092
rect 21177 24089 21189 24123
rect 21223 24089 21235 24123
rect 21177 24083 21235 24089
rect 23014 24080 23020 24132
rect 23072 24080 23078 24132
rect 18907 24024 19472 24052
rect 19521 24055 19579 24061
rect 18907 24021 18919 24024
rect 18861 24015 18919 24021
rect 19521 24021 19533 24055
rect 19567 24052 19579 24055
rect 19610 24052 19616 24064
rect 19567 24024 19616 24052
rect 19567 24021 19579 24024
rect 19521 24015 19579 24021
rect 19610 24012 19616 24024
rect 19668 24012 19674 24064
rect 19886 24012 19892 24064
rect 19944 24052 19950 24064
rect 20073 24055 20131 24061
rect 20073 24052 20085 24055
rect 19944 24024 20085 24052
rect 19944 24012 19950 24024
rect 20073 24021 20085 24024
rect 20119 24021 20131 24055
rect 20073 24015 20131 24021
rect 20162 24012 20168 24064
rect 20220 24052 20226 24064
rect 20533 24055 20591 24061
rect 20533 24052 20545 24055
rect 20220 24024 20545 24052
rect 20220 24012 20226 24024
rect 20533 24021 20545 24024
rect 20579 24021 20591 24055
rect 20533 24015 20591 24021
rect 21082 24012 21088 24064
rect 21140 24052 21146 24064
rect 21545 24055 21603 24061
rect 21545 24052 21557 24055
rect 21140 24024 21557 24052
rect 21140 24012 21146 24024
rect 21545 24021 21557 24024
rect 21591 24021 21603 24055
rect 21545 24015 21603 24021
rect 22738 24012 22744 24064
rect 22796 24052 22802 24064
rect 23308 24052 23336 24151
rect 22796 24024 23336 24052
rect 22796 24012 22802 24024
rect 1104 23962 25208 23984
rect 1104 23910 4874 23962
rect 4926 23910 4938 23962
rect 4990 23910 5002 23962
rect 5054 23910 5066 23962
rect 5118 23910 5130 23962
rect 5182 23910 25208 23962
rect 1104 23888 25208 23910
rect 1762 23808 1768 23860
rect 1820 23848 1826 23860
rect 1949 23851 2007 23857
rect 1949 23848 1961 23851
rect 1820 23820 1961 23848
rect 1820 23808 1826 23820
rect 1949 23817 1961 23820
rect 1995 23817 2007 23851
rect 1949 23811 2007 23817
rect 3234 23808 3240 23860
rect 3292 23848 3298 23860
rect 4157 23851 4215 23857
rect 4157 23848 4169 23851
rect 3292 23820 4169 23848
rect 3292 23808 3298 23820
rect 4157 23817 4169 23820
rect 4203 23817 4215 23851
rect 5813 23851 5871 23857
rect 5813 23848 5825 23851
rect 4157 23811 4215 23817
rect 4264 23820 5825 23848
rect 3326 23780 3332 23792
rect 2424 23752 3332 23780
rect 2424 23721 2452 23752
rect 3326 23740 3332 23752
rect 3384 23740 3390 23792
rect 4264 23780 4292 23820
rect 5813 23817 5825 23820
rect 5859 23817 5871 23851
rect 5813 23811 5871 23817
rect 7190 23808 7196 23860
rect 7248 23848 7254 23860
rect 7745 23851 7803 23857
rect 7745 23848 7757 23851
rect 7248 23820 7757 23848
rect 7248 23808 7254 23820
rect 7745 23817 7757 23820
rect 7791 23817 7803 23851
rect 7745 23811 7803 23817
rect 3620 23752 4292 23780
rect 2133 23715 2191 23721
rect 2133 23681 2145 23715
rect 2179 23681 2191 23715
rect 2133 23675 2191 23681
rect 2409 23715 2467 23721
rect 2409 23681 2421 23715
rect 2455 23681 2467 23715
rect 2409 23675 2467 23681
rect 2148 23576 2176 23675
rect 2866 23672 2872 23724
rect 2924 23712 2930 23724
rect 3620 23721 3648 23752
rect 4522 23740 4528 23792
rect 4580 23780 4586 23792
rect 5537 23783 5595 23789
rect 4580 23752 5488 23780
rect 4580 23740 4586 23752
rect 3053 23715 3111 23721
rect 3053 23712 3065 23715
rect 2924 23684 3065 23712
rect 2924 23672 2930 23684
rect 3053 23681 3065 23684
rect 3099 23681 3111 23715
rect 3053 23675 3111 23681
rect 3605 23715 3663 23721
rect 3605 23681 3617 23715
rect 3651 23681 3663 23715
rect 3605 23675 3663 23681
rect 3694 23672 3700 23724
rect 3752 23672 3758 23724
rect 3878 23672 3884 23724
rect 3936 23672 3942 23724
rect 4065 23715 4123 23721
rect 4065 23681 4077 23715
rect 4111 23712 4123 23715
rect 4154 23712 4160 23724
rect 4111 23684 4160 23712
rect 4111 23681 4123 23684
rect 4065 23675 4123 23681
rect 4154 23672 4160 23684
rect 4212 23712 4218 23724
rect 4801 23715 4859 23721
rect 4801 23712 4813 23715
rect 4212 23684 4813 23712
rect 4212 23672 4218 23684
rect 4801 23681 4813 23684
rect 4847 23712 4859 23715
rect 5077 23715 5135 23721
rect 4847 23684 5028 23712
rect 4847 23681 4859 23684
rect 4801 23675 4859 23681
rect 2317 23647 2375 23653
rect 2317 23613 2329 23647
rect 2363 23644 2375 23647
rect 3418 23644 3424 23656
rect 2363 23616 3424 23644
rect 2363 23613 2375 23616
rect 2317 23607 2375 23613
rect 3418 23604 3424 23616
rect 3476 23604 3482 23656
rect 3712 23576 3740 23672
rect 3789 23647 3847 23653
rect 3789 23613 3801 23647
rect 3835 23644 3847 23647
rect 4246 23644 4252 23656
rect 3835 23616 4252 23644
rect 3835 23613 3847 23616
rect 3789 23607 3847 23613
rect 4246 23604 4252 23616
rect 4304 23644 4310 23656
rect 4614 23644 4620 23656
rect 4304 23616 4620 23644
rect 4304 23604 4310 23616
rect 4614 23604 4620 23616
rect 4672 23604 4678 23656
rect 4893 23647 4951 23653
rect 4893 23644 4905 23647
rect 4724 23616 4905 23644
rect 4724 23576 4752 23616
rect 4893 23613 4905 23616
rect 4939 23613 4951 23647
rect 5000 23644 5028 23684
rect 5077 23681 5089 23715
rect 5123 23712 5135 23715
rect 5166 23712 5172 23724
rect 5123 23684 5172 23712
rect 5123 23681 5135 23684
rect 5077 23675 5135 23681
rect 5166 23672 5172 23684
rect 5224 23672 5230 23724
rect 5353 23715 5411 23721
rect 5353 23681 5365 23715
rect 5399 23681 5411 23715
rect 5460 23712 5488 23752
rect 5537 23749 5549 23783
rect 5583 23780 5595 23783
rect 5583 23752 5948 23780
rect 5583 23749 5595 23752
rect 5537 23743 5595 23749
rect 5920 23721 5948 23752
rect 6914 23740 6920 23792
rect 6972 23740 6978 23792
rect 7653 23783 7711 23789
rect 7653 23780 7665 23783
rect 7116 23752 7665 23780
rect 7116 23724 7144 23752
rect 7653 23749 7665 23752
rect 7699 23749 7711 23783
rect 7653 23743 7711 23749
rect 5629 23715 5687 23721
rect 5629 23712 5641 23715
rect 5460 23684 5641 23712
rect 5353 23675 5411 23681
rect 5629 23681 5641 23684
rect 5675 23681 5687 23715
rect 5629 23675 5687 23681
rect 5905 23715 5963 23721
rect 5905 23681 5917 23715
rect 5951 23712 5963 23715
rect 5994 23712 6000 23724
rect 5951 23684 6000 23712
rect 5951 23681 5963 23684
rect 5905 23675 5963 23681
rect 5258 23644 5264 23656
rect 5000 23616 5264 23644
rect 4893 23607 4951 23613
rect 5258 23604 5264 23616
rect 5316 23604 5322 23656
rect 5368 23644 5396 23675
rect 5994 23672 6000 23684
rect 6052 23672 6058 23724
rect 7098 23672 7104 23724
rect 7156 23672 7162 23724
rect 7561 23715 7619 23721
rect 7561 23681 7573 23715
rect 7607 23681 7619 23715
rect 7760 23712 7788 23811
rect 11238 23808 11244 23860
rect 11296 23848 11302 23860
rect 12158 23848 12164 23860
rect 11296 23820 12164 23848
rect 11296 23808 11302 23820
rect 12158 23808 12164 23820
rect 12216 23808 12222 23860
rect 12618 23808 12624 23860
rect 12676 23848 12682 23860
rect 12805 23851 12863 23857
rect 12805 23848 12817 23851
rect 12676 23820 12817 23848
rect 12676 23808 12682 23820
rect 12805 23817 12817 23820
rect 12851 23817 12863 23851
rect 12805 23811 12863 23817
rect 12894 23808 12900 23860
rect 12952 23848 12958 23860
rect 15746 23848 15752 23860
rect 12952 23820 15752 23848
rect 12952 23808 12958 23820
rect 15746 23808 15752 23820
rect 15804 23808 15810 23860
rect 16574 23808 16580 23860
rect 16632 23848 16638 23860
rect 19242 23848 19248 23860
rect 16632 23820 19248 23848
rect 16632 23808 16638 23820
rect 19242 23808 19248 23820
rect 19300 23808 19306 23860
rect 20806 23848 20812 23860
rect 19444 23820 20812 23848
rect 11885 23783 11943 23789
rect 11885 23749 11897 23783
rect 11931 23780 11943 23783
rect 12986 23780 12992 23792
rect 11931 23752 12992 23780
rect 11931 23749 11943 23752
rect 11885 23743 11943 23749
rect 12986 23740 12992 23752
rect 13044 23740 13050 23792
rect 13354 23740 13360 23792
rect 13412 23780 13418 23792
rect 15102 23780 15108 23792
rect 13412 23752 15108 23780
rect 13412 23740 13418 23752
rect 15102 23740 15108 23752
rect 15160 23740 15166 23792
rect 17770 23780 17776 23792
rect 16684 23752 17776 23780
rect 8386 23712 8392 23724
rect 7760 23684 8392 23712
rect 7561 23675 7619 23681
rect 5368 23616 5488 23644
rect 2148 23548 2774 23576
rect 3712 23548 4752 23576
rect 2406 23468 2412 23520
rect 2464 23508 2470 23520
rect 2501 23511 2559 23517
rect 2501 23508 2513 23511
rect 2464 23480 2513 23508
rect 2464 23468 2470 23480
rect 2501 23477 2513 23480
rect 2547 23477 2559 23511
rect 2746 23508 2774 23548
rect 4798 23536 4804 23588
rect 4856 23576 4862 23588
rect 5353 23579 5411 23585
rect 5353 23576 5365 23579
rect 4856 23548 5365 23576
rect 4856 23536 4862 23548
rect 5353 23545 5365 23548
rect 5399 23545 5411 23579
rect 5353 23539 5411 23545
rect 4338 23508 4344 23520
rect 2746 23480 4344 23508
rect 2501 23471 2559 23477
rect 4338 23468 4344 23480
rect 4396 23468 4402 23520
rect 4706 23468 4712 23520
rect 4764 23508 4770 23520
rect 5261 23511 5319 23517
rect 5261 23508 5273 23511
rect 4764 23480 5273 23508
rect 4764 23468 4770 23480
rect 5261 23477 5273 23480
rect 5307 23508 5319 23511
rect 5460 23508 5488 23616
rect 6086 23604 6092 23656
rect 6144 23644 6150 23656
rect 7374 23644 7380 23656
rect 6144 23616 7380 23644
rect 6144 23604 6150 23616
rect 7374 23604 7380 23616
rect 7432 23644 7438 23656
rect 7576 23644 7604 23675
rect 8386 23672 8392 23684
rect 8444 23672 8450 23724
rect 11054 23672 11060 23724
rect 11112 23672 11118 23724
rect 11149 23715 11207 23721
rect 11149 23681 11161 23715
rect 11195 23681 11207 23715
rect 11149 23675 11207 23681
rect 7432 23616 7604 23644
rect 7432 23604 7438 23616
rect 7650 23604 7656 23656
rect 7708 23644 7714 23656
rect 7929 23647 7987 23653
rect 7929 23644 7941 23647
rect 7708 23616 7941 23644
rect 7708 23604 7714 23616
rect 7929 23613 7941 23616
rect 7975 23613 7987 23647
rect 11164 23644 11192 23675
rect 11790 23672 11796 23724
rect 11848 23672 11854 23724
rect 11977 23715 12035 23721
rect 11977 23681 11989 23715
rect 12023 23712 12035 23715
rect 12345 23715 12403 23721
rect 12345 23712 12357 23715
rect 12023 23684 12357 23712
rect 12023 23681 12035 23684
rect 11977 23675 12035 23681
rect 12345 23681 12357 23684
rect 12391 23681 12403 23715
rect 12345 23675 12403 23681
rect 12434 23672 12440 23724
rect 12492 23712 12498 23724
rect 12559 23715 12617 23721
rect 12559 23712 12571 23715
rect 12492 23684 12571 23712
rect 12492 23672 12498 23684
rect 12559 23681 12571 23684
rect 12605 23681 12617 23715
rect 12559 23675 12617 23681
rect 12713 23715 12771 23721
rect 12713 23681 12725 23715
rect 12759 23712 12771 23715
rect 12894 23712 12900 23724
rect 12759 23684 12900 23712
rect 12759 23681 12771 23684
rect 12713 23675 12771 23681
rect 12894 23672 12900 23684
rect 12952 23672 12958 23724
rect 13078 23672 13084 23724
rect 13136 23672 13142 23724
rect 16684 23721 16712 23752
rect 17770 23740 17776 23752
rect 17828 23740 17834 23792
rect 17862 23740 17868 23792
rect 17920 23740 17926 23792
rect 19150 23740 19156 23792
rect 19208 23740 19214 23792
rect 16669 23715 16727 23721
rect 16669 23681 16681 23715
rect 16715 23681 16727 23715
rect 16669 23675 16727 23681
rect 16942 23672 16948 23724
rect 17000 23672 17006 23724
rect 19058 23712 19064 23724
rect 18524 23684 19064 23712
rect 18524 23656 18552 23684
rect 19058 23672 19064 23684
rect 19116 23712 19122 23724
rect 19444 23721 19472 23820
rect 20806 23808 20812 23820
rect 20864 23808 20870 23860
rect 21082 23808 21088 23860
rect 21140 23848 21146 23860
rect 22281 23851 22339 23857
rect 21140 23820 22232 23848
rect 21140 23808 21146 23820
rect 19610 23740 19616 23792
rect 19668 23740 19674 23792
rect 19886 23740 19892 23792
rect 19944 23740 19950 23792
rect 20073 23783 20131 23789
rect 20073 23749 20085 23783
rect 20119 23780 20131 23783
rect 20162 23780 20168 23792
rect 20119 23752 20168 23780
rect 20119 23749 20131 23752
rect 20073 23743 20131 23749
rect 20162 23740 20168 23752
rect 20220 23740 20226 23792
rect 20990 23740 20996 23792
rect 21048 23780 21054 23792
rect 21269 23783 21327 23789
rect 21269 23780 21281 23783
rect 21048 23752 21281 23780
rect 21048 23740 21054 23752
rect 21269 23749 21281 23752
rect 21315 23780 21327 23783
rect 21358 23780 21364 23792
rect 21315 23752 21364 23780
rect 21315 23749 21327 23752
rect 21269 23743 21327 23749
rect 21358 23740 21364 23752
rect 21416 23740 21422 23792
rect 22204 23789 22232 23820
rect 22281 23817 22293 23851
rect 22327 23848 22339 23851
rect 22370 23848 22376 23860
rect 22327 23820 22376 23848
rect 22327 23817 22339 23820
rect 22281 23811 22339 23817
rect 22370 23808 22376 23820
rect 22428 23808 22434 23860
rect 22646 23808 22652 23860
rect 22704 23848 22710 23860
rect 23017 23851 23075 23857
rect 23017 23848 23029 23851
rect 22704 23820 23029 23848
rect 22704 23808 22710 23820
rect 23017 23817 23029 23820
rect 23063 23817 23075 23851
rect 23017 23811 23075 23817
rect 21989 23783 22047 23789
rect 21989 23749 22001 23783
rect 22035 23780 22047 23783
rect 22189 23783 22247 23789
rect 22035 23752 22140 23780
rect 22035 23749 22047 23752
rect 21989 23743 22047 23749
rect 19245 23715 19303 23721
rect 19245 23712 19257 23715
rect 19116 23684 19257 23712
rect 19116 23672 19122 23684
rect 19245 23681 19257 23684
rect 19291 23681 19303 23715
rect 19245 23675 19303 23681
rect 19429 23715 19487 23721
rect 19429 23681 19441 23715
rect 19475 23681 19487 23715
rect 19429 23675 19487 23681
rect 19521 23715 19579 23721
rect 19521 23681 19533 23715
rect 19567 23712 19579 23715
rect 19702 23712 19708 23724
rect 19567 23684 19708 23712
rect 19567 23681 19579 23684
rect 19521 23675 19579 23681
rect 19702 23672 19708 23684
rect 19760 23672 19766 23724
rect 19904 23712 19932 23740
rect 20349 23715 20407 23721
rect 20349 23712 20361 23715
rect 19904 23684 20361 23712
rect 20349 23681 20361 23684
rect 20395 23681 20407 23715
rect 20349 23675 20407 23681
rect 20441 23715 20499 23721
rect 20441 23681 20453 23715
rect 20487 23712 20499 23715
rect 21174 23712 21180 23724
rect 20487 23684 21180 23712
rect 20487 23681 20499 23684
rect 20441 23675 20499 23681
rect 12253 23647 12311 23653
rect 12253 23644 12265 23647
rect 11164 23616 12265 23644
rect 7929 23607 7987 23613
rect 12253 23613 12265 23616
rect 12299 23613 12311 23647
rect 12805 23647 12863 23653
rect 12805 23644 12817 23647
rect 12253 23607 12311 23613
rect 12360 23616 12817 23644
rect 7834 23536 7840 23588
rect 7892 23576 7898 23588
rect 8754 23576 8760 23588
rect 7892 23548 8760 23576
rect 7892 23536 7898 23548
rect 8754 23536 8760 23548
rect 8812 23536 8818 23588
rect 10873 23579 10931 23585
rect 10873 23545 10885 23579
rect 10919 23576 10931 23579
rect 11054 23576 11060 23588
rect 10919 23548 11060 23576
rect 10919 23545 10931 23548
rect 10873 23539 10931 23545
rect 11054 23536 11060 23548
rect 11112 23536 11118 23588
rect 11146 23536 11152 23588
rect 11204 23576 11210 23588
rect 11517 23579 11575 23585
rect 11517 23576 11529 23579
rect 11204 23548 11529 23576
rect 11204 23536 11210 23548
rect 11517 23545 11529 23548
rect 11563 23545 11575 23579
rect 11517 23539 11575 23545
rect 12158 23536 12164 23588
rect 12216 23536 12222 23588
rect 5307 23480 5488 23508
rect 5307 23477 5319 23480
rect 5261 23471 5319 23477
rect 7282 23468 7288 23520
rect 7340 23468 7346 23520
rect 7374 23468 7380 23520
rect 7432 23468 7438 23520
rect 8849 23511 8907 23517
rect 8849 23477 8861 23511
rect 8895 23508 8907 23511
rect 9030 23508 9036 23520
rect 8895 23480 9036 23508
rect 8895 23477 8907 23480
rect 8849 23471 8907 23477
rect 9030 23468 9036 23480
rect 9088 23468 9094 23520
rect 10686 23468 10692 23520
rect 10744 23468 10750 23520
rect 10965 23511 11023 23517
rect 10965 23477 10977 23511
rect 11011 23508 11023 23511
rect 11238 23508 11244 23520
rect 11011 23480 11244 23508
rect 11011 23477 11023 23480
rect 10965 23471 11023 23477
rect 11238 23468 11244 23480
rect 11296 23468 11302 23520
rect 12268 23508 12296 23607
rect 12360 23588 12388 23616
rect 12805 23613 12817 23616
rect 12851 23644 12863 23647
rect 14090 23644 14096 23656
rect 12851 23616 14096 23644
rect 12851 23613 12863 23616
rect 12805 23607 12863 23613
rect 14090 23604 14096 23616
rect 14148 23604 14154 23656
rect 15286 23604 15292 23656
rect 15344 23644 15350 23656
rect 17037 23647 17095 23653
rect 17037 23644 17049 23647
rect 15344 23616 17049 23644
rect 15344 23604 15350 23616
rect 17037 23613 17049 23616
rect 17083 23644 17095 23647
rect 18506 23644 18512 23656
rect 17083 23616 18512 23644
rect 17083 23613 17095 23616
rect 17037 23607 17095 23613
rect 18506 23604 18512 23616
rect 18564 23604 18570 23656
rect 18874 23604 18880 23656
rect 18932 23644 18938 23656
rect 19794 23644 19800 23656
rect 18932 23616 19800 23644
rect 18932 23604 18938 23616
rect 19794 23604 19800 23616
rect 19852 23604 19858 23656
rect 19886 23604 19892 23656
rect 19944 23644 19950 23656
rect 20165 23647 20223 23653
rect 20165 23644 20177 23647
rect 19944 23616 20177 23644
rect 19944 23604 19950 23616
rect 20165 23613 20177 23616
rect 20211 23644 20223 23647
rect 20622 23644 20628 23656
rect 20211 23616 20628 23644
rect 20211 23613 20223 23616
rect 20165 23607 20223 23613
rect 20622 23604 20628 23616
rect 20680 23604 20686 23656
rect 12342 23536 12348 23588
rect 12400 23536 12406 23588
rect 16761 23579 16819 23585
rect 16761 23576 16773 23579
rect 12912 23548 16773 23576
rect 12526 23508 12532 23520
rect 12268 23480 12532 23508
rect 12526 23468 12532 23480
rect 12584 23508 12590 23520
rect 12912 23508 12940 23548
rect 16761 23545 16773 23548
rect 16807 23576 16819 23579
rect 17678 23576 17684 23588
rect 16807 23548 17684 23576
rect 16807 23545 16819 23548
rect 16761 23539 16819 23545
rect 17678 23536 17684 23548
rect 17736 23536 17742 23588
rect 17770 23536 17776 23588
rect 17828 23576 17834 23588
rect 18141 23579 18199 23585
rect 18141 23576 18153 23579
rect 17828 23548 18153 23576
rect 17828 23536 17834 23548
rect 18141 23545 18153 23548
rect 18187 23545 18199 23579
rect 18414 23576 18420 23588
rect 18141 23539 18199 23545
rect 18248 23548 18420 23576
rect 12584 23480 12940 23508
rect 12989 23511 13047 23517
rect 12584 23468 12590 23480
rect 12989 23477 13001 23511
rect 13035 23508 13047 23511
rect 13262 23508 13268 23520
rect 13035 23480 13268 23508
rect 13035 23477 13047 23480
rect 12989 23471 13047 23477
rect 13262 23468 13268 23480
rect 13320 23468 13326 23520
rect 15102 23468 15108 23520
rect 15160 23508 15166 23520
rect 18248 23508 18276 23548
rect 18414 23536 18420 23548
rect 18472 23536 18478 23588
rect 18966 23536 18972 23588
rect 19024 23576 19030 23588
rect 20257 23579 20315 23585
rect 20257 23576 20269 23579
rect 19024 23548 20269 23576
rect 19024 23536 19030 23548
rect 20257 23545 20269 23548
rect 20303 23545 20315 23579
rect 20257 23539 20315 23545
rect 15160 23480 18276 23508
rect 15160 23468 15166 23480
rect 18322 23468 18328 23520
rect 18380 23468 18386 23520
rect 19334 23468 19340 23520
rect 19392 23508 19398 23520
rect 19705 23511 19763 23517
rect 19705 23508 19717 23511
rect 19392 23480 19717 23508
rect 19392 23468 19398 23480
rect 19705 23477 19717 23480
rect 19751 23477 19763 23511
rect 19705 23471 19763 23477
rect 19794 23468 19800 23520
rect 19852 23508 19858 23520
rect 20732 23508 20760 23684
rect 21174 23672 21180 23684
rect 21232 23672 21238 23724
rect 22112 23712 22140 23752
rect 22189 23749 22201 23783
rect 22235 23780 22247 23783
rect 22235 23752 22600 23780
rect 22235 23749 22247 23752
rect 22189 23743 22247 23749
rect 22278 23712 22284 23724
rect 22112 23684 22284 23712
rect 22278 23672 22284 23684
rect 22336 23712 22342 23724
rect 22572 23721 22600 23752
rect 22465 23715 22523 23721
rect 22465 23712 22477 23715
rect 22336 23684 22477 23712
rect 22336 23672 22342 23684
rect 22465 23681 22477 23684
rect 22511 23681 22523 23715
rect 22465 23675 22523 23681
rect 22557 23715 22615 23721
rect 22557 23681 22569 23715
rect 22603 23712 22615 23715
rect 22741 23715 22799 23721
rect 22741 23712 22753 23715
rect 22603 23684 22753 23712
rect 22603 23681 22615 23684
rect 22557 23675 22615 23681
rect 22741 23681 22753 23684
rect 22787 23681 22799 23715
rect 22741 23675 22799 23681
rect 20898 23604 20904 23656
rect 20956 23644 20962 23656
rect 20956 23616 21220 23644
rect 20956 23604 20962 23616
rect 20993 23579 21051 23585
rect 20993 23545 21005 23579
rect 21039 23576 21051 23579
rect 21082 23576 21088 23588
rect 21039 23548 21088 23576
rect 21039 23545 21051 23548
rect 20993 23539 21051 23545
rect 21082 23536 21088 23548
rect 21140 23536 21146 23588
rect 21192 23576 21220 23616
rect 21821 23579 21879 23585
rect 21821 23576 21833 23579
rect 21192 23548 21833 23576
rect 21821 23545 21833 23548
rect 21867 23545 21879 23579
rect 22480 23576 22508 23675
rect 22922 23604 22928 23656
rect 22980 23644 22986 23656
rect 23017 23647 23075 23653
rect 23017 23644 23029 23647
rect 22980 23616 23029 23644
rect 22980 23604 22986 23616
rect 23017 23613 23029 23616
rect 23063 23644 23075 23647
rect 23198 23644 23204 23656
rect 23063 23616 23204 23644
rect 23063 23613 23075 23616
rect 23017 23607 23075 23613
rect 23198 23604 23204 23616
rect 23256 23604 23262 23656
rect 22833 23579 22891 23585
rect 22833 23576 22845 23579
rect 22480 23548 22845 23576
rect 21821 23539 21879 23545
rect 22833 23545 22845 23548
rect 22879 23545 22891 23579
rect 22833 23539 22891 23545
rect 19852 23480 20760 23508
rect 19852 23468 19858 23480
rect 20806 23468 20812 23520
rect 20864 23468 20870 23520
rect 21266 23468 21272 23520
rect 21324 23508 21330 23520
rect 22005 23511 22063 23517
rect 22005 23508 22017 23511
rect 21324 23480 22017 23508
rect 21324 23468 21330 23480
rect 22005 23477 22017 23480
rect 22051 23477 22063 23511
rect 22005 23471 22063 23477
rect 1104 23418 25208 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 25208 23418
rect 1104 23344 25208 23366
rect 3878 23264 3884 23316
rect 3936 23304 3942 23316
rect 4525 23307 4583 23313
rect 4525 23304 4537 23307
rect 3936 23276 4537 23304
rect 3936 23264 3942 23276
rect 4525 23273 4537 23276
rect 4571 23273 4583 23307
rect 4525 23267 4583 23273
rect 4709 23307 4767 23313
rect 4709 23273 4721 23307
rect 4755 23304 4767 23307
rect 5166 23304 5172 23316
rect 4755 23276 5172 23304
rect 4755 23273 4767 23276
rect 4709 23267 4767 23273
rect 5166 23264 5172 23276
rect 5224 23264 5230 23316
rect 7282 23264 7288 23316
rect 7340 23304 7346 23316
rect 7745 23307 7803 23313
rect 7745 23304 7757 23307
rect 7340 23276 7757 23304
rect 7340 23264 7346 23276
rect 7745 23273 7757 23276
rect 7791 23273 7803 23307
rect 7745 23267 7803 23273
rect 9582 23264 9588 23316
rect 9640 23304 9646 23316
rect 9640 23276 11008 23304
rect 9640 23264 9646 23276
rect 2774 23236 2780 23248
rect 2746 23196 2780 23236
rect 2832 23196 2838 23248
rect 8386 23196 8392 23248
rect 8444 23236 8450 23248
rect 8573 23239 8631 23245
rect 8573 23236 8585 23239
rect 8444 23208 8585 23236
rect 8444 23196 8450 23208
rect 8573 23205 8585 23208
rect 8619 23205 8631 23239
rect 9125 23239 9183 23245
rect 9125 23236 9137 23239
rect 8573 23199 8631 23205
rect 8680 23208 9137 23236
rect 1673 23171 1731 23177
rect 1673 23137 1685 23171
rect 1719 23168 1731 23171
rect 2746 23168 2774 23196
rect 1719 23140 2774 23168
rect 1719 23137 1731 23140
rect 1673 23131 1731 23137
rect 7098 23128 7104 23180
rect 7156 23168 7162 23180
rect 8680 23168 8708 23208
rect 9125 23205 9137 23208
rect 9171 23236 9183 23239
rect 9766 23236 9772 23248
rect 9171 23208 9772 23236
rect 9171 23205 9183 23208
rect 9125 23199 9183 23205
rect 9766 23196 9772 23208
rect 9824 23196 9830 23248
rect 10980 23245 11008 23276
rect 11054 23264 11060 23316
rect 11112 23264 11118 23316
rect 11238 23264 11244 23316
rect 11296 23264 11302 23316
rect 12158 23264 12164 23316
rect 12216 23304 12222 23316
rect 12526 23304 12532 23316
rect 12216 23276 12532 23304
rect 12216 23264 12222 23276
rect 12526 23264 12532 23276
rect 12584 23264 12590 23316
rect 14090 23264 14096 23316
rect 14148 23304 14154 23316
rect 14918 23304 14924 23316
rect 14148 23276 14924 23304
rect 14148 23264 14154 23276
rect 14918 23264 14924 23276
rect 14976 23264 14982 23316
rect 15930 23264 15936 23316
rect 15988 23304 15994 23316
rect 16025 23307 16083 23313
rect 16025 23304 16037 23307
rect 15988 23276 16037 23304
rect 15988 23264 15994 23276
rect 16025 23273 16037 23276
rect 16071 23304 16083 23307
rect 16666 23304 16672 23316
rect 16071 23276 16672 23304
rect 16071 23273 16083 23276
rect 16025 23267 16083 23273
rect 16666 23264 16672 23276
rect 16724 23264 16730 23316
rect 16942 23264 16948 23316
rect 17000 23264 17006 23316
rect 17313 23307 17371 23313
rect 17313 23273 17325 23307
rect 17359 23304 17371 23307
rect 20806 23304 20812 23316
rect 17359 23276 20812 23304
rect 17359 23273 17371 23276
rect 17313 23267 17371 23273
rect 20806 23264 20812 23276
rect 20864 23264 20870 23316
rect 10965 23239 11023 23245
rect 10965 23205 10977 23239
rect 11011 23236 11023 23239
rect 11425 23239 11483 23245
rect 11011 23208 11192 23236
rect 11011 23205 11023 23208
rect 10965 23199 11023 23205
rect 7156 23140 8708 23168
rect 8757 23171 8815 23177
rect 7156 23128 7162 23140
rect 8757 23137 8769 23171
rect 8803 23168 8815 23171
rect 10318 23168 10324 23180
rect 8803 23140 10324 23168
rect 8803 23137 8815 23140
rect 8757 23131 8815 23137
rect 10318 23128 10324 23140
rect 10376 23128 10382 23180
rect 10413 23171 10471 23177
rect 10413 23137 10425 23171
rect 10459 23168 10471 23171
rect 11054 23168 11060 23180
rect 10459 23140 11060 23168
rect 10459 23137 10471 23140
rect 10413 23131 10471 23137
rect 11054 23128 11060 23140
rect 11112 23128 11118 23180
rect 1394 23060 1400 23112
rect 1452 23060 1458 23112
rect 2774 23060 2780 23112
rect 2832 23060 2838 23112
rect 4154 23060 4160 23112
rect 4212 23060 4218 23112
rect 4614 23060 4620 23112
rect 4672 23060 4678 23112
rect 7374 23060 7380 23112
rect 7432 23060 7438 23112
rect 8662 23100 8668 23112
rect 7760 23072 8668 23100
rect 2958 22992 2964 23044
rect 3016 23032 3022 23044
rect 3421 23035 3479 23041
rect 3421 23032 3433 23035
rect 3016 23004 3433 23032
rect 3016 22992 3022 23004
rect 3421 23001 3433 23004
rect 3467 23001 3479 23035
rect 3421 22995 3479 23001
rect 3436 22964 3464 22995
rect 3510 22992 3516 23044
rect 3568 23032 3574 23044
rect 3789 23035 3847 23041
rect 3789 23032 3801 23035
rect 3568 23004 3801 23032
rect 3568 22992 3574 23004
rect 3789 23001 3801 23004
rect 3835 23001 3847 23035
rect 3789 22995 3847 23001
rect 4341 23035 4399 23041
rect 4341 23001 4353 23035
rect 4387 23032 4399 23035
rect 4632 23032 4660 23060
rect 7760 23041 7788 23072
rect 8662 23060 8668 23072
rect 8720 23060 8726 23112
rect 10229 23103 10287 23109
rect 10229 23069 10241 23103
rect 10275 23100 10287 23103
rect 10686 23100 10692 23112
rect 10275 23072 10692 23100
rect 10275 23069 10287 23072
rect 10229 23063 10287 23069
rect 10686 23060 10692 23072
rect 10744 23060 10750 23112
rect 4387 23004 4660 23032
rect 7745 23035 7803 23041
rect 4387 23001 4399 23004
rect 4341 22995 4399 23001
rect 7745 23001 7757 23035
rect 7791 23001 7803 23035
rect 7745 22995 7803 23001
rect 8297 23035 8355 23041
rect 8297 23001 8309 23035
rect 8343 23032 8355 23035
rect 8754 23032 8760 23044
rect 8343 23004 8760 23032
rect 8343 23001 8355 23004
rect 8297 22995 8355 23001
rect 3602 22964 3608 22976
rect 3436 22936 3608 22964
rect 3602 22924 3608 22936
rect 3660 22924 3666 22976
rect 3804 22964 3832 22995
rect 8754 22992 8760 23004
rect 8812 23032 8818 23044
rect 9306 23032 9312 23044
rect 8812 23004 9312 23032
rect 8812 22992 8818 23004
rect 9306 22992 9312 23004
rect 9364 22992 9370 23044
rect 9490 22992 9496 23044
rect 9548 22992 9554 23044
rect 9674 22992 9680 23044
rect 9732 23032 9738 23044
rect 10137 23035 10195 23041
rect 10137 23032 10149 23035
rect 9732 23004 10149 23032
rect 9732 22992 9738 23004
rect 10137 23001 10149 23004
rect 10183 23001 10195 23035
rect 10137 22995 10195 23001
rect 10597 23035 10655 23041
rect 10597 23001 10609 23035
rect 10643 23001 10655 23035
rect 10597 22995 10655 23001
rect 4541 22967 4599 22973
rect 4541 22964 4553 22967
rect 3804 22936 4553 22964
rect 4541 22933 4553 22936
rect 4587 22933 4599 22967
rect 4541 22927 4599 22933
rect 7929 22967 7987 22973
rect 7929 22933 7941 22967
rect 7975 22964 7987 22967
rect 8386 22964 8392 22976
rect 7975 22936 8392 22964
rect 7975 22933 7987 22936
rect 7929 22927 7987 22933
rect 8386 22924 8392 22936
rect 8444 22924 8450 22976
rect 9033 22967 9091 22973
rect 9033 22933 9045 22967
rect 9079 22964 9091 22967
rect 9122 22964 9128 22976
rect 9079 22936 9128 22964
rect 9079 22933 9091 22936
rect 9033 22927 9091 22933
rect 9122 22924 9128 22936
rect 9180 22924 9186 22976
rect 9858 22924 9864 22976
rect 9916 22924 9922 22976
rect 10042 22924 10048 22976
rect 10100 22924 10106 22976
rect 10612 22964 10640 22995
rect 10686 22964 10692 22976
rect 10612 22936 10692 22964
rect 10686 22924 10692 22936
rect 10744 22924 10750 22976
rect 11164 22964 11192 23208
rect 11425 23205 11437 23239
rect 11471 23236 11483 23239
rect 12802 23236 12808 23248
rect 11471 23208 12808 23236
rect 11471 23205 11483 23208
rect 11425 23199 11483 23205
rect 12802 23196 12808 23208
rect 12860 23196 12866 23248
rect 12986 23196 12992 23248
rect 13044 23196 13050 23248
rect 16758 23196 16764 23248
rect 16816 23196 16822 23248
rect 16960 23236 16988 23264
rect 17957 23239 18015 23245
rect 17957 23236 17969 23239
rect 16960 23208 17969 23236
rect 17957 23205 17969 23208
rect 18003 23205 18015 23239
rect 17957 23199 18015 23205
rect 14093 23171 14151 23177
rect 14093 23168 14105 23171
rect 13218 23140 14105 23168
rect 11422 23060 11428 23112
rect 11480 23100 11486 23112
rect 11701 23103 11759 23109
rect 11701 23100 11713 23103
rect 11480 23072 11713 23100
rect 11480 23060 11486 23072
rect 11701 23069 11713 23072
rect 11747 23100 11759 23103
rect 12434 23100 12440 23112
rect 11747 23072 12440 23100
rect 11747 23069 11759 23072
rect 11701 23063 11759 23069
rect 12434 23060 12440 23072
rect 12492 23060 12498 23112
rect 12894 23060 12900 23112
rect 12952 23100 12958 23112
rect 13218 23109 13246 23140
rect 14093 23137 14105 23140
rect 14139 23168 14151 23171
rect 14182 23168 14188 23180
rect 14139 23140 14188 23168
rect 14139 23137 14151 23140
rect 14093 23131 14151 23137
rect 14182 23128 14188 23140
rect 14240 23128 14246 23180
rect 14826 23168 14832 23180
rect 14476 23140 14832 23168
rect 14476 23112 14504 23140
rect 14826 23128 14832 23140
rect 14884 23128 14890 23180
rect 15470 23128 15476 23180
rect 15528 23168 15534 23180
rect 15841 23171 15899 23177
rect 15841 23168 15853 23171
rect 15528 23140 15853 23168
rect 15528 23128 15534 23140
rect 15841 23137 15853 23140
rect 15887 23137 15899 23171
rect 15841 23131 15899 23137
rect 16945 23171 17003 23177
rect 16945 23137 16957 23171
rect 16991 23168 17003 23171
rect 17497 23171 17555 23177
rect 17497 23168 17509 23171
rect 16991 23140 17509 23168
rect 16991 23137 17003 23140
rect 16945 23131 17003 23137
rect 17497 23137 17509 23140
rect 17543 23137 17555 23171
rect 17497 23131 17555 23137
rect 18325 23171 18383 23177
rect 18325 23137 18337 23171
rect 18371 23168 18383 23171
rect 18874 23168 18880 23180
rect 18371 23140 18880 23168
rect 18371 23137 18383 23140
rect 18325 23131 18383 23137
rect 18874 23128 18880 23140
rect 18932 23128 18938 23180
rect 13203 23103 13261 23109
rect 13203 23102 13215 23103
rect 13112 23100 13215 23102
rect 12952 23074 13215 23100
rect 12952 23072 13140 23074
rect 12952 23060 12958 23072
rect 13203 23069 13215 23074
rect 13249 23069 13261 23103
rect 13203 23063 13261 23069
rect 13357 23103 13415 23109
rect 13357 23069 13369 23103
rect 13403 23100 13415 23103
rect 13538 23100 13544 23112
rect 13403 23072 13544 23100
rect 13403 23069 13415 23072
rect 13357 23063 13415 23069
rect 13538 23060 13544 23072
rect 13596 23060 13602 23112
rect 14458 23060 14464 23112
rect 14516 23060 14522 23112
rect 15930 23060 15936 23112
rect 15988 23060 15994 23112
rect 17402 23060 17408 23112
rect 17460 23060 17466 23112
rect 17589 23103 17647 23109
rect 17589 23069 17601 23103
rect 17635 23100 17647 23103
rect 17678 23100 17684 23112
rect 17635 23072 17684 23100
rect 17635 23069 17647 23072
rect 17589 23063 17647 23069
rect 17678 23060 17684 23072
rect 17736 23060 17742 23112
rect 17773 23103 17831 23109
rect 17773 23069 17785 23103
rect 17819 23100 17831 23103
rect 17862 23100 17868 23112
rect 17819 23072 17868 23100
rect 17819 23069 17831 23072
rect 17773 23063 17831 23069
rect 17862 23060 17868 23072
rect 17920 23060 17926 23112
rect 14274 23032 14280 23044
rect 12406 23004 14280 23032
rect 12406 22964 12434 23004
rect 14274 22992 14280 23004
rect 14332 22992 14338 23044
rect 15565 23035 15623 23041
rect 15565 23001 15577 23035
rect 15611 23001 15623 23035
rect 15565 22995 15623 23001
rect 11164 22936 12434 22964
rect 13446 22924 13452 22976
rect 13504 22964 13510 22976
rect 15580 22964 15608 22995
rect 16482 22992 16488 23044
rect 16540 22992 16546 23044
rect 13504 22936 15608 22964
rect 17037 22967 17095 22973
rect 13504 22924 13510 22936
rect 17037 22933 17049 22967
rect 17083 22964 17095 22967
rect 17126 22964 17132 22976
rect 17083 22936 17132 22964
rect 17083 22933 17095 22936
rect 17037 22927 17095 22933
rect 17126 22924 17132 22936
rect 17184 22924 17190 22976
rect 17865 22967 17923 22973
rect 17865 22933 17877 22967
rect 17911 22964 17923 22967
rect 17954 22964 17960 22976
rect 17911 22936 17960 22964
rect 17911 22933 17923 22936
rect 17865 22927 17923 22933
rect 17954 22924 17960 22936
rect 18012 22924 18018 22976
rect 1104 22874 25208 22896
rect 1104 22822 4874 22874
rect 4926 22822 4938 22874
rect 4990 22822 5002 22874
rect 5054 22822 5066 22874
rect 5118 22822 5130 22874
rect 5182 22822 25208 22874
rect 1104 22800 25208 22822
rect 3605 22763 3663 22769
rect 3605 22729 3617 22763
rect 3651 22760 3663 22763
rect 3878 22760 3884 22772
rect 3651 22732 3884 22760
rect 3651 22729 3663 22732
rect 3605 22723 3663 22729
rect 3878 22720 3884 22732
rect 3936 22720 3942 22772
rect 6365 22763 6423 22769
rect 6365 22729 6377 22763
rect 6411 22760 6423 22763
rect 7098 22760 7104 22772
rect 6411 22732 7104 22760
rect 6411 22729 6423 22732
rect 6365 22723 6423 22729
rect 7098 22720 7104 22732
rect 7156 22720 7162 22772
rect 9490 22720 9496 22772
rect 9548 22760 9554 22772
rect 9548 22732 9812 22760
rect 9548 22720 9554 22732
rect 2133 22695 2191 22701
rect 2133 22661 2145 22695
rect 2179 22692 2191 22695
rect 2406 22692 2412 22704
rect 2179 22664 2412 22692
rect 2179 22661 2191 22664
rect 2133 22655 2191 22661
rect 2406 22652 2412 22664
rect 2464 22652 2470 22704
rect 3142 22652 3148 22704
rect 3200 22652 3206 22704
rect 6178 22652 6184 22704
rect 6236 22692 6242 22704
rect 9309 22695 9367 22701
rect 6236 22664 6670 22692
rect 6236 22652 6242 22664
rect 9309 22661 9321 22695
rect 9355 22692 9367 22695
rect 9674 22692 9680 22704
rect 9355 22664 9680 22692
rect 9355 22661 9367 22664
rect 9309 22655 9367 22661
rect 9674 22652 9680 22664
rect 9732 22652 9738 22704
rect 9784 22692 9812 22732
rect 10042 22720 10048 22772
rect 10100 22760 10106 22772
rect 10137 22763 10195 22769
rect 10137 22760 10149 22763
rect 10100 22732 10149 22760
rect 10100 22720 10106 22732
rect 10137 22729 10149 22732
rect 10183 22729 10195 22763
rect 10137 22723 10195 22729
rect 12526 22720 12532 22772
rect 12584 22760 12590 22772
rect 12986 22760 12992 22772
rect 12584 22732 12992 22760
rect 12584 22720 12590 22732
rect 12986 22720 12992 22732
rect 13044 22720 13050 22772
rect 13170 22720 13176 22772
rect 13228 22760 13234 22772
rect 13722 22760 13728 22772
rect 13228 22732 13728 22760
rect 13228 22720 13234 22732
rect 13722 22720 13728 22732
rect 13780 22760 13786 22772
rect 14343 22763 14401 22769
rect 14343 22760 14355 22763
rect 13780 22732 14355 22760
rect 13780 22720 13786 22732
rect 14343 22729 14355 22732
rect 14389 22729 14401 22763
rect 14343 22723 14401 22729
rect 15565 22763 15623 22769
rect 15565 22729 15577 22763
rect 15611 22760 15623 22763
rect 16022 22760 16028 22772
rect 15611 22732 16028 22760
rect 15611 22729 15623 22732
rect 15565 22723 15623 22729
rect 16022 22720 16028 22732
rect 16080 22760 16086 22772
rect 16298 22760 16304 22772
rect 16080 22732 16304 22760
rect 16080 22720 16086 22732
rect 16298 22720 16304 22732
rect 16356 22720 16362 22772
rect 17402 22720 17408 22772
rect 17460 22720 17466 22772
rect 22449 22763 22507 22769
rect 22449 22729 22461 22763
rect 22495 22760 22507 22763
rect 23106 22760 23112 22772
rect 22495 22732 23112 22760
rect 22495 22729 22507 22732
rect 22449 22723 22507 22729
rect 23106 22720 23112 22732
rect 23164 22720 23170 22772
rect 11882 22692 11888 22704
rect 9784 22664 11888 22692
rect 11882 22652 11888 22664
rect 11940 22652 11946 22704
rect 12894 22652 12900 22704
rect 12952 22692 12958 22704
rect 13449 22695 13507 22701
rect 13449 22692 13461 22695
rect 12952 22664 13461 22692
rect 12952 22652 12958 22664
rect 13449 22661 13461 22664
rect 13495 22661 13507 22695
rect 13449 22655 13507 22661
rect 13814 22652 13820 22704
rect 13872 22692 13878 22704
rect 13872 22664 14412 22692
rect 13872 22652 13878 22664
rect 8110 22584 8116 22636
rect 8168 22584 8174 22636
rect 8754 22584 8760 22636
rect 8812 22584 8818 22636
rect 8846 22584 8852 22636
rect 8904 22584 8910 22636
rect 9030 22584 9036 22636
rect 9088 22584 9094 22636
rect 9122 22584 9128 22636
rect 9180 22584 9186 22636
rect 9398 22584 9404 22636
rect 9456 22584 9462 22636
rect 9582 22584 9588 22636
rect 9640 22584 9646 22636
rect 9766 22584 9772 22636
rect 9824 22584 9830 22636
rect 9953 22627 10011 22633
rect 9953 22593 9965 22627
rect 9999 22593 10011 22627
rect 9953 22587 10011 22593
rect 10413 22627 10471 22633
rect 10413 22593 10425 22627
rect 10459 22624 10471 22627
rect 10686 22624 10692 22636
rect 10459 22596 10692 22624
rect 10459 22593 10471 22596
rect 10413 22587 10471 22593
rect 1394 22516 1400 22568
rect 1452 22556 1458 22568
rect 1857 22559 1915 22565
rect 1857 22556 1869 22559
rect 1452 22528 1869 22556
rect 1452 22516 1458 22528
rect 1857 22525 1869 22528
rect 1903 22525 1915 22559
rect 1857 22519 1915 22525
rect 7837 22559 7895 22565
rect 7837 22525 7849 22559
rect 7883 22556 7895 22559
rect 8386 22556 8392 22568
rect 7883 22528 8392 22556
rect 7883 22525 7895 22528
rect 7837 22519 7895 22525
rect 8386 22516 8392 22528
rect 8444 22556 8450 22568
rect 9214 22556 9220 22568
rect 8444 22528 9220 22556
rect 8444 22516 8450 22528
rect 9214 22516 9220 22528
rect 9272 22516 9278 22568
rect 9677 22559 9735 22565
rect 9677 22525 9689 22559
rect 9723 22525 9735 22559
rect 9968 22556 9996 22587
rect 10686 22584 10692 22596
rect 10744 22584 10750 22636
rect 12158 22584 12164 22636
rect 12216 22584 12222 22636
rect 12250 22584 12256 22636
rect 12308 22584 12314 22636
rect 12345 22627 12403 22633
rect 12345 22593 12357 22627
rect 12391 22624 12403 22627
rect 12526 22624 12532 22636
rect 12391 22596 12532 22624
rect 12391 22593 12403 22596
rect 12345 22587 12403 22593
rect 12526 22584 12532 22596
rect 12584 22584 12590 22636
rect 13170 22584 13176 22636
rect 13228 22584 13234 22636
rect 13265 22627 13323 22633
rect 13265 22593 13277 22627
rect 13311 22624 13323 22627
rect 13311 22596 13952 22624
rect 13311 22593 13323 22596
rect 13265 22587 13323 22593
rect 10502 22556 10508 22568
rect 9968 22528 10508 22556
rect 9677 22519 9735 22525
rect 9692 22488 9720 22519
rect 10502 22516 10508 22528
rect 10560 22516 10566 22568
rect 12710 22516 12716 22568
rect 12768 22556 12774 22568
rect 13280 22556 13308 22587
rect 13817 22559 13875 22565
rect 13817 22556 13829 22559
rect 12768 22528 13308 22556
rect 13648 22528 13829 22556
rect 12768 22516 12774 22528
rect 10321 22491 10379 22497
rect 10321 22488 10333 22491
rect 9692 22460 10333 22488
rect 10321 22457 10333 22460
rect 10367 22457 10379 22491
rect 10321 22451 10379 22457
rect 10428 22460 12112 22488
rect 8938 22380 8944 22432
rect 8996 22380 9002 22432
rect 9306 22380 9312 22432
rect 9364 22420 9370 22432
rect 10428 22420 10456 22460
rect 9364 22392 10456 22420
rect 9364 22380 9370 22392
rect 11974 22380 11980 22432
rect 12032 22380 12038 22432
rect 12084 22420 12112 22460
rect 12434 22448 12440 22500
rect 12492 22488 12498 22500
rect 12529 22491 12587 22497
rect 12529 22488 12541 22491
rect 12492 22460 12541 22488
rect 12492 22448 12498 22460
rect 12529 22457 12541 22460
rect 12575 22457 12587 22491
rect 12529 22451 12587 22457
rect 13449 22491 13507 22497
rect 13449 22457 13461 22491
rect 13495 22488 13507 22491
rect 13648 22488 13676 22528
rect 13817 22525 13829 22528
rect 13863 22525 13875 22559
rect 13924 22556 13952 22596
rect 14090 22584 14096 22636
rect 14148 22584 14154 22636
rect 14384 22624 14412 22664
rect 14458 22652 14464 22704
rect 14516 22692 14522 22704
rect 14553 22695 14611 22701
rect 14553 22692 14565 22695
rect 14516 22664 14565 22692
rect 14516 22652 14522 22664
rect 14553 22661 14565 22664
rect 14599 22692 14611 22695
rect 14734 22692 14740 22704
rect 14599 22664 14740 22692
rect 14599 22661 14611 22664
rect 14553 22655 14611 22661
rect 14734 22652 14740 22664
rect 14792 22652 14798 22704
rect 15930 22652 15936 22704
rect 15988 22692 15994 22704
rect 16945 22695 17003 22701
rect 16945 22692 16957 22695
rect 15988 22664 16957 22692
rect 15988 22652 15994 22664
rect 16945 22661 16957 22664
rect 16991 22692 17003 22695
rect 17494 22692 17500 22704
rect 16991 22664 17500 22692
rect 16991 22661 17003 22664
rect 16945 22655 17003 22661
rect 17494 22652 17500 22664
rect 17552 22652 17558 22704
rect 20990 22652 20996 22704
rect 21048 22692 21054 22704
rect 22649 22695 22707 22701
rect 22649 22692 22661 22695
rect 21048 22664 21220 22692
rect 21048 22652 21054 22664
rect 15473 22627 15531 22633
rect 15473 22624 15485 22627
rect 14384 22596 15485 22624
rect 15473 22593 15485 22596
rect 15519 22624 15531 22627
rect 16758 22624 16764 22636
rect 15519 22596 16764 22624
rect 15519 22593 15531 22596
rect 15473 22587 15531 22593
rect 16758 22584 16764 22596
rect 16816 22584 16822 22636
rect 21082 22584 21088 22636
rect 21140 22584 21146 22636
rect 21192 22633 21220 22664
rect 21929 22664 22661 22692
rect 21178 22627 21236 22633
rect 21178 22593 21190 22627
rect 21224 22593 21236 22627
rect 21178 22587 21236 22593
rect 21726 22584 21732 22636
rect 21784 22624 21790 22636
rect 21929 22633 21957 22664
rect 22649 22661 22661 22664
rect 22695 22692 22707 22695
rect 23014 22692 23020 22704
rect 22695 22664 23020 22692
rect 22695 22661 22707 22664
rect 22649 22655 22707 22661
rect 23014 22652 23020 22664
rect 23072 22652 23078 22704
rect 21821 22627 21879 22633
rect 21821 22624 21833 22627
rect 21784 22596 21833 22624
rect 21784 22584 21790 22596
rect 21821 22593 21833 22596
rect 21867 22593 21879 22627
rect 21821 22587 21879 22593
rect 21914 22627 21972 22633
rect 21914 22593 21926 22627
rect 21960 22593 21972 22627
rect 21914 22587 21972 22593
rect 14274 22556 14280 22568
rect 13924 22528 14280 22556
rect 13817 22519 13875 22525
rect 14274 22516 14280 22528
rect 14332 22516 14338 22568
rect 13495 22460 13676 22488
rect 13495 22457 13507 22460
rect 13449 22451 13507 22457
rect 16758 22448 16764 22500
rect 16816 22488 16822 22500
rect 17221 22491 17279 22497
rect 17221 22488 17233 22491
rect 16816 22460 17233 22488
rect 16816 22448 16822 22460
rect 17221 22457 17233 22460
rect 17267 22488 17279 22491
rect 17586 22488 17592 22500
rect 17267 22460 17592 22488
rect 17267 22457 17279 22460
rect 17221 22451 17279 22457
rect 17586 22448 17592 22460
rect 17644 22448 17650 22500
rect 21453 22491 21511 22497
rect 21453 22457 21465 22491
rect 21499 22488 21511 22491
rect 22094 22488 22100 22500
rect 21499 22460 22100 22488
rect 21499 22457 21511 22460
rect 21453 22451 21511 22457
rect 22094 22448 22100 22460
rect 22152 22448 22158 22500
rect 22186 22448 22192 22500
rect 22244 22448 22250 22500
rect 12986 22420 12992 22432
rect 12084 22392 12992 22420
rect 12986 22380 12992 22392
rect 13044 22380 13050 22432
rect 13538 22380 13544 22432
rect 13596 22380 13602 22432
rect 14001 22423 14059 22429
rect 14001 22389 14013 22423
rect 14047 22420 14059 22423
rect 14185 22423 14243 22429
rect 14185 22420 14197 22423
rect 14047 22392 14197 22420
rect 14047 22389 14059 22392
rect 14001 22383 14059 22389
rect 14185 22389 14197 22392
rect 14231 22389 14243 22423
rect 14185 22383 14243 22389
rect 14274 22380 14280 22432
rect 14332 22420 14338 22432
rect 14369 22423 14427 22429
rect 14369 22420 14381 22423
rect 14332 22392 14381 22420
rect 14332 22380 14338 22392
rect 14369 22389 14381 22392
rect 14415 22389 14427 22423
rect 14369 22383 14427 22389
rect 14918 22380 14924 22432
rect 14976 22420 14982 22432
rect 15930 22420 15936 22432
rect 14976 22392 15936 22420
rect 14976 22380 14982 22392
rect 15930 22380 15936 22392
rect 15988 22380 15994 22432
rect 22278 22380 22284 22432
rect 22336 22380 22342 22432
rect 22465 22423 22523 22429
rect 22465 22389 22477 22423
rect 22511 22420 22523 22423
rect 22830 22420 22836 22432
rect 22511 22392 22836 22420
rect 22511 22389 22523 22392
rect 22465 22383 22523 22389
rect 22830 22380 22836 22392
rect 22888 22380 22894 22432
rect 1104 22330 25208 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 25208 22330
rect 1104 22256 25208 22278
rect 8297 22219 8355 22225
rect 8297 22185 8309 22219
rect 8343 22216 8355 22219
rect 8938 22216 8944 22228
rect 8343 22188 8944 22216
rect 8343 22185 8355 22188
rect 8297 22179 8355 22185
rect 8938 22176 8944 22188
rect 8996 22176 9002 22228
rect 9950 22176 9956 22228
rect 10008 22216 10014 22228
rect 10502 22216 10508 22228
rect 10008 22188 10508 22216
rect 10008 22176 10014 22188
rect 10502 22176 10508 22188
rect 10560 22176 10566 22228
rect 11624 22188 12940 22216
rect 6365 22151 6423 22157
rect 6365 22117 6377 22151
rect 6411 22148 6423 22151
rect 8205 22151 8263 22157
rect 6411 22120 6868 22148
rect 6411 22117 6423 22120
rect 6365 22111 6423 22117
rect 5905 22083 5963 22089
rect 5905 22049 5917 22083
rect 5951 22080 5963 22083
rect 6840 22080 6868 22120
rect 8205 22117 8217 22151
rect 8251 22148 8263 22151
rect 8386 22148 8392 22160
rect 8251 22120 8392 22148
rect 8251 22117 8263 22120
rect 8205 22111 8263 22117
rect 8386 22108 8392 22120
rect 8444 22108 8450 22160
rect 8662 22080 8668 22092
rect 5951 22052 6776 22080
rect 6840 22052 8668 22080
rect 5951 22049 5963 22052
rect 5905 22043 5963 22049
rect 3602 21972 3608 22024
rect 3660 22012 3666 22024
rect 5629 22015 5687 22021
rect 5629 22012 5641 22015
rect 3660 21984 5641 22012
rect 3660 21972 3666 21984
rect 5629 21981 5641 21984
rect 5675 22012 5687 22015
rect 5994 22012 6000 22024
rect 5675 21984 6000 22012
rect 5675 21981 5687 21984
rect 5629 21975 5687 21981
rect 5994 21972 6000 21984
rect 6052 21972 6058 22024
rect 6181 22015 6239 22021
rect 6181 21981 6193 22015
rect 6227 22012 6239 22015
rect 6362 22012 6368 22024
rect 6227 21984 6368 22012
rect 6227 21981 6239 21984
rect 6181 21975 6239 21981
rect 6362 21972 6368 21984
rect 6420 21972 6426 22024
rect 6457 22015 6515 22021
rect 6457 21981 6469 22015
rect 6503 21981 6515 22015
rect 6457 21975 6515 21981
rect 5810 21904 5816 21956
rect 5868 21944 5874 21956
rect 6472 21944 6500 21975
rect 6546 21972 6552 22024
rect 6604 21972 6610 22024
rect 6748 22021 6776 22052
rect 8662 22040 8668 22052
rect 8720 22040 8726 22092
rect 9214 22040 9220 22092
rect 9272 22040 9278 22092
rect 9950 22040 9956 22092
rect 10008 22080 10014 22092
rect 11624 22080 11652 22188
rect 12066 22108 12072 22160
rect 12124 22148 12130 22160
rect 12710 22148 12716 22160
rect 12124 22120 12296 22148
rect 12124 22108 12130 22120
rect 10008 22052 11652 22080
rect 11977 22083 12035 22089
rect 10008 22040 10014 22052
rect 11977 22049 11989 22083
rect 12023 22080 12035 22083
rect 12158 22080 12164 22092
rect 12023 22052 12164 22080
rect 12023 22049 12035 22052
rect 11977 22043 12035 22049
rect 12158 22040 12164 22052
rect 12216 22040 12222 22092
rect 6733 22015 6791 22021
rect 6733 21981 6745 22015
rect 6779 22012 6791 22015
rect 9309 22015 9367 22021
rect 6779 21984 7972 22012
rect 6779 21981 6791 21984
rect 6733 21975 6791 21981
rect 5868 21916 6500 21944
rect 7837 21947 7895 21953
rect 5868 21904 5874 21916
rect 7837 21913 7849 21947
rect 7883 21913 7895 21947
rect 7944 21944 7972 21984
rect 9309 21981 9321 22015
rect 9355 22012 9367 22015
rect 9968 22012 9996 22040
rect 9355 21984 9996 22012
rect 9355 21981 9367 21984
rect 9309 21975 9367 21981
rect 10318 21972 10324 22024
rect 10376 22012 10382 22024
rect 11425 22015 11483 22021
rect 11425 22012 11437 22015
rect 10376 21984 11437 22012
rect 10376 21972 10382 21984
rect 11425 21981 11437 21984
rect 11471 21981 11483 22015
rect 11425 21975 11483 21981
rect 11514 21972 11520 22024
rect 11572 21972 11578 22024
rect 11785 22015 11843 22021
rect 11624 22010 11744 22014
rect 11785 22010 11797 22015
rect 11624 21986 11797 22010
rect 9858 21944 9864 21956
rect 7944 21916 9864 21944
rect 7837 21907 7895 21913
rect 5626 21836 5632 21888
rect 5684 21876 5690 21888
rect 6549 21879 6607 21885
rect 6549 21876 6561 21879
rect 5684 21848 6561 21876
rect 5684 21836 5690 21848
rect 6549 21845 6561 21848
rect 6595 21845 6607 21879
rect 6549 21839 6607 21845
rect 6914 21836 6920 21888
rect 6972 21876 6978 21888
rect 7852 21876 7880 21907
rect 9858 21904 9864 21916
rect 9916 21904 9922 21956
rect 10594 21904 10600 21956
rect 10652 21944 10658 21956
rect 11624 21944 11652 21986
rect 11716 21982 11797 21986
rect 11785 21981 11797 21982
rect 11831 21981 11843 22015
rect 11785 21975 11843 21981
rect 11882 21972 11888 22024
rect 11940 21972 11946 22024
rect 12066 21972 12072 22024
rect 12124 21972 12130 22024
rect 12268 22021 12296 22120
rect 12360 22120 12716 22148
rect 12360 22089 12388 22120
rect 12710 22108 12716 22120
rect 12768 22108 12774 22160
rect 12345 22083 12403 22089
rect 12345 22049 12357 22083
rect 12391 22049 12403 22083
rect 12345 22043 12403 22049
rect 12253 22015 12311 22021
rect 12253 21981 12265 22015
rect 12299 21981 12311 22015
rect 12253 21975 12311 21981
rect 10652 21916 11652 21944
rect 11701 21947 11759 21953
rect 10652 21904 10658 21916
rect 11701 21913 11713 21947
rect 11747 21944 11759 21947
rect 12268 21944 12296 21975
rect 11747 21916 12296 21944
rect 11747 21913 11759 21916
rect 11701 21907 11759 21913
rect 8570 21876 8576 21888
rect 6972 21848 8576 21876
rect 6972 21836 6978 21848
rect 8570 21836 8576 21848
rect 8628 21836 8634 21888
rect 9674 21836 9680 21888
rect 9732 21836 9738 21888
rect 11514 21836 11520 21888
rect 11572 21876 11578 21888
rect 12360 21876 12388 22043
rect 12526 22040 12532 22092
rect 12584 22080 12590 22092
rect 12805 22083 12863 22089
rect 12805 22080 12817 22083
rect 12584 22052 12817 22080
rect 12584 22040 12590 22052
rect 12805 22049 12817 22052
rect 12851 22049 12863 22083
rect 12912 22080 12940 22188
rect 12986 22176 12992 22228
rect 13044 22176 13050 22228
rect 13078 22176 13084 22228
rect 13136 22176 13142 22228
rect 13170 22176 13176 22228
rect 13228 22216 13234 22228
rect 13265 22219 13323 22225
rect 13265 22216 13277 22219
rect 13228 22188 13277 22216
rect 13228 22176 13234 22188
rect 13265 22185 13277 22188
rect 13311 22185 13323 22219
rect 15562 22216 15568 22228
rect 13265 22179 13323 22185
rect 13372 22188 15568 22216
rect 13004 22148 13032 22176
rect 13372 22148 13400 22188
rect 15562 22176 15568 22188
rect 15620 22176 15626 22228
rect 15749 22219 15807 22225
rect 15749 22185 15761 22219
rect 15795 22216 15807 22219
rect 15795 22188 17080 22216
rect 15795 22185 15807 22188
rect 15749 22179 15807 22185
rect 13004 22120 13400 22148
rect 13446 22108 13452 22160
rect 13504 22148 13510 22160
rect 13630 22148 13636 22160
rect 13504 22120 13636 22148
rect 13504 22108 13510 22120
rect 13630 22108 13636 22120
rect 13688 22148 13694 22160
rect 14918 22148 14924 22160
rect 13688 22120 14924 22148
rect 13688 22108 13694 22120
rect 14918 22108 14924 22120
rect 14976 22108 14982 22160
rect 15010 22108 15016 22160
rect 15068 22148 15074 22160
rect 15289 22151 15347 22157
rect 15289 22148 15301 22151
rect 15068 22120 15301 22148
rect 15068 22108 15074 22120
rect 15289 22117 15301 22120
rect 15335 22117 15347 22151
rect 15289 22111 15347 22117
rect 16206 22108 16212 22160
rect 16264 22108 16270 22160
rect 16853 22151 16911 22157
rect 16853 22148 16865 22151
rect 16684 22120 16865 22148
rect 12986 22080 12992 22092
rect 12912 22052 12992 22080
rect 12805 22043 12863 22049
rect 12986 22040 12992 22052
rect 13044 22040 13050 22092
rect 13078 22040 13084 22092
rect 13136 22080 13142 22092
rect 13262 22080 13268 22092
rect 13136 22052 13268 22080
rect 13136 22040 13142 22052
rect 13262 22040 13268 22052
rect 13320 22040 13326 22092
rect 13354 22040 13360 22092
rect 13412 22080 13418 22092
rect 13725 22083 13783 22089
rect 13725 22080 13737 22083
rect 13412 22052 13737 22080
rect 13412 22040 13418 22052
rect 13725 22049 13737 22052
rect 13771 22049 13783 22083
rect 13725 22043 13783 22049
rect 15197 22083 15255 22089
rect 15197 22049 15209 22083
rect 15243 22080 15255 22083
rect 16117 22083 16175 22089
rect 16117 22080 16129 22083
rect 15243 22052 16129 22080
rect 15243 22049 15255 22052
rect 15197 22043 15255 22049
rect 16117 22049 16129 22052
rect 16163 22049 16175 22083
rect 16577 22083 16635 22089
rect 16577 22080 16589 22083
rect 16117 22043 16175 22049
rect 16224 22052 16589 22080
rect 12437 22015 12495 22021
rect 12437 21981 12449 22015
rect 12483 22012 12495 22015
rect 12483 21984 12572 22012
rect 12483 21981 12495 21984
rect 12437 21975 12495 21981
rect 12544 21956 12572 21984
rect 12618 21972 12624 22024
rect 12676 22012 12682 22024
rect 13817 22015 13875 22021
rect 12676 21984 13308 22012
rect 12676 21972 12682 21984
rect 12526 21904 12532 21956
rect 12584 21944 12590 21956
rect 12897 21947 12955 21953
rect 12897 21944 12909 21947
rect 12584 21916 12909 21944
rect 12584 21904 12590 21916
rect 12897 21913 12909 21916
rect 12943 21913 12955 21947
rect 12897 21907 12955 21913
rect 11572 21848 12388 21876
rect 11572 21836 11578 21848
rect 12710 21836 12716 21888
rect 12768 21876 12774 21888
rect 13097 21879 13155 21885
rect 13097 21876 13109 21879
rect 12768 21848 13109 21876
rect 12768 21836 12774 21848
rect 13097 21845 13109 21848
rect 13143 21845 13155 21879
rect 13280 21876 13308 21984
rect 13817 21981 13829 22015
rect 13863 21981 13875 22015
rect 13817 21975 13875 21981
rect 13354 21904 13360 21956
rect 13412 21944 13418 21956
rect 13538 21944 13544 21956
rect 13412 21916 13544 21944
rect 13412 21904 13418 21916
rect 13538 21904 13544 21916
rect 13596 21944 13602 21956
rect 13832 21944 13860 21975
rect 15010 21972 15016 22024
rect 15068 22012 15074 22024
rect 15105 22015 15163 22021
rect 15105 22012 15117 22015
rect 15068 21984 15117 22012
rect 15068 21972 15074 21984
rect 15105 21981 15117 21984
rect 15151 21981 15163 22015
rect 15105 21975 15163 21981
rect 16022 21972 16028 22024
rect 16080 21972 16086 22024
rect 16224 22012 16252 22052
rect 16577 22049 16589 22052
rect 16623 22049 16635 22083
rect 16577 22043 16635 22049
rect 16132 21984 16252 22012
rect 13596 21916 13860 21944
rect 13924 21916 15148 21944
rect 13596 21904 13602 21916
rect 13924 21876 13952 21916
rect 13280 21848 13952 21876
rect 13097 21839 13155 21845
rect 15010 21836 15016 21888
rect 15068 21836 15074 21888
rect 15120 21876 15148 21916
rect 15654 21904 15660 21956
rect 15712 21904 15718 21956
rect 15746 21904 15752 21956
rect 15804 21944 15810 21956
rect 16132 21944 16160 21984
rect 16298 21972 16304 22024
rect 16356 21972 16362 22024
rect 16482 21972 16488 22024
rect 16540 21972 16546 22024
rect 15804 21916 16160 21944
rect 15804 21904 15810 21916
rect 16316 21876 16344 21972
rect 16390 21904 16396 21956
rect 16448 21944 16454 21956
rect 16684 21944 16712 22120
rect 16853 22117 16865 22120
rect 16899 22117 16911 22151
rect 17052 22148 17080 22188
rect 17126 22176 17132 22228
rect 17184 22176 17190 22228
rect 17954 22176 17960 22228
rect 18012 22176 18018 22228
rect 18141 22219 18199 22225
rect 18141 22185 18153 22219
rect 18187 22216 18199 22219
rect 19889 22219 19947 22225
rect 19889 22216 19901 22219
rect 18187 22188 19901 22216
rect 18187 22185 18199 22188
rect 18141 22179 18199 22185
rect 19889 22185 19901 22188
rect 19935 22185 19947 22219
rect 19889 22179 19947 22185
rect 22370 22176 22376 22228
rect 22428 22176 22434 22228
rect 22830 22216 22836 22228
rect 22480 22188 22836 22216
rect 18049 22151 18107 22157
rect 17052 22120 17172 22148
rect 16853 22111 16911 22117
rect 17144 22021 17172 22120
rect 18049 22117 18061 22151
rect 18095 22148 18107 22151
rect 18230 22148 18236 22160
rect 18095 22120 18236 22148
rect 18095 22117 18107 22120
rect 18049 22111 18107 22117
rect 18230 22108 18236 22120
rect 18288 22108 18294 22160
rect 19429 22151 19487 22157
rect 19429 22117 19441 22151
rect 19475 22148 19487 22151
rect 19794 22148 19800 22160
rect 19475 22120 19800 22148
rect 19475 22117 19487 22120
rect 19429 22111 19487 22117
rect 19794 22108 19800 22120
rect 19852 22108 19858 22160
rect 19978 22108 19984 22160
rect 20036 22108 20042 22160
rect 21269 22151 21327 22157
rect 21269 22148 21281 22151
rect 20824 22120 21281 22148
rect 17313 22083 17371 22089
rect 17313 22049 17325 22083
rect 17359 22080 17371 22083
rect 17681 22083 17739 22089
rect 17681 22080 17693 22083
rect 17359 22052 17693 22080
rect 17359 22049 17371 22052
rect 17313 22043 17371 22049
rect 17681 22049 17693 22052
rect 17727 22049 17739 22083
rect 17681 22043 17739 22049
rect 20438 22040 20444 22092
rect 20496 22040 20502 22092
rect 20824 22080 20852 22120
rect 21269 22117 21281 22120
rect 21315 22148 21327 22151
rect 22480 22148 22508 22188
rect 22830 22176 22836 22188
rect 22888 22176 22894 22228
rect 21315 22120 22508 22148
rect 22557 22151 22615 22157
rect 21315 22117 21327 22120
rect 21269 22111 21327 22117
rect 22557 22117 22569 22151
rect 22603 22117 22615 22151
rect 22557 22111 22615 22117
rect 20548 22052 20852 22080
rect 20901 22083 20959 22089
rect 17129 22015 17187 22021
rect 17129 21981 17141 22015
rect 17175 21981 17187 22015
rect 17129 21975 17187 21981
rect 17405 22015 17463 22021
rect 17405 21981 17417 22015
rect 17451 22012 17463 22015
rect 17954 22012 17960 22024
rect 17451 21984 17960 22012
rect 17451 21981 17463 21984
rect 17405 21975 17463 21981
rect 17954 21972 17960 21984
rect 18012 21972 18018 22024
rect 18233 22015 18291 22021
rect 18233 21981 18245 22015
rect 18279 21981 18291 22015
rect 18233 21975 18291 21981
rect 16448 21916 16712 21944
rect 16448 21904 16454 21916
rect 17770 21904 17776 21956
rect 17828 21944 17834 21956
rect 18248 21944 18276 21975
rect 18414 21972 18420 22024
rect 18472 21972 18478 22024
rect 20349 22015 20407 22021
rect 20349 21981 20361 22015
rect 20395 22012 20407 22015
rect 20548 22012 20576 22052
rect 20901 22049 20913 22083
rect 20947 22080 20959 22083
rect 22572 22080 22600 22111
rect 22922 22080 22928 22092
rect 20947 22052 22928 22080
rect 20947 22049 20959 22052
rect 20901 22043 20959 22049
rect 22922 22040 22928 22052
rect 22980 22040 22986 22092
rect 20395 21984 20576 22012
rect 20809 22015 20867 22021
rect 20395 21981 20407 21984
rect 20349 21975 20407 21981
rect 20809 21981 20821 22015
rect 20855 21981 20867 22015
rect 20809 21975 20867 21981
rect 22005 22015 22063 22021
rect 22005 21981 22017 22015
rect 22051 22012 22063 22015
rect 22278 22012 22284 22024
rect 22051 21984 22284 22012
rect 22051 21981 22063 21984
rect 22005 21975 22063 21981
rect 17828 21916 18276 21944
rect 19705 21947 19763 21953
rect 17828 21904 17834 21916
rect 19705 21913 19717 21947
rect 19751 21944 19763 21947
rect 20162 21944 20168 21956
rect 19751 21916 20168 21944
rect 19751 21913 19763 21916
rect 19705 21907 19763 21913
rect 20162 21904 20168 21916
rect 20220 21904 20226 21956
rect 20824 21944 20852 21975
rect 22278 21972 22284 21984
rect 22336 21972 22342 22024
rect 22830 21972 22836 22024
rect 22888 21972 22894 22024
rect 23106 21972 23112 22024
rect 23164 21972 23170 22024
rect 21545 21947 21603 21953
rect 21545 21944 21557 21947
rect 20824 21916 21557 21944
rect 15120 21848 16344 21876
rect 17037 21879 17095 21885
rect 17037 21845 17049 21879
rect 17083 21876 17095 21879
rect 17494 21876 17500 21888
rect 17083 21848 17500 21876
rect 17083 21845 17095 21848
rect 17037 21839 17095 21845
rect 17494 21836 17500 21848
rect 17552 21836 17558 21888
rect 17589 21879 17647 21885
rect 17589 21845 17601 21879
rect 17635 21876 17647 21879
rect 19058 21876 19064 21888
rect 17635 21848 19064 21876
rect 17635 21845 17647 21848
rect 17589 21839 17647 21845
rect 19058 21836 19064 21848
rect 19116 21836 19122 21888
rect 19242 21836 19248 21888
rect 19300 21836 19306 21888
rect 19426 21836 19432 21888
rect 19484 21876 19490 21888
rect 19886 21876 19892 21888
rect 19484 21848 19892 21876
rect 19484 21836 19490 21848
rect 19886 21836 19892 21848
rect 19944 21836 19950 21888
rect 19978 21836 19984 21888
rect 20036 21876 20042 21888
rect 20824 21876 20852 21916
rect 21545 21913 21557 21916
rect 21591 21913 21603 21947
rect 21545 21907 21603 21913
rect 22462 21904 22468 21956
rect 22520 21944 22526 21956
rect 23198 21944 23204 21956
rect 22520 21916 23204 21944
rect 22520 21904 22526 21916
rect 23198 21904 23204 21916
rect 23256 21904 23262 21956
rect 20036 21848 20852 21876
rect 20036 21836 20042 21848
rect 20990 21836 20996 21888
rect 21048 21876 21054 21888
rect 21085 21879 21143 21885
rect 21085 21876 21097 21879
rect 21048 21848 21097 21876
rect 21048 21836 21054 21848
rect 21085 21845 21097 21848
rect 21131 21845 21143 21879
rect 21085 21839 21143 21845
rect 22373 21879 22431 21885
rect 22373 21845 22385 21879
rect 22419 21876 22431 21879
rect 22649 21879 22707 21885
rect 22649 21876 22661 21879
rect 22419 21848 22661 21876
rect 22419 21845 22431 21848
rect 22373 21839 22431 21845
rect 22649 21845 22661 21848
rect 22695 21845 22707 21879
rect 22649 21839 22707 21845
rect 23014 21836 23020 21888
rect 23072 21836 23078 21888
rect 1104 21786 25208 21808
rect 1104 21734 4874 21786
rect 4926 21734 4938 21786
rect 4990 21734 5002 21786
rect 5054 21734 5066 21786
rect 5118 21734 5130 21786
rect 5182 21734 25208 21786
rect 1104 21712 25208 21734
rect 4801 21675 4859 21681
rect 4801 21641 4813 21675
rect 4847 21672 4859 21675
rect 4982 21672 4988 21684
rect 4847 21644 4988 21672
rect 4847 21641 4859 21644
rect 4801 21635 4859 21641
rect 4982 21632 4988 21644
rect 5040 21672 5046 21684
rect 8297 21675 8355 21681
rect 5040 21644 6500 21672
rect 5040 21632 5046 21644
rect 4154 21564 4160 21616
rect 4212 21604 4218 21616
rect 4341 21607 4399 21613
rect 4341 21604 4353 21607
rect 4212 21576 4353 21604
rect 4212 21564 4218 21576
rect 4341 21573 4353 21576
rect 4387 21573 4399 21607
rect 4341 21567 4399 21573
rect 5077 21607 5135 21613
rect 5077 21573 5089 21607
rect 5123 21604 5135 21607
rect 5445 21607 5503 21613
rect 5445 21604 5457 21607
rect 5123 21576 5457 21604
rect 5123 21573 5135 21576
rect 5077 21567 5135 21573
rect 5445 21573 5457 21576
rect 5491 21604 5503 21607
rect 6086 21604 6092 21616
rect 5491 21576 6092 21604
rect 5491 21573 5503 21576
rect 5445 21567 5503 21573
rect 6086 21564 6092 21576
rect 6144 21564 6150 21616
rect 6472 21604 6500 21644
rect 8297 21641 8309 21675
rect 8343 21672 8355 21675
rect 9398 21672 9404 21684
rect 8343 21644 9404 21672
rect 8343 21641 8355 21644
rect 8297 21635 8355 21641
rect 9398 21632 9404 21644
rect 9456 21632 9462 21684
rect 12066 21672 12072 21684
rect 10336 21644 12072 21672
rect 8757 21607 8815 21613
rect 6472 21576 8432 21604
rect 4614 21496 4620 21548
rect 4672 21536 4678 21548
rect 4893 21539 4951 21545
rect 4893 21536 4905 21539
rect 4672 21508 4905 21536
rect 4672 21496 4678 21508
rect 4893 21505 4905 21508
rect 4939 21505 4951 21539
rect 4893 21499 4951 21505
rect 5626 21496 5632 21548
rect 5684 21496 5690 21548
rect 5994 21496 6000 21548
rect 6052 21496 6058 21548
rect 6181 21539 6239 21545
rect 6181 21505 6193 21539
rect 6227 21536 6239 21539
rect 6472 21536 6500 21576
rect 8404 21548 8432 21576
rect 8757 21573 8769 21607
rect 8803 21604 8815 21607
rect 10336 21604 10364 21644
rect 12066 21632 12072 21644
rect 12124 21632 12130 21684
rect 12250 21632 12256 21684
rect 12308 21632 12314 21684
rect 12345 21675 12403 21681
rect 12345 21641 12357 21675
rect 12391 21672 12403 21675
rect 12434 21672 12440 21684
rect 12391 21644 12440 21672
rect 12391 21641 12403 21644
rect 12345 21635 12403 21641
rect 12434 21632 12440 21644
rect 12492 21632 12498 21684
rect 12529 21675 12587 21681
rect 12529 21641 12541 21675
rect 12575 21672 12587 21675
rect 12618 21672 12624 21684
rect 12575 21644 12624 21672
rect 12575 21641 12587 21644
rect 12529 21635 12587 21641
rect 12618 21632 12624 21644
rect 12676 21632 12682 21684
rect 12986 21632 12992 21684
rect 13044 21672 13050 21684
rect 15565 21675 15623 21681
rect 13044 21644 13124 21672
rect 13044 21632 13050 21644
rect 8803 21576 10364 21604
rect 8803 21573 8815 21576
rect 8757 21567 8815 21573
rect 11882 21564 11888 21616
rect 11940 21604 11946 21616
rect 13096 21604 13124 21644
rect 15565 21641 15577 21675
rect 15611 21672 15623 21675
rect 16022 21672 16028 21684
rect 15611 21644 16028 21672
rect 15611 21641 15623 21644
rect 15565 21635 15623 21641
rect 16022 21632 16028 21644
rect 16080 21632 16086 21684
rect 17954 21632 17960 21684
rect 18012 21632 18018 21684
rect 18414 21672 18420 21684
rect 18156 21644 18420 21672
rect 11940 21576 13032 21604
rect 13096 21576 15056 21604
rect 11940 21564 11946 21576
rect 6227 21508 6500 21536
rect 6227 21505 6239 21508
rect 6181 21499 6239 21505
rect 6914 21496 6920 21548
rect 6972 21496 6978 21548
rect 7650 21496 7656 21548
rect 7708 21536 7714 21548
rect 7929 21539 7987 21545
rect 7929 21536 7941 21539
rect 7708 21508 7941 21536
rect 7708 21496 7714 21508
rect 7929 21505 7941 21508
rect 7975 21536 7987 21539
rect 7975 21508 8340 21536
rect 7975 21505 7987 21508
rect 7929 21499 7987 21505
rect 5810 21468 5816 21480
rect 5644 21440 5816 21468
rect 4341 21403 4399 21409
rect 4341 21369 4353 21403
rect 4387 21400 4399 21403
rect 4706 21400 4712 21412
rect 4387 21372 4712 21400
rect 4387 21369 4399 21372
rect 4341 21363 4399 21369
rect 4706 21360 4712 21372
rect 4764 21360 4770 21412
rect 2958 21292 2964 21344
rect 3016 21332 3022 21344
rect 5644 21332 5672 21440
rect 5810 21428 5816 21440
rect 5868 21428 5874 21480
rect 5905 21471 5963 21477
rect 5905 21437 5917 21471
rect 5951 21468 5963 21471
rect 6454 21468 6460 21480
rect 5951 21440 6460 21468
rect 5951 21437 5963 21440
rect 5905 21431 5963 21437
rect 6454 21428 6460 21440
rect 6512 21468 6518 21480
rect 6825 21471 6883 21477
rect 6825 21468 6837 21471
rect 6512 21440 6837 21468
rect 6512 21428 6518 21440
rect 6825 21437 6837 21440
rect 6871 21437 6883 21471
rect 6825 21431 6883 21437
rect 8018 21428 8024 21480
rect 8076 21428 8082 21480
rect 8312 21468 8340 21508
rect 8386 21496 8392 21548
rect 8444 21496 8450 21548
rect 8570 21545 8576 21548
rect 8543 21539 8576 21545
rect 8543 21505 8555 21539
rect 8628 21536 8634 21548
rect 10778 21536 10784 21548
rect 8628 21508 10784 21536
rect 8543 21499 8576 21505
rect 8570 21496 8576 21499
rect 8628 21496 8634 21508
rect 10778 21496 10784 21508
rect 10836 21496 10842 21548
rect 11514 21496 11520 21548
rect 11572 21496 11578 21548
rect 11698 21496 11704 21548
rect 11756 21496 11762 21548
rect 11793 21539 11851 21545
rect 11793 21505 11805 21539
rect 11839 21536 11851 21539
rect 12069 21539 12127 21545
rect 11839 21508 12020 21536
rect 11839 21505 11851 21508
rect 11793 21499 11851 21505
rect 9766 21468 9772 21480
rect 8312 21440 9772 21468
rect 9766 21428 9772 21440
rect 9824 21428 9830 21480
rect 11885 21471 11943 21477
rect 11885 21468 11897 21471
rect 9968 21440 11897 21468
rect 5721 21403 5779 21409
rect 5721 21369 5733 21403
rect 5767 21400 5779 21403
rect 5997 21403 6055 21409
rect 5997 21400 6009 21403
rect 5767 21372 6009 21400
rect 5767 21369 5779 21372
rect 5721 21363 5779 21369
rect 5997 21369 6009 21372
rect 6043 21369 6055 21403
rect 5997 21363 6055 21369
rect 6546 21360 6552 21412
rect 6604 21400 6610 21412
rect 9858 21400 9864 21412
rect 6604 21372 9864 21400
rect 6604 21360 6610 21372
rect 9858 21360 9864 21372
rect 9916 21360 9922 21412
rect 3016 21304 5672 21332
rect 3016 21292 3022 21304
rect 7282 21292 7288 21344
rect 7340 21292 7346 21344
rect 8754 21292 8760 21344
rect 8812 21332 8818 21344
rect 9968 21332 9996 21440
rect 11885 21437 11897 21440
rect 11931 21437 11943 21471
rect 11992 21468 12020 21508
rect 12069 21505 12081 21539
rect 12115 21536 12127 21539
rect 12158 21536 12164 21548
rect 12115 21508 12164 21536
rect 12115 21505 12127 21508
rect 12069 21499 12127 21505
rect 12158 21496 12164 21508
rect 12216 21496 12222 21548
rect 12526 21536 12532 21548
rect 12487 21508 12532 21536
rect 12526 21496 12532 21508
rect 12584 21496 12590 21548
rect 13004 21545 13032 21576
rect 15028 21548 15056 21576
rect 15654 21564 15660 21616
rect 15712 21604 15718 21616
rect 18046 21604 18052 21616
rect 15712 21576 18052 21604
rect 15712 21564 15718 21576
rect 18046 21564 18052 21576
rect 18104 21604 18110 21616
rect 18156 21604 18184 21644
rect 18414 21632 18420 21644
rect 18472 21632 18478 21684
rect 18506 21632 18512 21684
rect 18564 21672 18570 21684
rect 18601 21675 18659 21681
rect 18601 21672 18613 21675
rect 18564 21644 18613 21672
rect 18564 21632 18570 21644
rect 18601 21641 18613 21644
rect 18647 21641 18659 21675
rect 18601 21635 18659 21641
rect 22005 21675 22063 21681
rect 22005 21641 22017 21675
rect 22051 21672 22063 21675
rect 22186 21672 22192 21684
rect 22051 21644 22192 21672
rect 22051 21641 22063 21644
rect 22005 21635 22063 21641
rect 22186 21632 22192 21644
rect 22244 21632 22250 21684
rect 22830 21632 22836 21684
rect 22888 21672 22894 21684
rect 24397 21675 24455 21681
rect 24397 21672 24409 21675
rect 22888 21644 24409 21672
rect 22888 21632 22894 21644
rect 24397 21641 24409 21644
rect 24443 21641 24455 21675
rect 24397 21635 24455 21641
rect 19242 21604 19248 21616
rect 18104 21576 18184 21604
rect 18248 21576 19248 21604
rect 18104 21564 18110 21576
rect 12989 21539 13047 21545
rect 12989 21505 13001 21539
rect 13035 21536 13047 21539
rect 13262 21536 13268 21548
rect 13035 21508 13268 21536
rect 13035 21505 13047 21508
rect 12989 21499 13047 21505
rect 13262 21496 13268 21508
rect 13320 21496 13326 21548
rect 13354 21496 13360 21548
rect 13412 21496 13418 21548
rect 13446 21496 13452 21548
rect 13504 21496 13510 21548
rect 13630 21496 13636 21548
rect 13688 21496 13694 21548
rect 13722 21496 13728 21548
rect 13780 21496 13786 21548
rect 15010 21496 15016 21548
rect 15068 21536 15074 21548
rect 15068 21508 15240 21536
rect 15068 21496 15074 21508
rect 12894 21468 12900 21480
rect 11992 21440 12900 21468
rect 11885 21431 11943 21437
rect 12894 21428 12900 21440
rect 12952 21428 12958 21480
rect 15102 21428 15108 21480
rect 15160 21428 15166 21480
rect 15212 21468 15240 21508
rect 15470 21496 15476 21548
rect 15528 21536 15534 21548
rect 16117 21539 16175 21545
rect 16117 21536 16129 21539
rect 15528 21508 16129 21536
rect 15528 21496 15534 21508
rect 16117 21505 16129 21508
rect 16163 21536 16175 21539
rect 16298 21536 16304 21548
rect 16163 21508 16304 21536
rect 16163 21505 16175 21508
rect 16117 21499 16175 21505
rect 16298 21496 16304 21508
rect 16356 21496 16362 21548
rect 16666 21496 16672 21548
rect 16724 21496 16730 21548
rect 16758 21496 16764 21548
rect 16816 21496 16822 21548
rect 16942 21496 16948 21548
rect 17000 21496 17006 21548
rect 17034 21496 17040 21548
rect 17092 21496 17098 21548
rect 17126 21496 17132 21548
rect 17184 21496 17190 21548
rect 17770 21536 17776 21548
rect 17236 21508 17776 21536
rect 17236 21468 17264 21508
rect 17770 21496 17776 21508
rect 17828 21496 17834 21548
rect 18248 21545 18276 21576
rect 19242 21564 19248 21576
rect 19300 21564 19306 21616
rect 22922 21564 22928 21616
rect 22980 21564 22986 21616
rect 23198 21564 23204 21616
rect 23256 21604 23262 21616
rect 23256 21576 23414 21604
rect 23256 21564 23262 21576
rect 18233 21539 18291 21545
rect 18233 21505 18245 21539
rect 18279 21505 18291 21539
rect 18233 21499 18291 21505
rect 18322 21496 18328 21548
rect 18380 21496 18386 21548
rect 18693 21539 18751 21545
rect 18693 21505 18705 21539
rect 18739 21536 18751 21539
rect 18874 21536 18880 21548
rect 18739 21508 18880 21536
rect 18739 21505 18751 21508
rect 18693 21499 18751 21505
rect 18874 21496 18880 21508
rect 18932 21496 18938 21548
rect 20349 21539 20407 21545
rect 20349 21536 20361 21539
rect 18984 21508 20361 21536
rect 15212 21440 17264 21468
rect 17494 21428 17500 21480
rect 17552 21468 17558 21480
rect 18417 21471 18475 21477
rect 18417 21468 18429 21471
rect 17552 21440 18429 21468
rect 17552 21428 17558 21440
rect 18417 21437 18429 21440
rect 18463 21437 18475 21471
rect 18417 21431 18475 21437
rect 10042 21360 10048 21412
rect 10100 21400 10106 21412
rect 11974 21400 11980 21412
rect 10100 21372 11980 21400
rect 10100 21360 10106 21372
rect 11974 21360 11980 21372
rect 12032 21360 12038 21412
rect 15473 21403 15531 21409
rect 12912 21372 13308 21400
rect 8812 21304 9996 21332
rect 8812 21292 8818 21304
rect 10594 21292 10600 21344
rect 10652 21332 10658 21344
rect 12912 21341 12940 21372
rect 12897 21335 12955 21341
rect 12897 21332 12909 21335
rect 10652 21304 12909 21332
rect 10652 21292 10658 21304
rect 12897 21301 12909 21304
rect 12943 21301 12955 21335
rect 12897 21295 12955 21301
rect 12986 21292 12992 21344
rect 13044 21332 13050 21344
rect 13173 21335 13231 21341
rect 13173 21332 13185 21335
rect 13044 21304 13185 21332
rect 13044 21292 13050 21304
rect 13173 21301 13185 21304
rect 13219 21301 13231 21335
rect 13280 21332 13308 21372
rect 15473 21369 15485 21403
rect 15519 21400 15531 21403
rect 15562 21400 15568 21412
rect 15519 21372 15568 21400
rect 15519 21369 15531 21372
rect 15473 21363 15531 21369
rect 15562 21360 15568 21372
rect 15620 21360 15626 21412
rect 17405 21403 17463 21409
rect 17405 21369 17417 21403
rect 17451 21400 17463 21403
rect 18984 21400 19012 21508
rect 20349 21505 20361 21508
rect 20395 21505 20407 21539
rect 20349 21499 20407 21505
rect 20714 21496 20720 21548
rect 20772 21536 20778 21548
rect 20993 21539 21051 21545
rect 20993 21536 21005 21539
rect 20772 21508 21005 21536
rect 20772 21496 20778 21508
rect 20993 21505 21005 21508
rect 21039 21536 21051 21539
rect 21542 21536 21548 21548
rect 21039 21508 21548 21536
rect 21039 21505 21051 21508
rect 20993 21499 21051 21505
rect 21542 21496 21548 21508
rect 21600 21496 21606 21548
rect 21637 21539 21695 21545
rect 21637 21505 21649 21539
rect 21683 21536 21695 21539
rect 21683 21508 22032 21536
rect 21683 21505 21695 21508
rect 21637 21499 21695 21505
rect 19886 21468 19892 21480
rect 17451 21372 19012 21400
rect 19168 21440 19892 21468
rect 17451 21369 17463 21372
rect 17405 21363 17463 21369
rect 19168 21332 19196 21440
rect 19886 21428 19892 21440
rect 19944 21428 19950 21480
rect 20070 21428 20076 21480
rect 20128 21428 20134 21480
rect 20916 21440 21404 21468
rect 13280 21304 19196 21332
rect 13173 21295 13231 21301
rect 19242 21292 19248 21344
rect 19300 21332 19306 21344
rect 19797 21335 19855 21341
rect 19797 21332 19809 21335
rect 19300 21304 19809 21332
rect 19300 21292 19306 21304
rect 19797 21301 19809 21304
rect 19843 21301 19855 21335
rect 19797 21295 19855 21301
rect 20257 21335 20315 21341
rect 20257 21301 20269 21335
rect 20303 21332 20315 21335
rect 20916 21332 20944 21440
rect 21269 21403 21327 21409
rect 21269 21369 21281 21403
rect 21315 21369 21327 21403
rect 21376 21400 21404 21440
rect 21910 21428 21916 21480
rect 21968 21428 21974 21480
rect 22004 21468 22032 21508
rect 22094 21496 22100 21548
rect 22152 21496 22158 21548
rect 22370 21496 22376 21548
rect 22428 21496 22434 21548
rect 22004 21440 22600 21468
rect 21821 21403 21879 21409
rect 21821 21400 21833 21403
rect 21376 21372 21833 21400
rect 21269 21363 21327 21369
rect 21821 21369 21833 21372
rect 21867 21369 21879 21403
rect 22462 21400 22468 21412
rect 21821 21363 21879 21369
rect 21928 21372 22468 21400
rect 20303 21304 20944 21332
rect 20303 21301 20315 21304
rect 20257 21295 20315 21301
rect 21174 21292 21180 21344
rect 21232 21292 21238 21344
rect 21284 21332 21312 21363
rect 21726 21332 21732 21344
rect 21284 21304 21732 21332
rect 21726 21292 21732 21304
rect 21784 21332 21790 21344
rect 21928 21332 21956 21372
rect 22462 21360 22468 21372
rect 22520 21360 22526 21412
rect 21784 21304 21956 21332
rect 21784 21292 21790 21304
rect 22094 21292 22100 21344
rect 22152 21332 22158 21344
rect 22281 21335 22339 21341
rect 22281 21332 22293 21335
rect 22152 21304 22293 21332
rect 22152 21292 22158 21304
rect 22281 21301 22293 21304
rect 22327 21301 22339 21335
rect 22572 21332 22600 21440
rect 22646 21428 22652 21480
rect 22704 21428 22710 21480
rect 23014 21332 23020 21344
rect 22572 21304 23020 21332
rect 22281 21295 22339 21301
rect 23014 21292 23020 21304
rect 23072 21292 23078 21344
rect 1104 21242 25208 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 25208 21242
rect 1104 21168 25208 21190
rect 4982 21088 4988 21140
rect 5040 21088 5046 21140
rect 8294 21088 8300 21140
rect 8352 21088 8358 21140
rect 9674 21088 9680 21140
rect 9732 21128 9738 21140
rect 10137 21131 10195 21137
rect 10137 21128 10149 21131
rect 9732 21100 10149 21128
rect 9732 21088 9738 21100
rect 10137 21097 10149 21100
rect 10183 21097 10195 21131
rect 10137 21091 10195 21097
rect 10410 21088 10416 21140
rect 10468 21128 10474 21140
rect 10781 21131 10839 21137
rect 10781 21128 10793 21131
rect 10468 21100 10793 21128
rect 10468 21088 10474 21100
rect 10781 21097 10793 21100
rect 10827 21097 10839 21131
rect 10781 21091 10839 21097
rect 10965 21131 11023 21137
rect 10965 21097 10977 21131
rect 11011 21097 11023 21131
rect 10965 21091 11023 21097
rect 13541 21131 13599 21137
rect 13541 21097 13553 21131
rect 13587 21128 13599 21131
rect 13722 21128 13728 21140
rect 13587 21100 13728 21128
rect 13587 21097 13599 21100
rect 13541 21091 13599 21097
rect 2774 21020 2780 21072
rect 2832 21060 2838 21072
rect 4522 21060 4528 21072
rect 2832 21032 4528 21060
rect 2832 21020 2838 21032
rect 4522 21020 4528 21032
rect 4580 21020 4586 21072
rect 7282 21020 7288 21072
rect 7340 21060 7346 21072
rect 9953 21063 10011 21069
rect 7340 21032 8432 21060
rect 7340 21020 7346 21032
rect 1394 20952 1400 21004
rect 1452 20952 1458 21004
rect 2792 20910 2820 21020
rect 3145 20995 3203 21001
rect 3145 20961 3157 20995
rect 3191 20992 3203 20995
rect 4706 20992 4712 21004
rect 3191 20964 4712 20992
rect 3191 20961 3203 20964
rect 3145 20955 3203 20961
rect 3050 20884 3056 20936
rect 3108 20924 3114 20936
rect 3467 20927 3525 20933
rect 3467 20924 3479 20927
rect 3108 20896 3479 20924
rect 3108 20884 3114 20896
rect 3466 20893 3479 20896
rect 3513 20893 3525 20927
rect 3466 20887 3525 20893
rect 1670 20816 1676 20868
rect 1728 20816 1734 20868
rect 3466 20856 3494 20887
rect 3602 20884 3608 20936
rect 3660 20884 3666 20936
rect 3804 20933 3832 20964
rect 4706 20952 4712 20964
rect 4764 20952 4770 21004
rect 6362 20952 6368 21004
rect 6420 20992 6426 21004
rect 6733 20995 6791 21001
rect 6733 20992 6745 20995
rect 6420 20964 6745 20992
rect 6420 20952 6426 20964
rect 6733 20961 6745 20964
rect 6779 20992 6791 20995
rect 8110 20992 8116 21004
rect 6779 20964 8116 20992
rect 6779 20961 6791 20964
rect 6733 20955 6791 20961
rect 8110 20952 8116 20964
rect 8168 20952 8174 21004
rect 8404 21001 8432 21032
rect 9953 21029 9965 21063
rect 9999 21060 10011 21063
rect 10980 21060 11008 21091
rect 13722 21088 13728 21100
rect 13780 21088 13786 21140
rect 18230 21088 18236 21140
rect 18288 21088 18294 21140
rect 21634 21088 21640 21140
rect 21692 21128 21698 21140
rect 22646 21128 22652 21140
rect 21692 21100 22652 21128
rect 21692 21088 21698 21100
rect 22646 21088 22652 21100
rect 22704 21088 22710 21140
rect 9999 21032 11008 21060
rect 15565 21063 15623 21069
rect 9999 21029 10011 21032
rect 9953 21023 10011 21029
rect 15565 21029 15577 21063
rect 15611 21060 15623 21063
rect 16942 21060 16948 21072
rect 15611 21032 16948 21060
rect 15611 21029 15623 21032
rect 15565 21023 15623 21029
rect 16942 21020 16948 21032
rect 17000 21020 17006 21072
rect 17954 21020 17960 21072
rect 18012 21060 18018 21072
rect 18049 21063 18107 21069
rect 18049 21060 18061 21063
rect 18012 21032 18061 21060
rect 18012 21020 18018 21032
rect 18049 21029 18061 21032
rect 18095 21029 18107 21063
rect 18049 21023 18107 21029
rect 20349 21063 20407 21069
rect 20349 21029 20361 21063
rect 20395 21060 20407 21063
rect 21910 21060 21916 21072
rect 20395 21032 21916 21060
rect 20395 21029 20407 21032
rect 20349 21023 20407 21029
rect 21910 21020 21916 21032
rect 21968 21020 21974 21072
rect 23106 21020 23112 21072
rect 23164 21060 23170 21072
rect 23474 21060 23480 21072
rect 23164 21032 23480 21060
rect 23164 21020 23170 21032
rect 23474 21020 23480 21032
rect 23532 21020 23538 21072
rect 8389 20995 8447 21001
rect 8389 20961 8401 20995
rect 8435 20961 8447 20995
rect 8389 20955 8447 20961
rect 9677 20995 9735 21001
rect 9677 20961 9689 20995
rect 9723 20992 9735 20995
rect 9858 20992 9864 21004
rect 9723 20964 9864 20992
rect 9723 20961 9735 20964
rect 9677 20955 9735 20961
rect 9858 20952 9864 20964
rect 9916 20952 9922 21004
rect 10226 20952 10232 21004
rect 10284 20992 10290 21004
rect 10321 20995 10379 21001
rect 10321 20992 10333 20995
rect 10284 20964 10333 20992
rect 10284 20952 10290 20964
rect 10321 20961 10333 20964
rect 10367 20961 10379 20995
rect 11057 20995 11115 21001
rect 11057 20992 11069 20995
rect 10321 20955 10379 20961
rect 10428 20964 11069 20992
rect 3789 20927 3847 20933
rect 3789 20893 3801 20927
rect 3835 20893 3847 20927
rect 3789 20887 3847 20893
rect 4154 20884 4160 20936
rect 4212 20884 4218 20936
rect 4614 20884 4620 20936
rect 4672 20884 4678 20936
rect 8570 20884 8576 20936
rect 8628 20884 8634 20936
rect 9582 20884 9588 20936
rect 9640 20884 9646 20936
rect 4062 20856 4068 20868
rect 3466 20828 4068 20856
rect 4062 20816 4068 20828
rect 4120 20816 4126 20868
rect 6178 20856 6184 20868
rect 6026 20828 6184 20856
rect 3234 20748 3240 20800
rect 3292 20748 3298 20800
rect 3602 20748 3608 20800
rect 3660 20788 3666 20800
rect 3881 20791 3939 20797
rect 3881 20788 3893 20791
rect 3660 20760 3893 20788
rect 3660 20748 3666 20760
rect 3881 20757 3893 20760
rect 3927 20757 3939 20791
rect 3881 20751 3939 20757
rect 4522 20748 4528 20800
rect 4580 20788 4586 20800
rect 4798 20788 4804 20800
rect 4580 20760 4804 20788
rect 4580 20748 4586 20760
rect 4798 20748 4804 20760
rect 4856 20788 4862 20800
rect 6104 20788 6132 20828
rect 6178 20816 6184 20828
rect 6236 20816 6242 20868
rect 6454 20816 6460 20868
rect 6512 20816 6518 20868
rect 8294 20816 8300 20868
rect 8352 20816 8358 20868
rect 10042 20816 10048 20868
rect 10100 20816 10106 20868
rect 4856 20760 6132 20788
rect 8757 20791 8815 20797
rect 4856 20748 4862 20760
rect 8757 20757 8769 20791
rect 8803 20788 8815 20791
rect 10428 20788 10456 20964
rect 11057 20961 11069 20964
rect 11103 20961 11115 20995
rect 11057 20955 11115 20961
rect 13354 20952 13360 21004
rect 13412 20952 13418 21004
rect 16390 20992 16396 21004
rect 15212 20964 16396 20992
rect 10502 20884 10508 20936
rect 10560 20884 10566 20936
rect 10965 20927 11023 20933
rect 10965 20924 10977 20927
rect 10704 20896 10977 20924
rect 10704 20797 10732 20896
rect 10965 20893 10977 20896
rect 11011 20893 11023 20927
rect 10965 20887 11023 20893
rect 11241 20927 11299 20933
rect 11241 20893 11253 20927
rect 11287 20924 11299 20927
rect 12986 20924 12992 20936
rect 11287 20896 12992 20924
rect 11287 20893 11299 20896
rect 11241 20887 11299 20893
rect 12986 20884 12992 20896
rect 13044 20884 13050 20936
rect 13265 20927 13323 20933
rect 13265 20893 13277 20927
rect 13311 20924 13323 20927
rect 13814 20924 13820 20936
rect 13311 20896 13820 20924
rect 13311 20893 13323 20896
rect 13265 20887 13323 20893
rect 13814 20884 13820 20896
rect 13872 20884 13878 20936
rect 15212 20933 15240 20964
rect 16390 20952 16396 20964
rect 16448 20952 16454 21004
rect 19058 20952 19064 21004
rect 19116 20992 19122 21004
rect 19116 20964 19472 20992
rect 19116 20952 19122 20964
rect 15197 20927 15255 20933
rect 15197 20893 15209 20927
rect 15243 20893 15255 20927
rect 15197 20887 15255 20893
rect 15351 20927 15409 20933
rect 15351 20893 15363 20927
rect 15397 20924 15409 20927
rect 15746 20924 15752 20936
rect 15397 20896 15752 20924
rect 15397 20893 15409 20896
rect 15351 20887 15409 20893
rect 15746 20884 15752 20896
rect 15804 20924 15810 20936
rect 16022 20924 16028 20936
rect 15804 20896 16028 20924
rect 15804 20884 15810 20896
rect 16022 20884 16028 20896
rect 16080 20884 16086 20936
rect 16758 20884 16764 20936
rect 16816 20924 16822 20936
rect 17405 20927 17463 20933
rect 17405 20924 17417 20927
rect 16816 20896 17417 20924
rect 16816 20884 16822 20896
rect 17405 20893 17417 20896
rect 17451 20924 17463 20927
rect 17451 20896 19196 20924
rect 17451 20893 17463 20896
rect 17405 20887 17463 20893
rect 10778 20816 10784 20868
rect 10836 20856 10842 20868
rect 13906 20856 13912 20868
rect 10836 20828 13912 20856
rect 10836 20816 10842 20828
rect 13906 20816 13912 20828
rect 13964 20856 13970 20868
rect 15838 20856 15844 20868
rect 13964 20828 15844 20856
rect 13964 20816 13970 20828
rect 15838 20816 15844 20828
rect 15896 20816 15902 20868
rect 17494 20816 17500 20868
rect 17552 20856 17558 20868
rect 17773 20859 17831 20865
rect 17773 20856 17785 20859
rect 17552 20828 17785 20856
rect 17552 20816 17558 20828
rect 17773 20825 17785 20828
rect 17819 20856 17831 20859
rect 17862 20856 17868 20868
rect 17819 20828 17868 20856
rect 17819 20825 17831 20828
rect 17773 20819 17831 20825
rect 17862 20816 17868 20828
rect 17920 20816 17926 20868
rect 18877 20859 18935 20865
rect 18877 20825 18889 20859
rect 18923 20825 18935 20859
rect 18877 20819 18935 20825
rect 8803 20760 10456 20788
rect 10689 20791 10747 20797
rect 8803 20757 8815 20760
rect 8757 20751 8815 20757
rect 10689 20757 10701 20791
rect 10735 20757 10747 20791
rect 10689 20751 10747 20757
rect 16117 20791 16175 20797
rect 16117 20757 16129 20791
rect 16163 20788 16175 20791
rect 16298 20788 16304 20800
rect 16163 20760 16304 20788
rect 16163 20757 16175 20760
rect 16117 20751 16175 20757
rect 16298 20748 16304 20760
rect 16356 20748 16362 20800
rect 18690 20748 18696 20800
rect 18748 20748 18754 20800
rect 18892 20788 18920 20819
rect 19058 20816 19064 20868
rect 19116 20816 19122 20868
rect 19168 20856 19196 20896
rect 19242 20884 19248 20936
rect 19300 20884 19306 20936
rect 19444 20933 19472 20964
rect 22370 20952 22376 21004
rect 22428 20992 22434 21004
rect 23124 20992 23152 21020
rect 23569 20995 23627 21001
rect 23569 20992 23581 20995
rect 22428 20964 23152 20992
rect 22428 20952 22434 20964
rect 19429 20927 19487 20933
rect 19429 20893 19441 20927
rect 19475 20893 19487 20927
rect 19429 20887 19487 20893
rect 19702 20884 19708 20936
rect 19760 20884 19766 20936
rect 19794 20884 19800 20936
rect 19852 20924 19858 20936
rect 20162 20933 20168 20936
rect 19981 20927 20039 20933
rect 19981 20924 19993 20927
rect 19852 20896 19993 20924
rect 19852 20884 19858 20896
rect 19981 20893 19993 20896
rect 20027 20893 20039 20927
rect 19981 20887 20039 20893
rect 20135 20927 20168 20933
rect 20135 20893 20147 20927
rect 20135 20887 20168 20893
rect 20162 20884 20168 20887
rect 20220 20884 20226 20936
rect 23014 20884 23020 20936
rect 23072 20884 23078 20936
rect 23124 20933 23152 20964
rect 23216 20964 23581 20992
rect 23216 20933 23244 20964
rect 23569 20961 23581 20964
rect 23615 20961 23627 20995
rect 23569 20955 23627 20961
rect 23109 20927 23167 20933
rect 23109 20893 23121 20927
rect 23155 20893 23167 20927
rect 23109 20887 23167 20893
rect 23201 20927 23259 20933
rect 23201 20893 23213 20927
rect 23247 20893 23259 20927
rect 23201 20887 23259 20893
rect 23382 20884 23388 20936
rect 23440 20884 23446 20936
rect 23474 20884 23480 20936
rect 23532 20884 23538 20936
rect 23658 20884 23664 20936
rect 23716 20884 23722 20936
rect 20533 20859 20591 20865
rect 20533 20856 20545 20859
rect 19168 20828 20545 20856
rect 20533 20825 20545 20828
rect 20579 20825 20591 20859
rect 23032 20856 23060 20884
rect 23676 20856 23704 20884
rect 23032 20828 23704 20856
rect 20533 20819 20591 20825
rect 19242 20788 19248 20800
rect 18892 20760 19248 20788
rect 19242 20748 19248 20760
rect 19300 20748 19306 20800
rect 19426 20748 19432 20800
rect 19484 20788 19490 20800
rect 19889 20791 19947 20797
rect 19889 20788 19901 20791
rect 19484 20760 19901 20788
rect 19484 20748 19490 20760
rect 19889 20757 19901 20760
rect 19935 20757 19947 20791
rect 19889 20751 19947 20757
rect 21634 20748 21640 20800
rect 21692 20788 21698 20800
rect 21821 20791 21879 20797
rect 21821 20788 21833 20791
rect 21692 20760 21833 20788
rect 21692 20748 21698 20760
rect 21821 20757 21833 20760
rect 21867 20757 21879 20791
rect 21821 20751 21879 20757
rect 22738 20748 22744 20800
rect 22796 20748 22802 20800
rect 1104 20698 25208 20720
rect 1104 20646 4874 20698
rect 4926 20646 4938 20698
rect 4990 20646 5002 20698
rect 5054 20646 5066 20698
rect 5118 20646 5130 20698
rect 5182 20646 25208 20698
rect 1104 20624 25208 20646
rect 1670 20544 1676 20596
rect 1728 20584 1734 20596
rect 2317 20587 2375 20593
rect 2317 20584 2329 20587
rect 1728 20556 2329 20584
rect 1728 20544 1734 20556
rect 2317 20553 2329 20556
rect 2363 20553 2375 20587
rect 3602 20584 3608 20596
rect 2317 20547 2375 20553
rect 2516 20556 3608 20584
rect 2516 20457 2544 20556
rect 3602 20544 3608 20556
rect 3660 20544 3666 20596
rect 4062 20544 4068 20596
rect 4120 20584 4126 20596
rect 5445 20587 5503 20593
rect 5445 20584 5457 20587
rect 4120 20556 5457 20584
rect 4120 20544 4126 20556
rect 5445 20553 5457 20556
rect 5491 20553 5503 20587
rect 9861 20587 9919 20593
rect 5445 20547 5503 20553
rect 7024 20556 8432 20584
rect 2958 20516 2964 20528
rect 2608 20488 2964 20516
rect 2608 20457 2636 20488
rect 2958 20476 2964 20488
rect 3016 20476 3022 20528
rect 3234 20476 3240 20528
rect 3292 20476 3298 20528
rect 4522 20516 4528 20528
rect 4462 20488 4528 20516
rect 4522 20476 4528 20488
rect 4580 20476 4586 20528
rect 4985 20519 5043 20525
rect 4985 20485 4997 20519
rect 5031 20485 5043 20519
rect 4985 20479 5043 20485
rect 2501 20451 2559 20457
rect 2501 20417 2513 20451
rect 2547 20417 2559 20451
rect 2501 20411 2559 20417
rect 2593 20451 2651 20457
rect 2593 20417 2605 20451
rect 2639 20417 2651 20451
rect 2593 20411 2651 20417
rect 2774 20408 2780 20460
rect 2832 20408 2838 20460
rect 2866 20408 2872 20460
rect 2924 20408 2930 20460
rect 4614 20408 4620 20460
rect 4672 20448 4678 20460
rect 5000 20448 5028 20479
rect 6178 20476 6184 20528
rect 6236 20516 6242 20528
rect 6733 20519 6791 20525
rect 6733 20516 6745 20519
rect 6236 20488 6745 20516
rect 6236 20476 6242 20488
rect 6733 20485 6745 20488
rect 6779 20485 6791 20519
rect 6733 20479 6791 20485
rect 5442 20448 5448 20460
rect 4672 20420 5448 20448
rect 4672 20408 4678 20420
rect 2682 20340 2688 20392
rect 2740 20380 2746 20392
rect 4724 20389 4752 20420
rect 5442 20408 5448 20420
rect 5500 20448 5506 20460
rect 7024 20457 7052 20556
rect 8404 20528 8432 20556
rect 9861 20553 9873 20587
rect 9907 20584 9919 20587
rect 10042 20584 10048 20596
rect 9907 20556 10048 20584
rect 9907 20553 9919 20556
rect 9861 20547 9919 20553
rect 10042 20544 10048 20556
rect 10100 20544 10106 20596
rect 13354 20544 13360 20596
rect 13412 20584 13418 20596
rect 13633 20587 13691 20593
rect 13633 20584 13645 20587
rect 13412 20556 13645 20584
rect 13412 20544 13418 20556
rect 13633 20553 13645 20556
rect 13679 20553 13691 20587
rect 13633 20547 13691 20553
rect 7374 20476 7380 20528
rect 7432 20516 7438 20528
rect 8202 20525 8208 20528
rect 8173 20519 8208 20525
rect 8173 20516 8185 20519
rect 7432 20488 8185 20516
rect 7432 20476 7438 20488
rect 8173 20485 8185 20488
rect 8173 20479 8208 20485
rect 8202 20476 8208 20479
rect 8260 20476 8266 20528
rect 8386 20476 8392 20528
rect 8444 20476 8450 20528
rect 8662 20476 8668 20528
rect 8720 20476 8726 20528
rect 10594 20516 10600 20528
rect 10244 20488 10600 20516
rect 5629 20451 5687 20457
rect 5629 20448 5641 20451
rect 5500 20420 5641 20448
rect 5500 20408 5506 20420
rect 5629 20417 5641 20420
rect 5675 20417 5687 20451
rect 5629 20411 5687 20417
rect 5997 20451 6055 20457
rect 5997 20417 6009 20451
rect 6043 20417 6055 20451
rect 5997 20411 6055 20417
rect 7009 20451 7067 20457
rect 7009 20417 7021 20451
rect 7055 20417 7067 20451
rect 7009 20411 7067 20417
rect 7561 20451 7619 20457
rect 7561 20417 7573 20451
rect 7607 20448 7619 20451
rect 7650 20448 7656 20460
rect 7607 20420 7656 20448
rect 7607 20417 7619 20420
rect 7561 20411 7619 20417
rect 2961 20383 3019 20389
rect 2961 20380 2973 20383
rect 2740 20352 2973 20380
rect 2740 20340 2746 20352
rect 2961 20349 2973 20352
rect 3007 20349 3019 20383
rect 2961 20343 3019 20349
rect 4709 20383 4767 20389
rect 4709 20349 4721 20383
rect 4755 20349 4767 20383
rect 6012 20380 6040 20411
rect 7650 20408 7656 20420
rect 7708 20408 7714 20460
rect 10244 20457 10272 20488
rect 10594 20476 10600 20488
rect 10652 20476 10658 20528
rect 13078 20476 13084 20528
rect 13136 20516 13142 20528
rect 13265 20519 13323 20525
rect 13265 20516 13277 20519
rect 13136 20488 13277 20516
rect 13136 20476 13142 20488
rect 13265 20485 13277 20488
rect 13311 20485 13323 20519
rect 13265 20479 13323 20485
rect 10229 20451 10287 20457
rect 10229 20417 10241 20451
rect 10275 20417 10287 20451
rect 10229 20411 10287 20417
rect 12802 20408 12808 20460
rect 12860 20408 12866 20460
rect 13446 20408 13452 20460
rect 13504 20408 13510 20460
rect 13648 20448 13676 20547
rect 15562 20544 15568 20596
rect 15620 20584 15626 20596
rect 15930 20584 15936 20596
rect 15620 20556 15936 20584
rect 15620 20544 15626 20556
rect 15930 20544 15936 20556
rect 15988 20544 15994 20596
rect 16206 20544 16212 20596
rect 16264 20584 16270 20596
rect 16669 20587 16727 20593
rect 16669 20584 16681 20587
rect 16264 20556 16681 20584
rect 16264 20544 16270 20556
rect 16669 20553 16681 20556
rect 16715 20553 16727 20587
rect 16669 20547 16727 20553
rect 17034 20544 17040 20596
rect 17092 20584 17098 20596
rect 17221 20587 17279 20593
rect 17221 20584 17233 20587
rect 17092 20556 17233 20584
rect 17092 20544 17098 20556
rect 17221 20553 17233 20556
rect 17267 20553 17279 20587
rect 19702 20584 19708 20596
rect 17221 20547 17279 20553
rect 18616 20556 19708 20584
rect 14642 20476 14648 20528
rect 14700 20516 14706 20528
rect 14700 20488 15700 20516
rect 14700 20476 14706 20488
rect 13725 20451 13783 20457
rect 13725 20448 13737 20451
rect 13648 20420 13737 20448
rect 13725 20417 13737 20420
rect 13771 20417 13783 20451
rect 13725 20411 13783 20417
rect 15562 20408 15568 20460
rect 15620 20408 15626 20460
rect 15672 20448 15700 20488
rect 15838 20476 15844 20528
rect 15896 20516 15902 20528
rect 18616 20525 18644 20556
rect 19702 20544 19708 20556
rect 19760 20544 19766 20596
rect 20070 20544 20076 20596
rect 20128 20584 20134 20596
rect 20533 20587 20591 20593
rect 20533 20584 20545 20587
rect 20128 20556 20545 20584
rect 20128 20544 20134 20556
rect 20533 20553 20545 20556
rect 20579 20553 20591 20587
rect 20533 20547 20591 20553
rect 21177 20587 21235 20593
rect 21177 20553 21189 20587
rect 21223 20584 21235 20587
rect 22002 20584 22008 20596
rect 21223 20556 22008 20584
rect 21223 20553 21235 20556
rect 21177 20547 21235 20553
rect 22002 20544 22008 20556
rect 22060 20584 22066 20596
rect 22060 20544 22094 20584
rect 23658 20544 23664 20596
rect 23716 20584 23722 20596
rect 24765 20587 24823 20593
rect 24765 20584 24777 20587
rect 23716 20556 24777 20584
rect 23716 20544 23722 20556
rect 24765 20553 24777 20556
rect 24811 20553 24823 20587
rect 24765 20547 24823 20553
rect 17129 20519 17187 20525
rect 17129 20516 17141 20519
rect 15896 20488 17141 20516
rect 15896 20476 15902 20488
rect 17129 20485 17141 20488
rect 17175 20516 17187 20519
rect 18601 20519 18659 20525
rect 17175 20488 18092 20516
rect 17175 20485 17187 20488
rect 17129 20479 17187 20485
rect 15672 20420 15792 20448
rect 4709 20343 4767 20349
rect 5276 20352 6040 20380
rect 6733 20383 6791 20389
rect 4614 20272 4620 20324
rect 4672 20312 4678 20324
rect 4672 20284 5028 20312
rect 4672 20272 4678 20284
rect 3602 20204 3608 20256
rect 3660 20244 3666 20256
rect 5000 20253 5028 20284
rect 5276 20256 5304 20352
rect 6733 20349 6745 20383
rect 6779 20349 6791 20383
rect 6733 20343 6791 20349
rect 5350 20272 5356 20324
rect 5408 20312 5414 20324
rect 5408 20284 5672 20312
rect 5408 20272 5414 20284
rect 4801 20247 4859 20253
rect 4801 20244 4813 20247
rect 3660 20216 4813 20244
rect 3660 20204 3666 20216
rect 4801 20213 4813 20216
rect 4847 20213 4859 20247
rect 4801 20207 4859 20213
rect 4985 20247 5043 20253
rect 4985 20213 4997 20247
rect 5031 20244 5043 20247
rect 5258 20244 5264 20256
rect 5031 20216 5264 20244
rect 5031 20213 5043 20216
rect 4985 20207 5043 20213
rect 5258 20204 5264 20216
rect 5316 20204 5322 20256
rect 5644 20253 5672 20284
rect 5629 20247 5687 20253
rect 5629 20213 5641 20247
rect 5675 20213 5687 20247
rect 6748 20244 6776 20343
rect 7098 20340 7104 20392
rect 7156 20380 7162 20392
rect 7469 20383 7527 20389
rect 7469 20380 7481 20383
rect 7156 20352 7481 20380
rect 7156 20340 7162 20352
rect 7469 20349 7481 20352
rect 7515 20349 7527 20383
rect 7469 20343 7527 20349
rect 7929 20383 7987 20389
rect 7929 20349 7941 20383
rect 7975 20380 7987 20383
rect 8570 20380 8576 20392
rect 7975 20352 8576 20380
rect 7975 20349 7987 20352
rect 7929 20343 7987 20349
rect 8570 20340 8576 20352
rect 8628 20340 8634 20392
rect 10321 20383 10379 20389
rect 10321 20349 10333 20383
rect 10367 20380 10379 20383
rect 10594 20380 10600 20392
rect 10367 20352 10600 20380
rect 10367 20349 10379 20352
rect 10321 20343 10379 20349
rect 10594 20340 10600 20352
rect 10652 20340 10658 20392
rect 12894 20340 12900 20392
rect 12952 20340 12958 20392
rect 13173 20383 13231 20389
rect 13173 20349 13185 20383
rect 13219 20380 13231 20383
rect 13630 20380 13636 20392
rect 13219 20352 13636 20380
rect 13219 20349 13231 20352
rect 13173 20343 13231 20349
rect 13630 20340 13636 20352
rect 13688 20340 13694 20392
rect 15654 20340 15660 20392
rect 15712 20340 15718 20392
rect 15764 20380 15792 20420
rect 15930 20408 15936 20460
rect 15988 20448 15994 20460
rect 16025 20451 16083 20457
rect 16025 20448 16037 20451
rect 15988 20420 16037 20448
rect 15988 20408 15994 20420
rect 16025 20417 16037 20420
rect 16071 20417 16083 20451
rect 17494 20448 17500 20460
rect 16025 20411 16083 20417
rect 16224 20420 17356 20448
rect 17455 20420 17500 20448
rect 16224 20380 16252 20420
rect 15764 20352 16252 20380
rect 16485 20383 16543 20389
rect 16485 20349 16497 20383
rect 16531 20380 16543 20383
rect 17328 20380 17356 20420
rect 17494 20408 17500 20420
rect 17552 20408 17558 20460
rect 17589 20451 17647 20457
rect 17589 20417 17601 20451
rect 17635 20448 17647 20451
rect 17954 20448 17960 20460
rect 17635 20420 17960 20448
rect 17635 20417 17647 20420
rect 17589 20411 17647 20417
rect 17604 20380 17632 20411
rect 17954 20408 17960 20420
rect 18012 20408 18018 20460
rect 18064 20457 18092 20488
rect 18601 20485 18613 20519
rect 18647 20485 18659 20519
rect 18601 20479 18659 20485
rect 18690 20476 18696 20528
rect 18748 20516 18754 20528
rect 22066 20516 22094 20544
rect 22186 20516 22192 20528
rect 18748 20488 18920 20516
rect 22066 20488 22192 20516
rect 18748 20476 18754 20488
rect 18049 20451 18107 20457
rect 18049 20417 18061 20451
rect 18095 20417 18107 20451
rect 18049 20411 18107 20417
rect 18782 20408 18788 20460
rect 18840 20408 18846 20460
rect 18892 20457 18920 20488
rect 22186 20476 22192 20488
rect 22244 20476 22250 20528
rect 23198 20476 23204 20528
rect 23256 20516 23262 20528
rect 23256 20488 23782 20516
rect 23256 20476 23262 20488
rect 18877 20451 18935 20457
rect 18877 20417 18889 20451
rect 18923 20417 18935 20451
rect 18877 20411 18935 20417
rect 19613 20451 19671 20457
rect 19613 20417 19625 20451
rect 19659 20448 19671 20451
rect 19794 20448 19800 20460
rect 19659 20420 19800 20448
rect 19659 20417 19671 20420
rect 19613 20411 19671 20417
rect 19794 20408 19800 20420
rect 19852 20408 19858 20460
rect 20990 20408 20996 20460
rect 21048 20408 21054 20460
rect 21269 20451 21327 20457
rect 21269 20417 21281 20451
rect 21315 20448 21327 20451
rect 22094 20448 22100 20460
rect 21315 20420 22100 20448
rect 21315 20417 21327 20420
rect 21269 20411 21327 20417
rect 22094 20408 22100 20420
rect 22152 20408 22158 20460
rect 22462 20408 22468 20460
rect 22520 20408 22526 20460
rect 22646 20408 22652 20460
rect 22704 20448 22710 20460
rect 23017 20451 23075 20457
rect 23017 20448 23029 20451
rect 22704 20420 23029 20448
rect 22704 20408 22710 20420
rect 23017 20417 23029 20420
rect 23063 20417 23075 20451
rect 23017 20411 23075 20417
rect 16531 20352 17080 20380
rect 17328 20352 17632 20380
rect 16531 20349 16543 20352
rect 16485 20343 16543 20349
rect 6917 20315 6975 20321
rect 6917 20281 6929 20315
rect 6963 20312 6975 20315
rect 7374 20312 7380 20324
rect 6963 20284 7380 20312
rect 6963 20281 6975 20284
rect 6917 20275 6975 20281
rect 7374 20272 7380 20284
rect 7432 20272 7438 20324
rect 7484 20284 8616 20312
rect 7484 20244 7512 20284
rect 6748 20216 7512 20244
rect 5629 20207 5687 20213
rect 7650 20204 7656 20256
rect 7708 20244 7714 20256
rect 8021 20247 8079 20253
rect 8021 20244 8033 20247
rect 7708 20216 8033 20244
rect 7708 20204 7714 20216
rect 8021 20213 8033 20216
rect 8067 20213 8079 20247
rect 8021 20207 8079 20213
rect 8110 20204 8116 20256
rect 8168 20244 8174 20256
rect 8588 20253 8616 20284
rect 15102 20272 15108 20324
rect 15160 20312 15166 20324
rect 16301 20315 16359 20321
rect 16301 20312 16313 20315
rect 15160 20284 16313 20312
rect 15160 20272 15166 20284
rect 16301 20281 16313 20284
rect 16347 20281 16359 20315
rect 16301 20275 16359 20281
rect 16666 20272 16672 20324
rect 16724 20312 16730 20324
rect 16761 20315 16819 20321
rect 16761 20312 16773 20315
rect 16724 20284 16773 20312
rect 16724 20272 16730 20284
rect 16761 20281 16773 20284
rect 16807 20281 16819 20315
rect 17052 20312 17080 20352
rect 18138 20340 18144 20392
rect 18196 20380 18202 20392
rect 19705 20383 19763 20389
rect 18196 20352 18644 20380
rect 18196 20340 18202 20352
rect 18616 20321 18644 20352
rect 19705 20349 19717 20383
rect 19751 20380 19763 20383
rect 20714 20380 20720 20392
rect 19751 20352 20720 20380
rect 19751 20349 19763 20352
rect 19705 20343 19763 20349
rect 20714 20340 20720 20352
rect 20772 20340 20778 20392
rect 20809 20383 20867 20389
rect 20809 20349 20821 20383
rect 20855 20380 20867 20383
rect 21174 20380 21180 20392
rect 20855 20352 21180 20380
rect 20855 20349 20867 20352
rect 20809 20343 20867 20349
rect 21174 20340 21180 20352
rect 21232 20340 21238 20392
rect 22557 20383 22615 20389
rect 22557 20349 22569 20383
rect 22603 20380 22615 20383
rect 22738 20380 22744 20392
rect 22603 20352 22744 20380
rect 22603 20349 22615 20352
rect 22557 20343 22615 20349
rect 22738 20340 22744 20352
rect 22796 20380 22802 20392
rect 23293 20383 23351 20389
rect 23293 20380 23305 20383
rect 22796 20352 23305 20380
rect 22796 20340 22802 20352
rect 23293 20349 23305 20352
rect 23339 20349 23351 20383
rect 23293 20343 23351 20349
rect 18601 20315 18659 20321
rect 17052 20284 18552 20312
rect 16761 20275 16819 20281
rect 8205 20247 8263 20253
rect 8205 20244 8217 20247
rect 8168 20216 8217 20244
rect 8168 20204 8174 20216
rect 8205 20213 8217 20216
rect 8251 20213 8263 20247
rect 8205 20207 8263 20213
rect 8573 20247 8631 20253
rect 8573 20213 8585 20247
rect 8619 20244 8631 20247
rect 9306 20244 9312 20256
rect 8619 20216 9312 20244
rect 8619 20213 8631 20216
rect 8573 20207 8631 20213
rect 9306 20204 9312 20216
rect 9364 20204 9370 20256
rect 13814 20204 13820 20256
rect 13872 20204 13878 20256
rect 15930 20204 15936 20256
rect 15988 20204 15994 20256
rect 18414 20204 18420 20256
rect 18472 20204 18478 20256
rect 18524 20244 18552 20284
rect 18601 20281 18613 20315
rect 18647 20281 18659 20315
rect 20901 20315 20959 20321
rect 20901 20312 20913 20315
rect 18601 20275 18659 20281
rect 18708 20284 20913 20312
rect 18708 20244 18736 20284
rect 20901 20281 20913 20284
rect 20947 20281 20959 20315
rect 20901 20275 20959 20281
rect 18524 20216 18736 20244
rect 19978 20204 19984 20256
rect 20036 20204 20042 20256
rect 20990 20204 20996 20256
rect 21048 20244 21054 20256
rect 22097 20247 22155 20253
rect 22097 20244 22109 20247
rect 21048 20216 22109 20244
rect 21048 20204 21054 20216
rect 22097 20213 22109 20216
rect 22143 20213 22155 20247
rect 22097 20207 22155 20213
rect 1104 20154 25208 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 25208 20154
rect 1104 20080 25208 20102
rect 11885 20043 11943 20049
rect 11885 20009 11897 20043
rect 11931 20040 11943 20043
rect 13446 20040 13452 20052
rect 11931 20012 13452 20040
rect 11931 20009 11943 20012
rect 11885 20003 11943 20009
rect 13446 20000 13452 20012
rect 13504 20000 13510 20052
rect 13814 20000 13820 20052
rect 13872 20000 13878 20052
rect 18782 20000 18788 20052
rect 18840 20040 18846 20052
rect 19245 20043 19303 20049
rect 19245 20040 19257 20043
rect 18840 20012 19257 20040
rect 18840 20000 18846 20012
rect 19245 20009 19257 20012
rect 19291 20009 19303 20043
rect 19245 20003 19303 20009
rect 19978 20000 19984 20052
rect 20036 20040 20042 20052
rect 20073 20043 20131 20049
rect 20073 20040 20085 20043
rect 20036 20012 20085 20040
rect 20036 20000 20042 20012
rect 20073 20009 20085 20012
rect 20119 20009 20131 20043
rect 20073 20003 20131 20009
rect 2774 19932 2780 19984
rect 2832 19972 2838 19984
rect 3418 19972 3424 19984
rect 2832 19944 3424 19972
rect 2832 19932 2838 19944
rect 3418 19932 3424 19944
rect 3476 19932 3482 19984
rect 8205 19975 8263 19981
rect 8205 19941 8217 19975
rect 8251 19972 8263 19975
rect 8386 19972 8392 19984
rect 8251 19944 8392 19972
rect 8251 19941 8263 19944
rect 8205 19935 8263 19941
rect 8386 19932 8392 19944
rect 8444 19972 8450 19984
rect 10137 19975 10195 19981
rect 8444 19944 9352 19972
rect 8444 19932 8450 19944
rect 1394 19864 1400 19916
rect 1452 19904 1458 19916
rect 2682 19904 2688 19916
rect 1452 19876 2688 19904
rect 1452 19864 1458 19876
rect 2682 19864 2688 19876
rect 2740 19904 2746 19916
rect 4893 19907 4951 19913
rect 2740 19876 3832 19904
rect 2740 19864 2746 19876
rect 3326 19836 3332 19848
rect 2806 19808 3332 19836
rect 3326 19796 3332 19808
rect 3384 19796 3390 19848
rect 3418 19796 3424 19848
rect 3476 19796 3482 19848
rect 3602 19796 3608 19848
rect 3660 19796 3666 19848
rect 3804 19845 3832 19876
rect 4893 19873 4905 19907
rect 4939 19904 4951 19907
rect 5442 19904 5448 19916
rect 4939 19876 5448 19904
rect 4939 19873 4951 19876
rect 4893 19867 4951 19873
rect 5442 19864 5448 19876
rect 5500 19864 5506 19916
rect 6362 19864 6368 19916
rect 6420 19864 6426 19916
rect 6641 19907 6699 19913
rect 6641 19873 6653 19907
rect 6687 19904 6699 19907
rect 7098 19904 7104 19916
rect 6687 19876 7104 19904
rect 6687 19873 6699 19876
rect 6641 19867 6699 19873
rect 7098 19864 7104 19876
rect 7156 19864 7162 19916
rect 7282 19864 7288 19916
rect 7340 19904 7346 19916
rect 9324 19913 9352 19944
rect 10137 19941 10149 19975
rect 10183 19972 10195 19975
rect 11514 19972 11520 19984
rect 10183 19944 11520 19972
rect 10183 19941 10195 19944
rect 10137 19935 10195 19941
rect 11514 19932 11520 19944
rect 11572 19932 11578 19984
rect 12066 19932 12072 19984
rect 12124 19932 12130 19984
rect 12161 19975 12219 19981
rect 12161 19941 12173 19975
rect 12207 19972 12219 19975
rect 12526 19972 12532 19984
rect 12207 19944 12532 19972
rect 12207 19941 12219 19944
rect 12161 19935 12219 19941
rect 9309 19907 9367 19913
rect 7340 19876 7972 19904
rect 7340 19864 7346 19876
rect 7944 19848 7972 19876
rect 9309 19873 9321 19907
rect 9355 19904 9367 19907
rect 9677 19907 9735 19913
rect 9677 19904 9689 19907
rect 9355 19876 9689 19904
rect 9355 19873 9367 19876
rect 9309 19867 9367 19873
rect 9677 19873 9689 19876
rect 9723 19873 9735 19907
rect 9677 19867 9735 19873
rect 11793 19907 11851 19913
rect 11793 19873 11805 19907
rect 11839 19904 11851 19907
rect 12084 19904 12112 19932
rect 11839 19876 12112 19904
rect 11839 19873 11851 19876
rect 11793 19867 11851 19873
rect 3789 19839 3847 19845
rect 3789 19805 3801 19839
rect 3835 19836 3847 19839
rect 4154 19836 4160 19848
rect 3835 19808 4160 19836
rect 3835 19805 3847 19808
rect 3789 19799 3847 19805
rect 4154 19796 4160 19808
rect 4212 19796 4218 19848
rect 5350 19836 5356 19848
rect 5092 19808 5356 19836
rect 1673 19771 1731 19777
rect 1673 19737 1685 19771
rect 1719 19737 1731 19771
rect 3237 19771 3295 19777
rect 3237 19768 3249 19771
rect 1673 19731 1731 19737
rect 2976 19740 3249 19768
rect 1688 19700 1716 19731
rect 2976 19700 3004 19740
rect 3237 19737 3249 19740
rect 3283 19737 3295 19771
rect 3237 19731 3295 19737
rect 4706 19728 4712 19780
rect 4764 19768 4770 19780
rect 4985 19771 5043 19777
rect 4985 19768 4997 19771
rect 4764 19740 4997 19768
rect 4764 19728 4770 19740
rect 4985 19737 4997 19740
rect 5031 19737 5043 19771
rect 4985 19731 5043 19737
rect 1688 19672 3004 19700
rect 3142 19660 3148 19712
rect 3200 19700 3206 19712
rect 4062 19700 4068 19712
rect 3200 19672 4068 19700
rect 3200 19660 3206 19672
rect 4062 19660 4068 19672
rect 4120 19700 4126 19712
rect 5092 19700 5120 19808
rect 5350 19796 5356 19808
rect 5408 19796 5414 19848
rect 7926 19796 7932 19848
rect 7984 19836 7990 19848
rect 8941 19839 8999 19845
rect 8941 19836 8953 19839
rect 7984 19808 8953 19836
rect 7984 19796 7990 19808
rect 8941 19805 8953 19808
rect 8987 19805 8999 19839
rect 8941 19799 8999 19805
rect 9125 19839 9183 19845
rect 9125 19805 9137 19839
rect 9171 19805 9183 19839
rect 9125 19799 9183 19805
rect 5258 19728 5264 19780
rect 5316 19768 5322 19780
rect 5445 19771 5503 19777
rect 5445 19768 5457 19771
rect 5316 19740 5457 19768
rect 5316 19728 5322 19740
rect 5445 19737 5457 19740
rect 5491 19768 5503 19771
rect 5810 19768 5816 19780
rect 5491 19740 5816 19768
rect 5491 19737 5503 19740
rect 5445 19731 5503 19737
rect 5810 19728 5816 19740
rect 5868 19728 5874 19780
rect 7098 19728 7104 19780
rect 7156 19728 7162 19780
rect 8202 19728 8208 19780
rect 8260 19768 8266 19780
rect 8573 19771 8631 19777
rect 8573 19768 8585 19771
rect 8260 19740 8585 19768
rect 8260 19728 8266 19740
rect 8573 19737 8585 19740
rect 8619 19768 8631 19771
rect 9140 19768 9168 19799
rect 9766 19796 9772 19848
rect 9824 19796 9830 19848
rect 8619 19740 9168 19768
rect 8619 19737 8631 19740
rect 8573 19731 8631 19737
rect 9306 19728 9312 19780
rect 9364 19768 9370 19780
rect 11808 19768 11836 19867
rect 11977 19839 12035 19845
rect 11977 19805 11989 19839
rect 12023 19805 12035 19839
rect 11977 19799 12035 19805
rect 12069 19839 12127 19845
rect 12069 19805 12081 19839
rect 12115 19836 12127 19839
rect 12176 19836 12204 19935
rect 12526 19932 12532 19944
rect 12584 19932 12590 19984
rect 13633 19907 13691 19913
rect 13633 19873 13645 19907
rect 13679 19904 13691 19907
rect 13832 19904 13860 20000
rect 15930 19932 15936 19984
rect 15988 19972 15994 19984
rect 15988 19944 20208 19972
rect 15988 19932 15994 19944
rect 13679 19876 13860 19904
rect 13679 19873 13691 19876
rect 13633 19867 13691 19873
rect 15838 19864 15844 19916
rect 15896 19904 15902 19916
rect 16485 19907 16543 19913
rect 15896 19876 16252 19904
rect 15896 19864 15902 19876
rect 12115 19808 12204 19836
rect 12115 19805 12127 19808
rect 12069 19799 12127 19805
rect 9364 19740 11836 19768
rect 9364 19728 9370 19740
rect 4120 19672 5120 19700
rect 4120 19660 4126 19672
rect 5994 19660 6000 19712
rect 6052 19700 6058 19712
rect 7282 19700 7288 19712
rect 6052 19672 7288 19700
rect 6052 19660 6058 19672
rect 7282 19660 7288 19672
rect 7340 19660 7346 19712
rect 7466 19660 7472 19712
rect 7524 19700 7530 19712
rect 8110 19700 8116 19712
rect 7524 19672 8116 19700
rect 7524 19660 7530 19672
rect 8110 19660 8116 19672
rect 8168 19700 8174 19712
rect 8389 19703 8447 19709
rect 8389 19700 8401 19703
rect 8168 19672 8401 19700
rect 8168 19660 8174 19672
rect 8389 19669 8401 19672
rect 8435 19669 8447 19703
rect 8389 19663 8447 19669
rect 8481 19703 8539 19709
rect 8481 19669 8493 19703
rect 8527 19700 8539 19703
rect 8662 19700 8668 19712
rect 8527 19672 8668 19700
rect 8527 19669 8539 19672
rect 8481 19663 8539 19669
rect 8662 19660 8668 19672
rect 8720 19660 8726 19712
rect 8757 19703 8815 19709
rect 8757 19669 8769 19703
rect 8803 19700 8815 19703
rect 9674 19700 9680 19712
rect 8803 19672 9680 19700
rect 8803 19669 8815 19672
rect 8757 19663 8815 19669
rect 9674 19660 9680 19672
rect 9732 19660 9738 19712
rect 11992 19700 12020 19799
rect 13906 19796 13912 19848
rect 13964 19796 13970 19848
rect 16224 19845 16252 19876
rect 16485 19873 16497 19907
rect 16531 19904 16543 19907
rect 17126 19904 17132 19916
rect 16531 19876 17132 19904
rect 16531 19873 16543 19876
rect 16485 19867 16543 19873
rect 17126 19864 17132 19876
rect 17184 19864 17190 19916
rect 18414 19864 18420 19916
rect 18472 19904 18478 19916
rect 20180 19913 20208 19944
rect 20165 19907 20223 19913
rect 18472 19876 20116 19904
rect 18472 19864 18478 19876
rect 16117 19839 16175 19845
rect 16117 19805 16129 19839
rect 16163 19805 16175 19839
rect 16117 19799 16175 19805
rect 16210 19839 16268 19845
rect 16210 19805 16222 19839
rect 16256 19805 16268 19839
rect 16210 19799 16268 19805
rect 13998 19768 14004 19780
rect 13202 19740 14004 19768
rect 13998 19728 14004 19740
rect 14056 19768 14062 19780
rect 14826 19768 14832 19780
rect 14056 19740 14832 19768
rect 14056 19728 14062 19740
rect 14826 19728 14832 19740
rect 14884 19728 14890 19780
rect 16132 19768 16160 19799
rect 19610 19796 19616 19848
rect 19668 19836 19674 19848
rect 20088 19845 20116 19876
rect 20165 19873 20177 19907
rect 20211 19873 20223 19907
rect 20165 19867 20223 19873
rect 19797 19839 19855 19845
rect 19797 19836 19809 19839
rect 19668 19808 19809 19836
rect 19668 19796 19674 19808
rect 19797 19805 19809 19808
rect 19843 19805 19855 19839
rect 19797 19799 19855 19805
rect 20073 19839 20131 19845
rect 20073 19805 20085 19839
rect 20119 19805 20131 19839
rect 20073 19799 20131 19805
rect 20349 19839 20407 19845
rect 20349 19805 20361 19839
rect 20395 19836 20407 19839
rect 20438 19836 20444 19848
rect 20395 19808 20444 19836
rect 20395 19805 20407 19808
rect 20349 19799 20407 19805
rect 20438 19796 20444 19808
rect 20496 19796 20502 19848
rect 16666 19768 16672 19780
rect 16132 19740 16672 19768
rect 16666 19728 16672 19740
rect 16724 19728 16730 19780
rect 19426 19728 19432 19780
rect 19484 19768 19490 19780
rect 22002 19768 22008 19780
rect 19484 19740 22008 19768
rect 19484 19728 19490 19740
rect 22002 19728 22008 19740
rect 22060 19728 22066 19780
rect 12710 19700 12716 19712
rect 11992 19672 12716 19700
rect 12710 19660 12716 19672
rect 12768 19660 12774 19712
rect 19886 19660 19892 19712
rect 19944 19700 19950 19712
rect 20533 19703 20591 19709
rect 20533 19700 20545 19703
rect 19944 19672 20545 19700
rect 19944 19660 19950 19672
rect 20533 19669 20545 19672
rect 20579 19669 20591 19703
rect 20533 19663 20591 19669
rect 1104 19610 25208 19632
rect 1104 19558 4874 19610
rect 4926 19558 4938 19610
rect 4990 19558 5002 19610
rect 5054 19558 5066 19610
rect 5118 19558 5130 19610
rect 5182 19558 25208 19610
rect 1104 19536 25208 19558
rect 2774 19456 2780 19508
rect 2832 19456 2838 19508
rect 2866 19456 2872 19508
rect 2924 19456 2930 19508
rect 3142 19496 3148 19508
rect 2976 19468 3148 19496
rect 2593 19431 2651 19437
rect 2593 19397 2605 19431
rect 2639 19428 2651 19431
rect 2976 19428 3004 19468
rect 3142 19456 3148 19468
rect 3200 19456 3206 19508
rect 7101 19499 7159 19505
rect 7101 19465 7113 19499
rect 7147 19496 7159 19499
rect 7190 19496 7196 19508
rect 7147 19468 7196 19496
rect 7147 19465 7159 19468
rect 7101 19459 7159 19465
rect 7190 19456 7196 19468
rect 7248 19456 7254 19508
rect 7285 19499 7343 19505
rect 7285 19465 7297 19499
rect 7331 19496 7343 19499
rect 9306 19496 9312 19508
rect 7331 19468 9312 19496
rect 7331 19465 7343 19468
rect 7285 19459 7343 19465
rect 9306 19456 9312 19468
rect 9364 19456 9370 19508
rect 10870 19456 10876 19508
rect 10928 19496 10934 19508
rect 12158 19496 12164 19508
rect 10928 19468 12164 19496
rect 10928 19456 10934 19468
rect 12158 19456 12164 19468
rect 12216 19496 12222 19508
rect 12269 19499 12327 19505
rect 12269 19496 12281 19499
rect 12216 19468 12281 19496
rect 12216 19456 12222 19468
rect 12269 19465 12281 19468
rect 12315 19465 12327 19499
rect 12269 19459 12327 19465
rect 12437 19499 12495 19505
rect 12437 19465 12449 19499
rect 12483 19496 12495 19499
rect 12729 19499 12787 19505
rect 12729 19496 12741 19499
rect 12483 19468 12741 19496
rect 12483 19465 12495 19468
rect 12437 19459 12495 19465
rect 12729 19465 12741 19468
rect 12775 19465 12787 19499
rect 12729 19459 12787 19465
rect 12897 19499 12955 19505
rect 12897 19465 12909 19499
rect 12943 19496 12955 19499
rect 13078 19496 13084 19508
rect 12943 19468 13084 19496
rect 12943 19465 12955 19468
rect 12897 19459 12955 19465
rect 13078 19456 13084 19468
rect 13136 19456 13142 19508
rect 16206 19456 16212 19508
rect 16264 19456 16270 19508
rect 17862 19456 17868 19508
rect 17920 19456 17926 19508
rect 17954 19456 17960 19508
rect 18012 19496 18018 19508
rect 18230 19496 18236 19508
rect 18012 19468 18236 19496
rect 18012 19456 18018 19468
rect 18230 19456 18236 19468
rect 18288 19456 18294 19508
rect 19518 19456 19524 19508
rect 19576 19456 19582 19508
rect 20717 19499 20775 19505
rect 20717 19496 20729 19499
rect 19996 19468 20729 19496
rect 2639 19400 3004 19428
rect 2639 19397 2651 19400
rect 2593 19391 2651 19397
rect 3418 19388 3424 19440
rect 3476 19428 3482 19440
rect 3605 19431 3663 19437
rect 3605 19428 3617 19431
rect 3476 19400 3617 19428
rect 3476 19388 3482 19400
rect 3605 19397 3617 19400
rect 3651 19397 3663 19431
rect 3605 19391 3663 19397
rect 3789 19431 3847 19437
rect 3789 19397 3801 19431
rect 3835 19428 3847 19431
rect 3835 19400 7236 19428
rect 3835 19397 3847 19400
rect 3789 19391 3847 19397
rect 3053 19363 3111 19369
rect 3053 19360 3065 19363
rect 2746 19332 3065 19360
rect 2222 19184 2228 19236
rect 2280 19184 2286 19236
rect 2593 19159 2651 19165
rect 2593 19125 2605 19159
rect 2639 19156 2651 19159
rect 2746 19156 2774 19332
rect 3053 19329 3065 19332
rect 3099 19360 3111 19363
rect 3099 19332 3924 19360
rect 3099 19329 3111 19332
rect 3053 19323 3111 19329
rect 3142 19252 3148 19304
rect 3200 19252 3206 19304
rect 3896 19292 3924 19332
rect 5442 19320 5448 19372
rect 5500 19360 5506 19372
rect 5629 19363 5687 19369
rect 5629 19360 5641 19363
rect 5500 19332 5641 19360
rect 5500 19320 5506 19332
rect 5629 19329 5641 19332
rect 5675 19329 5687 19363
rect 5629 19323 5687 19329
rect 5810 19320 5816 19372
rect 5868 19320 5874 19372
rect 5994 19320 6000 19372
rect 6052 19320 6058 19372
rect 6178 19320 6184 19372
rect 6236 19320 6242 19372
rect 6362 19320 6368 19372
rect 6420 19360 6426 19372
rect 6733 19363 6791 19369
rect 6733 19360 6745 19363
rect 6420 19332 6745 19360
rect 6420 19320 6426 19332
rect 6733 19329 6745 19332
rect 6779 19329 6791 19363
rect 7208 19360 7236 19400
rect 11422 19388 11428 19440
rect 11480 19428 11486 19440
rect 11882 19428 11888 19440
rect 11480 19400 11888 19428
rect 11480 19388 11486 19400
rect 11882 19388 11888 19400
rect 11940 19428 11946 19440
rect 12069 19431 12127 19437
rect 12069 19428 12081 19431
rect 11940 19400 12081 19428
rect 11940 19388 11946 19400
rect 12069 19397 12081 19400
rect 12115 19397 12127 19431
rect 12069 19391 12127 19397
rect 12526 19388 12532 19440
rect 12584 19388 12590 19440
rect 16025 19431 16083 19437
rect 16025 19397 16037 19431
rect 16071 19428 16083 19431
rect 16666 19428 16672 19440
rect 16071 19400 16672 19428
rect 16071 19397 16083 19400
rect 16025 19391 16083 19397
rect 7837 19363 7895 19369
rect 7837 19360 7849 19363
rect 7208 19332 7849 19360
rect 6733 19323 6791 19329
rect 7837 19329 7849 19332
rect 7883 19360 7895 19363
rect 8938 19360 8944 19372
rect 7883 19332 8944 19360
rect 7883 19329 7895 19332
rect 7837 19323 7895 19329
rect 5721 19295 5779 19301
rect 5721 19292 5733 19295
rect 3896 19264 5733 19292
rect 5721 19261 5733 19264
rect 5767 19261 5779 19295
rect 6748 19292 6776 19323
rect 8938 19320 8944 19332
rect 8996 19320 9002 19372
rect 9766 19320 9772 19372
rect 9824 19360 9830 19372
rect 9861 19363 9919 19369
rect 9861 19360 9873 19363
rect 9824 19332 9873 19360
rect 9824 19320 9830 19332
rect 9861 19329 9873 19332
rect 9907 19360 9919 19363
rect 14642 19360 14648 19372
rect 9907 19332 14648 19360
rect 9907 19329 9919 19332
rect 9861 19323 9919 19329
rect 14642 19320 14648 19332
rect 14700 19320 14706 19372
rect 15102 19320 15108 19372
rect 15160 19360 15166 19372
rect 15841 19363 15899 19369
rect 15841 19360 15853 19363
rect 15160 19332 15853 19360
rect 15160 19320 15166 19332
rect 15841 19329 15853 19332
rect 15887 19329 15899 19363
rect 15841 19323 15899 19329
rect 16117 19363 16175 19369
rect 16117 19329 16129 19363
rect 16163 19329 16175 19363
rect 16117 19323 16175 19329
rect 16209 19363 16267 19369
rect 16209 19329 16221 19363
rect 16255 19358 16267 19363
rect 16316 19358 16344 19400
rect 16666 19388 16672 19400
rect 16724 19388 16730 19440
rect 17880 19428 17908 19456
rect 19996 19428 20024 19468
rect 20717 19465 20729 19468
rect 20763 19496 20775 19499
rect 20806 19496 20812 19508
rect 20763 19468 20812 19496
rect 20763 19465 20775 19468
rect 20717 19459 20775 19465
rect 20806 19456 20812 19468
rect 20864 19456 20870 19508
rect 21821 19499 21879 19505
rect 21821 19465 21833 19499
rect 21867 19496 21879 19499
rect 22278 19496 22284 19508
rect 21867 19468 22284 19496
rect 21867 19465 21879 19468
rect 21821 19459 21879 19465
rect 22278 19456 22284 19468
rect 22336 19456 22342 19508
rect 17880 19400 20024 19428
rect 20162 19388 20168 19440
rect 20220 19428 20226 19440
rect 20220 19400 20944 19428
rect 20220 19388 20226 19400
rect 16255 19330 16344 19358
rect 16255 19329 16267 19330
rect 16209 19323 16267 19329
rect 8662 19292 8668 19304
rect 6748 19264 8668 19292
rect 5721 19255 5779 19261
rect 8662 19252 8668 19264
rect 8720 19292 8726 19304
rect 9953 19295 10011 19301
rect 8720 19264 9168 19292
rect 8720 19252 8726 19264
rect 3234 19184 3240 19236
rect 3292 19224 3298 19236
rect 3605 19227 3663 19233
rect 3605 19224 3617 19227
rect 3292 19196 3617 19224
rect 3292 19184 3298 19196
rect 3605 19193 3617 19196
rect 3651 19193 3663 19227
rect 3605 19187 3663 19193
rect 4154 19184 4160 19236
rect 4212 19224 4218 19236
rect 4614 19224 4620 19236
rect 4212 19196 4620 19224
rect 4212 19184 4218 19196
rect 4614 19184 4620 19196
rect 4672 19224 4678 19236
rect 5077 19227 5135 19233
rect 5077 19224 5089 19227
rect 4672 19196 5089 19224
rect 4672 19184 4678 19196
rect 5077 19193 5089 19196
rect 5123 19193 5135 19227
rect 5077 19187 5135 19193
rect 6181 19227 6239 19233
rect 6181 19193 6193 19227
rect 6227 19224 6239 19227
rect 6822 19224 6828 19236
rect 6227 19196 6828 19224
rect 6227 19193 6239 19196
rect 6181 19187 6239 19193
rect 6822 19184 6828 19196
rect 6880 19224 6886 19236
rect 6880 19196 7512 19224
rect 6880 19184 6886 19196
rect 2639 19128 2774 19156
rect 7285 19159 7343 19165
rect 2639 19125 2651 19128
rect 2593 19119 2651 19125
rect 7285 19125 7297 19159
rect 7331 19156 7343 19159
rect 7374 19156 7380 19168
rect 7331 19128 7380 19156
rect 7331 19125 7343 19128
rect 7285 19119 7343 19125
rect 7374 19116 7380 19128
rect 7432 19116 7438 19168
rect 7484 19156 7512 19196
rect 7650 19184 7656 19236
rect 7708 19184 7714 19236
rect 9140 19233 9168 19264
rect 9953 19261 9965 19295
rect 9999 19261 10011 19295
rect 9953 19255 10011 19261
rect 10229 19295 10287 19301
rect 10229 19261 10241 19295
rect 10275 19292 10287 19295
rect 10502 19292 10508 19304
rect 10275 19264 10508 19292
rect 10275 19261 10287 19264
rect 10229 19255 10287 19261
rect 9125 19227 9183 19233
rect 9125 19193 9137 19227
rect 9171 19193 9183 19227
rect 9125 19187 9183 19193
rect 9968 19156 9996 19255
rect 10502 19252 10508 19264
rect 10560 19252 10566 19304
rect 12434 19252 12440 19304
rect 12492 19292 12498 19304
rect 12710 19292 12716 19304
rect 12492 19264 12716 19292
rect 12492 19252 12498 19264
rect 12710 19252 12716 19264
rect 12768 19292 12774 19304
rect 13078 19292 13084 19304
rect 12768 19264 13084 19292
rect 12768 19252 12774 19264
rect 13078 19252 13084 19264
rect 13136 19252 13142 19304
rect 15194 19252 15200 19304
rect 15252 19292 15258 19304
rect 16132 19292 16160 19323
rect 16390 19320 16396 19372
rect 16448 19320 16454 19372
rect 19886 19320 19892 19372
rect 19944 19320 19950 19372
rect 20622 19320 20628 19372
rect 20680 19320 20686 19372
rect 20916 19369 20944 19400
rect 22002 19388 22008 19440
rect 22060 19388 22066 19440
rect 20901 19363 20959 19369
rect 20901 19329 20913 19363
rect 20947 19329 20959 19363
rect 20901 19323 20959 19329
rect 21266 19320 21272 19372
rect 21324 19320 21330 19372
rect 21453 19363 21511 19369
rect 21453 19329 21465 19363
rect 21499 19360 21511 19363
rect 22094 19360 22100 19372
rect 21499 19332 22100 19360
rect 21499 19329 21511 19332
rect 21453 19323 21511 19329
rect 22094 19320 22100 19332
rect 22152 19320 22158 19372
rect 16408 19292 16436 19320
rect 15252 19264 16436 19292
rect 19797 19295 19855 19301
rect 15252 19252 15258 19264
rect 19797 19261 19809 19295
rect 19843 19292 19855 19295
rect 20990 19292 20996 19304
rect 19843 19264 20996 19292
rect 19843 19261 19855 19264
rect 19797 19255 19855 19261
rect 20990 19252 20996 19264
rect 21048 19252 21054 19304
rect 21637 19227 21695 19233
rect 21637 19193 21649 19227
rect 21683 19224 21695 19227
rect 21683 19196 22048 19224
rect 21683 19193 21695 19196
rect 21637 19187 21695 19193
rect 7484 19128 9996 19156
rect 12066 19116 12072 19168
rect 12124 19156 12130 19168
rect 12253 19159 12311 19165
rect 12253 19156 12265 19159
rect 12124 19128 12265 19156
rect 12124 19116 12130 19128
rect 12253 19125 12265 19128
rect 12299 19125 12311 19159
rect 12253 19119 12311 19125
rect 12713 19159 12771 19165
rect 12713 19125 12725 19159
rect 12759 19156 12771 19159
rect 12802 19156 12808 19168
rect 12759 19128 12808 19156
rect 12759 19125 12771 19128
rect 12713 19119 12771 19125
rect 12802 19116 12808 19128
rect 12860 19116 12866 19168
rect 15657 19159 15715 19165
rect 15657 19125 15669 19159
rect 15703 19156 15715 19159
rect 15838 19156 15844 19168
rect 15703 19128 15844 19156
rect 15703 19125 15715 19128
rect 15657 19119 15715 19125
rect 15838 19116 15844 19128
rect 15896 19116 15902 19168
rect 19702 19116 19708 19168
rect 19760 19116 19766 19168
rect 20898 19116 20904 19168
rect 20956 19156 20962 19168
rect 22020 19165 22048 19196
rect 22370 19184 22376 19236
rect 22428 19184 22434 19236
rect 21085 19159 21143 19165
rect 21085 19156 21097 19159
rect 20956 19128 21097 19156
rect 20956 19116 20962 19128
rect 21085 19125 21097 19128
rect 21131 19125 21143 19159
rect 21085 19119 21143 19125
rect 22005 19159 22063 19165
rect 22005 19125 22017 19159
rect 22051 19125 22063 19159
rect 22005 19119 22063 19125
rect 1104 19066 25208 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 25208 19066
rect 1104 18992 25208 19014
rect 3142 18912 3148 18964
rect 3200 18952 3206 18964
rect 3927 18955 3985 18961
rect 3927 18952 3939 18955
rect 3200 18924 3939 18952
rect 3200 18912 3206 18924
rect 3927 18921 3939 18924
rect 3973 18921 3985 18955
rect 3927 18915 3985 18921
rect 4798 18912 4804 18964
rect 4856 18952 4862 18964
rect 6086 18952 6092 18964
rect 4856 18924 6092 18952
rect 4856 18912 4862 18924
rect 6086 18912 6092 18924
rect 6144 18912 6150 18964
rect 7558 18912 7564 18964
rect 7616 18952 7622 18964
rect 8481 18955 8539 18961
rect 8481 18952 8493 18955
rect 7616 18924 8493 18952
rect 7616 18912 7622 18924
rect 8481 18921 8493 18924
rect 8527 18921 8539 18955
rect 8481 18915 8539 18921
rect 9858 18912 9864 18964
rect 9916 18952 9922 18964
rect 9916 18924 12388 18952
rect 9916 18912 9922 18924
rect 3326 18844 3332 18896
rect 3384 18884 3390 18896
rect 3384 18856 3740 18884
rect 3384 18844 3390 18856
rect 3602 18816 3608 18828
rect 3252 18788 3608 18816
rect 3252 18760 3280 18788
rect 3602 18776 3608 18788
rect 3660 18776 3666 18828
rect 3712 18816 3740 18856
rect 8294 18844 8300 18896
rect 8352 18884 8358 18896
rect 8941 18887 8999 18893
rect 8941 18884 8953 18887
rect 8352 18856 8953 18884
rect 8352 18844 8358 18856
rect 8941 18853 8953 18856
rect 8987 18853 8999 18887
rect 9306 18884 9312 18896
rect 8941 18847 8999 18853
rect 9140 18856 9312 18884
rect 4798 18816 4804 18828
rect 3712 18788 4804 18816
rect 4798 18776 4804 18788
rect 4856 18776 4862 18828
rect 5721 18819 5779 18825
rect 5721 18785 5733 18819
rect 5767 18816 5779 18819
rect 6362 18816 6368 18828
rect 5767 18788 6368 18816
rect 5767 18785 5779 18788
rect 5721 18779 5779 18785
rect 6362 18776 6368 18788
rect 6420 18816 6426 18828
rect 6549 18819 6607 18825
rect 6549 18816 6561 18819
rect 6420 18788 6561 18816
rect 6420 18776 6426 18788
rect 6549 18785 6561 18788
rect 6595 18785 6607 18819
rect 6549 18779 6607 18785
rect 6822 18776 6828 18828
rect 6880 18776 6886 18828
rect 8665 18819 8723 18825
rect 8665 18785 8677 18819
rect 8711 18816 8723 18819
rect 9140 18816 9168 18856
rect 9306 18844 9312 18856
rect 9364 18844 9370 18896
rect 9585 18887 9643 18893
rect 9585 18853 9597 18887
rect 9631 18853 9643 18887
rect 9585 18847 9643 18853
rect 8711 18788 9168 18816
rect 8711 18785 8723 18788
rect 8665 18779 8723 18785
rect 9214 18776 9220 18828
rect 9272 18816 9278 18828
rect 9600 18816 9628 18847
rect 11882 18844 11888 18896
rect 11940 18884 11946 18896
rect 12360 18884 12388 18924
rect 12434 18912 12440 18964
rect 12492 18912 12498 18964
rect 12710 18912 12716 18964
rect 12768 18912 12774 18964
rect 15194 18912 15200 18964
rect 15252 18912 15258 18964
rect 15746 18952 15752 18964
rect 15488 18924 15752 18952
rect 15488 18893 15516 18924
rect 15746 18912 15752 18924
rect 15804 18912 15810 18964
rect 15841 18955 15899 18961
rect 15841 18921 15853 18955
rect 15887 18952 15899 18955
rect 15930 18952 15936 18964
rect 15887 18924 15936 18952
rect 15887 18921 15899 18924
rect 15841 18915 15899 18921
rect 15930 18912 15936 18924
rect 15988 18912 15994 18964
rect 17773 18955 17831 18961
rect 17773 18921 17785 18955
rect 17819 18952 17831 18955
rect 18782 18952 18788 18964
rect 17819 18924 18788 18952
rect 17819 18921 17831 18924
rect 17773 18915 17831 18921
rect 18782 18912 18788 18924
rect 18840 18912 18846 18964
rect 18874 18912 18880 18964
rect 18932 18961 18938 18964
rect 18932 18915 18944 18961
rect 18932 18912 18938 18915
rect 19058 18912 19064 18964
rect 19116 18952 19122 18964
rect 19245 18955 19303 18961
rect 19245 18952 19257 18955
rect 19116 18924 19257 18952
rect 19116 18912 19122 18924
rect 19245 18921 19257 18924
rect 19291 18921 19303 18955
rect 19245 18915 19303 18921
rect 19702 18912 19708 18964
rect 19760 18912 19766 18964
rect 20162 18912 20168 18964
rect 20220 18952 20226 18964
rect 20257 18955 20315 18961
rect 20257 18952 20269 18955
rect 20220 18924 20269 18952
rect 20220 18912 20226 18924
rect 20257 18921 20269 18924
rect 20303 18921 20315 18955
rect 20257 18915 20315 18921
rect 20898 18912 20904 18964
rect 20956 18912 20962 18964
rect 21729 18955 21787 18961
rect 21729 18921 21741 18955
rect 21775 18952 21787 18955
rect 22370 18952 22376 18964
rect 21775 18924 22376 18952
rect 21775 18921 21787 18924
rect 21729 18915 21787 18921
rect 22370 18912 22376 18924
rect 22428 18912 22434 18964
rect 12529 18887 12587 18893
rect 12529 18884 12541 18887
rect 11940 18856 12312 18884
rect 12360 18856 12541 18884
rect 11940 18844 11946 18856
rect 9272 18788 9628 18816
rect 12284 18816 12312 18856
rect 12529 18853 12541 18856
rect 12575 18853 12587 18887
rect 12529 18847 12587 18853
rect 15381 18887 15439 18893
rect 15381 18853 15393 18887
rect 15427 18884 15439 18887
rect 15473 18887 15531 18893
rect 15473 18884 15485 18887
rect 15427 18856 15485 18884
rect 15427 18853 15439 18856
rect 15381 18847 15439 18853
rect 15473 18853 15485 18856
rect 15519 18853 15531 18887
rect 15473 18847 15531 18853
rect 15654 18844 15660 18896
rect 15712 18884 15718 18896
rect 16025 18887 16083 18893
rect 16025 18884 16037 18887
rect 15712 18856 16037 18884
rect 15712 18844 15718 18856
rect 16025 18853 16037 18856
rect 16071 18853 16083 18887
rect 16025 18847 16083 18853
rect 16669 18887 16727 18893
rect 16669 18853 16681 18887
rect 16715 18884 16727 18887
rect 20441 18887 20499 18893
rect 16715 18856 19564 18884
rect 16715 18853 16727 18856
rect 16669 18847 16727 18853
rect 12284 18788 13400 18816
rect 9272 18776 9278 18788
rect 2961 18751 3019 18757
rect 2961 18717 2973 18751
rect 3007 18748 3019 18751
rect 3050 18748 3056 18760
rect 3007 18720 3056 18748
rect 3007 18717 3019 18720
rect 2961 18711 3019 18717
rect 3050 18708 3056 18720
rect 3108 18708 3114 18760
rect 3142 18708 3148 18760
rect 3200 18708 3206 18760
rect 3234 18708 3240 18760
rect 3292 18708 3298 18760
rect 3329 18751 3387 18757
rect 3329 18717 3341 18751
rect 3375 18748 3387 18751
rect 3375 18720 4200 18748
rect 3375 18717 3387 18720
rect 3329 18711 3387 18717
rect 2222 18640 2228 18692
rect 2280 18680 2286 18692
rect 3344 18680 3372 18711
rect 2280 18652 3372 18680
rect 2280 18640 2286 18652
rect 3605 18615 3663 18621
rect 3605 18581 3617 18615
rect 3651 18612 3663 18615
rect 3694 18612 3700 18624
rect 3651 18584 3700 18612
rect 3651 18581 3663 18584
rect 3605 18575 3663 18581
rect 3694 18572 3700 18584
rect 3752 18572 3758 18624
rect 4172 18612 4200 18720
rect 5350 18708 5356 18760
rect 5408 18708 5414 18760
rect 8389 18751 8447 18757
rect 8389 18717 8401 18751
rect 8435 18748 8447 18751
rect 8754 18748 8760 18760
rect 8435 18720 8760 18748
rect 8435 18717 8447 18720
rect 8389 18711 8447 18717
rect 8754 18708 8760 18720
rect 8812 18708 8818 18760
rect 8846 18708 8852 18760
rect 8904 18748 8910 18760
rect 9309 18751 9367 18757
rect 9309 18748 9321 18751
rect 8904 18720 9321 18748
rect 8904 18708 8910 18720
rect 9309 18717 9321 18720
rect 9355 18717 9367 18751
rect 9309 18711 9367 18717
rect 9585 18751 9643 18757
rect 9585 18717 9597 18751
rect 9631 18717 9643 18751
rect 9585 18711 9643 18717
rect 4798 18640 4804 18692
rect 4856 18640 4862 18692
rect 8110 18680 8116 18692
rect 8050 18652 8116 18680
rect 8110 18640 8116 18652
rect 8168 18640 8174 18692
rect 8665 18683 8723 18689
rect 8665 18649 8677 18683
rect 8711 18680 8723 18683
rect 9600 18680 9628 18711
rect 9674 18708 9680 18760
rect 9732 18748 9738 18760
rect 9769 18751 9827 18757
rect 9769 18748 9781 18751
rect 9732 18720 9781 18748
rect 9732 18708 9738 18720
rect 9769 18717 9781 18720
rect 9815 18717 9827 18751
rect 9769 18711 9827 18717
rect 8711 18652 9628 18680
rect 8711 18649 8723 18652
rect 8665 18643 8723 18649
rect 5258 18612 5264 18624
rect 4172 18584 5264 18612
rect 5258 18572 5264 18584
rect 5316 18572 5322 18624
rect 7098 18572 7104 18624
rect 7156 18612 7162 18624
rect 8128 18612 8156 18640
rect 7156 18584 8156 18612
rect 8297 18615 8355 18621
rect 7156 18572 7162 18584
rect 8297 18581 8309 18615
rect 8343 18612 8355 18615
rect 8386 18612 8392 18624
rect 8343 18584 8392 18612
rect 8343 18581 8355 18584
rect 8297 18575 8355 18581
rect 8386 18572 8392 18584
rect 8444 18572 8450 18624
rect 9784 18612 9812 18711
rect 12066 18708 12072 18760
rect 12124 18708 12130 18760
rect 12158 18708 12164 18760
rect 12216 18708 12222 18760
rect 12268 18720 12756 18748
rect 10962 18640 10968 18692
rect 11020 18680 11026 18692
rect 12268 18680 12296 18720
rect 12728 18689 12756 18720
rect 13078 18708 13084 18760
rect 13136 18708 13142 18760
rect 13372 18757 13400 18788
rect 16114 18776 16120 18828
rect 16172 18816 16178 18828
rect 16209 18819 16267 18825
rect 16209 18816 16221 18819
rect 16172 18788 16221 18816
rect 16172 18776 16178 18788
rect 16209 18785 16221 18788
rect 16255 18785 16267 18819
rect 16209 18779 16267 18785
rect 17402 18776 17408 18828
rect 17460 18776 17466 18828
rect 18325 18819 18383 18825
rect 18325 18785 18337 18819
rect 18371 18785 18383 18819
rect 18325 18779 18383 18785
rect 18601 18819 18659 18825
rect 18601 18785 18613 18819
rect 18647 18816 18659 18819
rect 19337 18819 19395 18825
rect 19337 18816 19349 18819
rect 18647 18788 19349 18816
rect 18647 18785 18659 18788
rect 18601 18779 18659 18785
rect 19337 18785 19349 18788
rect 19383 18785 19395 18819
rect 19337 18779 19395 18785
rect 13357 18751 13415 18757
rect 13357 18717 13369 18751
rect 13403 18748 13415 18751
rect 13630 18748 13636 18760
rect 13403 18720 13636 18748
rect 13403 18717 13415 18720
rect 13357 18711 13415 18717
rect 13630 18708 13636 18720
rect 13688 18708 13694 18760
rect 15746 18708 15752 18760
rect 15804 18748 15810 18760
rect 15804 18720 15976 18748
rect 15804 18708 15810 18720
rect 11020 18652 12296 18680
rect 12713 18683 12771 18689
rect 11020 18640 11026 18652
rect 12713 18649 12725 18683
rect 12759 18649 12771 18683
rect 13446 18680 13452 18692
rect 12713 18643 12771 18649
rect 12820 18652 13452 18680
rect 12820 18624 12848 18652
rect 13446 18640 13452 18652
rect 13504 18680 13510 18692
rect 13541 18683 13599 18689
rect 13541 18680 13553 18683
rect 13504 18652 13553 18680
rect 13504 18640 13510 18652
rect 13541 18649 13553 18652
rect 13587 18649 13599 18683
rect 13541 18643 13599 18649
rect 15013 18683 15071 18689
rect 15013 18649 15025 18683
rect 15059 18649 15071 18683
rect 15013 18643 15071 18649
rect 12253 18615 12311 18621
rect 12253 18612 12265 18615
rect 9784 18584 12265 18612
rect 12253 18581 12265 18584
rect 12299 18612 12311 18615
rect 12802 18612 12808 18624
rect 12299 18584 12808 18612
rect 12299 18581 12311 18584
rect 12253 18575 12311 18581
rect 12802 18572 12808 18584
rect 12860 18572 12866 18624
rect 12894 18572 12900 18624
rect 12952 18612 12958 18624
rect 13173 18615 13231 18621
rect 13173 18612 13185 18615
rect 12952 18584 13185 18612
rect 12952 18572 12958 18584
rect 13173 18581 13185 18584
rect 13219 18581 13231 18615
rect 15028 18612 15056 18643
rect 15102 18640 15108 18692
rect 15160 18680 15166 18692
rect 15213 18683 15271 18689
rect 15213 18680 15225 18683
rect 15160 18652 15225 18680
rect 15160 18640 15166 18652
rect 15213 18649 15225 18652
rect 15259 18649 15271 18683
rect 15213 18643 15271 18649
rect 15838 18640 15844 18692
rect 15896 18640 15902 18692
rect 15948 18680 15976 18720
rect 16022 18708 16028 18760
rect 16080 18748 16086 18760
rect 16301 18751 16359 18757
rect 16301 18748 16313 18751
rect 16080 18720 16313 18748
rect 16080 18708 16086 18720
rect 16301 18717 16313 18720
rect 16347 18717 16359 18751
rect 16301 18711 16359 18717
rect 17497 18751 17555 18757
rect 17497 18717 17509 18751
rect 17543 18748 17555 18751
rect 17770 18748 17776 18760
rect 17543 18720 17776 18748
rect 17543 18717 17555 18720
rect 17497 18711 17555 18717
rect 17770 18708 17776 18720
rect 17828 18708 17834 18760
rect 18230 18708 18236 18760
rect 18288 18708 18294 18760
rect 16761 18683 16819 18689
rect 16761 18680 16773 18683
rect 15948 18652 16773 18680
rect 16761 18649 16773 18652
rect 16807 18649 16819 18683
rect 16761 18643 16819 18649
rect 16945 18683 17003 18689
rect 16945 18649 16957 18683
rect 16991 18680 17003 18683
rect 17034 18680 17040 18692
rect 16991 18652 17040 18680
rect 16991 18649 17003 18652
rect 16945 18643 17003 18649
rect 17034 18640 17040 18652
rect 17092 18680 17098 18692
rect 18046 18680 18052 18692
rect 17092 18652 18052 18680
rect 17092 18640 17098 18652
rect 18046 18640 18052 18652
rect 18104 18640 18110 18692
rect 18340 18680 18368 18779
rect 18690 18708 18696 18760
rect 18748 18748 18754 18760
rect 19536 18757 19564 18856
rect 20441 18853 20453 18887
rect 20487 18884 20499 18887
rect 20533 18887 20591 18893
rect 20533 18884 20545 18887
rect 20487 18856 20545 18884
rect 20487 18853 20499 18856
rect 20441 18847 20499 18853
rect 20533 18853 20545 18856
rect 20579 18884 20591 18887
rect 21266 18884 21272 18896
rect 20579 18856 21272 18884
rect 20579 18853 20591 18856
rect 20533 18847 20591 18853
rect 21266 18844 21272 18856
rect 21324 18844 21330 18896
rect 20622 18776 20628 18828
rect 20680 18816 20686 18828
rect 20680 18788 21588 18816
rect 20680 18776 20686 18788
rect 19521 18751 19579 18757
rect 18748 18720 19104 18748
rect 18748 18708 18754 18720
rect 19076 18689 19104 18720
rect 19521 18717 19533 18751
rect 19567 18717 19579 18751
rect 19521 18711 19579 18717
rect 20162 18708 20168 18760
rect 20220 18748 20226 18760
rect 21560 18757 21588 18788
rect 22278 18776 22284 18828
rect 22336 18776 22342 18828
rect 21361 18751 21419 18757
rect 21361 18748 21373 18751
rect 20220 18720 21373 18748
rect 20220 18708 20226 18720
rect 21361 18717 21373 18720
rect 21407 18717 21419 18751
rect 21361 18711 21419 18717
rect 21545 18751 21603 18757
rect 21545 18717 21557 18751
rect 21591 18717 21603 18751
rect 21545 18711 21603 18717
rect 21634 18708 21640 18760
rect 21692 18748 21698 18760
rect 22005 18751 22063 18757
rect 22005 18748 22017 18751
rect 21692 18720 22017 18748
rect 21692 18708 21698 18720
rect 22005 18717 22017 18720
rect 22051 18717 22063 18751
rect 22005 18711 22063 18717
rect 19061 18683 19119 18689
rect 18340 18652 19012 18680
rect 16666 18612 16672 18624
rect 15028 18584 16672 18612
rect 13173 18575 13231 18581
rect 16666 18572 16672 18584
rect 16724 18572 16730 18624
rect 16850 18572 16856 18624
rect 16908 18612 16914 18624
rect 18708 18621 18736 18652
rect 18874 18621 18880 18624
rect 17129 18615 17187 18621
rect 17129 18612 17141 18615
rect 16908 18584 17141 18612
rect 16908 18572 16914 18584
rect 17129 18581 17141 18584
rect 17175 18581 17187 18615
rect 17129 18575 17187 18581
rect 18693 18615 18751 18621
rect 18693 18581 18705 18615
rect 18739 18581 18751 18615
rect 18693 18575 18751 18581
rect 18861 18615 18880 18621
rect 18861 18581 18873 18615
rect 18861 18575 18880 18581
rect 18874 18572 18880 18575
rect 18932 18572 18938 18624
rect 18984 18612 19012 18652
rect 19061 18649 19073 18683
rect 19107 18680 19119 18683
rect 19150 18680 19156 18692
rect 19107 18652 19156 18680
rect 19107 18649 19119 18652
rect 19061 18643 19119 18649
rect 19150 18640 19156 18652
rect 19208 18640 19214 18692
rect 19245 18683 19303 18689
rect 19245 18649 19257 18683
rect 19291 18680 19303 18683
rect 19978 18680 19984 18692
rect 19291 18652 19984 18680
rect 19291 18649 19303 18652
rect 19245 18643 19303 18649
rect 19978 18640 19984 18652
rect 20036 18640 20042 18692
rect 20073 18683 20131 18689
rect 20073 18649 20085 18683
rect 20119 18649 20131 18683
rect 20073 18643 20131 18649
rect 19518 18612 19524 18624
rect 18984 18584 19524 18612
rect 19518 18572 19524 18584
rect 19576 18572 19582 18624
rect 20088 18612 20116 18643
rect 20254 18640 20260 18692
rect 20312 18689 20318 18692
rect 20312 18683 20347 18689
rect 20335 18680 20347 18683
rect 20622 18680 20628 18692
rect 20335 18652 20628 18680
rect 20335 18649 20347 18652
rect 20312 18643 20347 18649
rect 20312 18640 20318 18643
rect 20622 18640 20628 18652
rect 20680 18640 20686 18692
rect 20714 18640 20720 18692
rect 20772 18680 20778 18692
rect 20772 18652 21128 18680
rect 20772 18640 20778 18652
rect 21100 18624 21128 18652
rect 21174 18640 21180 18692
rect 21232 18640 21238 18692
rect 21453 18683 21511 18689
rect 21453 18649 21465 18683
rect 21499 18680 21511 18683
rect 21499 18652 21864 18680
rect 21499 18649 21511 18652
rect 21453 18643 21511 18649
rect 20806 18612 20812 18624
rect 20088 18584 20812 18612
rect 20806 18572 20812 18584
rect 20864 18572 20870 18624
rect 20898 18572 20904 18624
rect 20956 18572 20962 18624
rect 21082 18572 21088 18624
rect 21140 18572 21146 18624
rect 21836 18612 21864 18652
rect 23290 18640 23296 18692
rect 23348 18640 23354 18692
rect 22094 18612 22100 18624
rect 21836 18584 22100 18612
rect 22094 18572 22100 18584
rect 22152 18612 22158 18624
rect 23753 18615 23811 18621
rect 23753 18612 23765 18615
rect 22152 18584 23765 18612
rect 22152 18572 22158 18584
rect 23753 18581 23765 18584
rect 23799 18581 23811 18615
rect 23753 18575 23811 18581
rect 1104 18522 25208 18544
rect 1104 18470 4874 18522
rect 4926 18470 4938 18522
rect 4990 18470 5002 18522
rect 5054 18470 5066 18522
rect 5118 18470 5130 18522
rect 5182 18470 25208 18522
rect 1104 18448 25208 18470
rect 2961 18411 3019 18417
rect 2961 18377 2973 18411
rect 3007 18408 3019 18411
rect 3142 18408 3148 18420
rect 3007 18380 3148 18408
rect 3007 18377 3019 18380
rect 2961 18371 3019 18377
rect 3142 18368 3148 18380
rect 3200 18368 3206 18420
rect 5350 18368 5356 18420
rect 5408 18368 5414 18420
rect 7285 18411 7343 18417
rect 7285 18377 7297 18411
rect 7331 18408 7343 18411
rect 7374 18408 7380 18420
rect 7331 18380 7380 18408
rect 7331 18377 7343 18380
rect 7285 18371 7343 18377
rect 7374 18368 7380 18380
rect 7432 18368 7438 18420
rect 8110 18368 8116 18420
rect 8168 18368 8174 18420
rect 8754 18368 8760 18420
rect 8812 18408 8818 18420
rect 10413 18411 10471 18417
rect 10413 18408 10425 18411
rect 8812 18380 10425 18408
rect 8812 18368 8818 18380
rect 10413 18377 10425 18380
rect 10459 18377 10471 18411
rect 10413 18371 10471 18377
rect 10594 18368 10600 18420
rect 10652 18408 10658 18420
rect 11701 18411 11759 18417
rect 11701 18408 11713 18411
rect 10652 18380 11713 18408
rect 10652 18368 10658 18380
rect 11701 18377 11713 18380
rect 11747 18377 11759 18411
rect 11701 18371 11759 18377
rect 11885 18411 11943 18417
rect 11885 18377 11897 18411
rect 11931 18408 11943 18411
rect 12897 18411 12955 18417
rect 12897 18408 12909 18411
rect 11931 18380 12909 18408
rect 11931 18377 11943 18380
rect 11885 18371 11943 18377
rect 12897 18377 12909 18380
rect 12943 18377 12955 18411
rect 12897 18371 12955 18377
rect 13262 18368 13268 18420
rect 13320 18368 13326 18420
rect 14461 18411 14519 18417
rect 14461 18377 14473 18411
rect 14507 18408 14519 18411
rect 15102 18408 15108 18420
rect 14507 18380 15108 18408
rect 14507 18377 14519 18380
rect 14461 18371 14519 18377
rect 15102 18368 15108 18380
rect 15160 18408 15166 18420
rect 16945 18411 17003 18417
rect 16945 18408 16957 18411
rect 15160 18380 16957 18408
rect 15160 18368 15166 18380
rect 16945 18377 16957 18380
rect 16991 18377 17003 18411
rect 16945 18371 17003 18377
rect 17034 18368 17040 18420
rect 17092 18368 17098 18420
rect 19521 18411 19579 18417
rect 19521 18408 19533 18411
rect 17512 18380 19533 18408
rect 3694 18300 3700 18352
rect 3752 18300 3758 18352
rect 4982 18340 4988 18352
rect 4922 18312 4988 18340
rect 4982 18300 4988 18312
rect 5040 18340 5046 18352
rect 7098 18340 7104 18352
rect 5040 18312 7104 18340
rect 5040 18300 5046 18312
rect 7098 18300 7104 18312
rect 7156 18300 7162 18352
rect 7466 18300 7472 18352
rect 7524 18300 7530 18352
rect 7653 18343 7711 18349
rect 7653 18309 7665 18343
rect 7699 18340 7711 18343
rect 7926 18340 7932 18352
rect 7699 18312 7932 18340
rect 7699 18309 7711 18312
rect 7653 18303 7711 18309
rect 7926 18300 7932 18312
rect 7984 18300 7990 18352
rect 8941 18343 8999 18349
rect 8941 18309 8953 18343
rect 8987 18340 8999 18343
rect 9214 18340 9220 18352
rect 8987 18312 9220 18340
rect 8987 18309 8999 18312
rect 8941 18303 8999 18309
rect 9214 18300 9220 18312
rect 9272 18300 9278 18352
rect 10962 18300 10968 18352
rect 11020 18300 11026 18352
rect 11146 18300 11152 18352
rect 11204 18340 11210 18352
rect 12158 18340 12164 18352
rect 11204 18312 12164 18340
rect 11204 18300 11210 18312
rect 12158 18300 12164 18312
rect 12216 18300 12222 18352
rect 12434 18300 12440 18352
rect 12492 18300 12498 18352
rect 12653 18343 12711 18349
rect 12653 18309 12665 18343
rect 12699 18340 12711 18343
rect 13541 18343 13599 18349
rect 13541 18340 13553 18343
rect 12699 18312 13553 18340
rect 12699 18309 12711 18312
rect 12653 18303 12711 18309
rect 2866 18232 2872 18284
rect 2924 18232 2930 18284
rect 3053 18275 3111 18281
rect 3053 18241 3065 18275
rect 3099 18272 3111 18275
rect 3234 18272 3240 18284
rect 3099 18244 3240 18272
rect 3099 18241 3111 18244
rect 3053 18235 3111 18241
rect 3234 18232 3240 18244
rect 3292 18232 3298 18284
rect 6086 18232 6092 18284
rect 6144 18272 6150 18284
rect 7837 18275 7895 18281
rect 7837 18272 7849 18275
rect 6144 18244 7849 18272
rect 6144 18232 6150 18244
rect 7837 18241 7849 18244
rect 7883 18241 7895 18275
rect 7837 18235 7895 18241
rect 8662 18232 8668 18284
rect 8720 18232 8726 18284
rect 10042 18232 10048 18284
rect 10100 18232 10106 18284
rect 11333 18275 11391 18281
rect 11333 18241 11345 18275
rect 11379 18272 11391 18275
rect 12253 18275 12311 18281
rect 12253 18272 12265 18275
rect 11379 18244 12265 18272
rect 11379 18241 11391 18244
rect 11333 18235 11391 18241
rect 12253 18241 12265 18244
rect 12299 18272 12311 18275
rect 12897 18275 12955 18281
rect 12299 18244 12434 18272
rect 12299 18241 12311 18244
rect 12253 18235 12311 18241
rect 2774 18164 2780 18216
rect 2832 18204 2838 18216
rect 3421 18207 3479 18213
rect 3421 18204 3433 18207
rect 2832 18176 3433 18204
rect 2832 18164 2838 18176
rect 3421 18173 3433 18176
rect 3467 18173 3479 18207
rect 5905 18207 5963 18213
rect 5905 18204 5917 18207
rect 3421 18167 3479 18173
rect 3528 18176 5917 18204
rect 3418 18028 3424 18080
rect 3476 18068 3482 18080
rect 3528 18068 3556 18176
rect 5905 18173 5917 18176
rect 5951 18173 5963 18207
rect 5905 18167 5963 18173
rect 12406 18136 12434 18244
rect 12897 18241 12909 18275
rect 12943 18241 12955 18275
rect 13004 18270 13032 18312
rect 13541 18309 13553 18312
rect 13587 18340 13599 18343
rect 13587 18312 13768 18340
rect 13587 18309 13599 18312
rect 13541 18303 13599 18309
rect 13081 18275 13139 18281
rect 13081 18270 13093 18275
rect 13004 18242 13093 18270
rect 12897 18235 12955 18241
rect 13081 18241 13093 18242
rect 13127 18241 13139 18275
rect 13081 18235 13139 18241
rect 12912 18204 12940 18235
rect 13170 18232 13176 18284
rect 13228 18270 13234 18284
rect 13228 18242 13271 18270
rect 13228 18232 13234 18242
rect 13446 18232 13452 18284
rect 13504 18232 13510 18284
rect 13630 18232 13636 18284
rect 13688 18232 13694 18284
rect 13740 18281 13768 18312
rect 15470 18300 15476 18352
rect 15528 18300 15534 18352
rect 15654 18300 15660 18352
rect 15712 18340 15718 18352
rect 15933 18343 15991 18349
rect 15933 18340 15945 18343
rect 15712 18312 15945 18340
rect 15712 18300 15718 18312
rect 15933 18309 15945 18312
rect 15979 18309 15991 18343
rect 15933 18303 15991 18309
rect 16666 18300 16672 18352
rect 16724 18340 16730 18352
rect 17512 18349 17540 18380
rect 19521 18377 19533 18380
rect 19567 18408 19579 18411
rect 19610 18408 19616 18420
rect 19567 18380 19616 18408
rect 19567 18377 19579 18380
rect 19521 18371 19579 18377
rect 19610 18368 19616 18380
rect 19668 18368 19674 18420
rect 19978 18368 19984 18420
rect 20036 18408 20042 18420
rect 21821 18411 21879 18417
rect 21821 18408 21833 18411
rect 20036 18380 21833 18408
rect 20036 18368 20042 18380
rect 21821 18377 21833 18380
rect 21867 18377 21879 18411
rect 21821 18371 21879 18377
rect 17497 18343 17555 18349
rect 17497 18340 17509 18343
rect 16724 18312 17509 18340
rect 16724 18300 16730 18312
rect 17497 18309 17509 18312
rect 17543 18309 17555 18343
rect 17497 18303 17555 18309
rect 18049 18343 18107 18349
rect 18049 18309 18061 18343
rect 18095 18340 18107 18343
rect 18138 18340 18144 18352
rect 18095 18312 18144 18340
rect 18095 18309 18107 18312
rect 18049 18303 18107 18309
rect 18138 18300 18144 18312
rect 18196 18300 18202 18352
rect 20070 18340 20076 18352
rect 19274 18312 20076 18340
rect 20070 18300 20076 18312
rect 20128 18340 20134 18352
rect 20128 18312 20194 18340
rect 20128 18300 20134 18312
rect 21082 18300 21088 18352
rect 21140 18340 21146 18352
rect 21361 18343 21419 18349
rect 21361 18340 21373 18343
rect 21140 18312 21373 18340
rect 21140 18300 21146 18312
rect 21361 18309 21373 18312
rect 21407 18309 21419 18343
rect 21361 18303 21419 18309
rect 13725 18275 13783 18281
rect 13725 18241 13737 18275
rect 13771 18241 13783 18275
rect 13725 18235 13783 18241
rect 13909 18275 13967 18281
rect 13909 18241 13921 18275
rect 13955 18241 13967 18275
rect 13909 18235 13967 18241
rect 13354 18204 13360 18216
rect 12912 18176 13360 18204
rect 13354 18164 13360 18176
rect 13412 18204 13418 18216
rect 13924 18204 13952 18235
rect 16390 18232 16396 18284
rect 16448 18272 16454 18284
rect 16853 18275 16911 18281
rect 16853 18272 16865 18275
rect 16448 18244 16865 18272
rect 16448 18232 16454 18244
rect 16853 18241 16865 18244
rect 16899 18272 16911 18275
rect 17313 18275 17371 18281
rect 17313 18272 17325 18275
rect 16899 18244 17325 18272
rect 16899 18241 16911 18244
rect 16853 18235 16911 18241
rect 17313 18241 17325 18244
rect 17359 18241 17371 18275
rect 17313 18235 17371 18241
rect 22186 18232 22192 18284
rect 22244 18232 22250 18284
rect 13412 18176 13952 18204
rect 16209 18207 16267 18213
rect 13412 18164 13418 18176
rect 16209 18173 16221 18207
rect 16255 18204 16267 18207
rect 16298 18204 16304 18216
rect 16255 18176 16304 18204
rect 16255 18173 16267 18176
rect 16209 18167 16267 18173
rect 16298 18164 16304 18176
rect 16356 18204 16362 18216
rect 17773 18207 17831 18213
rect 17773 18204 17785 18207
rect 16356 18176 17785 18204
rect 16356 18164 16362 18176
rect 17773 18173 17785 18176
rect 17819 18173 17831 18207
rect 17773 18167 17831 18173
rect 19889 18207 19947 18213
rect 19889 18173 19901 18207
rect 19935 18204 19947 18207
rect 20162 18204 20168 18216
rect 19935 18176 20168 18204
rect 19935 18173 19947 18176
rect 19889 18167 19947 18173
rect 20162 18164 20168 18176
rect 20220 18164 20226 18216
rect 21634 18164 21640 18216
rect 21692 18164 21698 18216
rect 22278 18164 22284 18216
rect 22336 18164 22342 18216
rect 13725 18139 13783 18145
rect 13725 18136 13737 18139
rect 12406 18108 13737 18136
rect 13725 18105 13737 18108
rect 13771 18105 13783 18139
rect 13725 18099 13783 18105
rect 19058 18096 19064 18148
rect 19116 18136 19122 18148
rect 20254 18136 20260 18148
rect 19116 18108 20260 18136
rect 19116 18096 19122 18108
rect 20254 18096 20260 18108
rect 20312 18096 20318 18148
rect 3476 18040 3556 18068
rect 5169 18071 5227 18077
rect 3476 18028 3482 18040
rect 5169 18037 5181 18071
rect 5215 18068 5227 18071
rect 5258 18068 5264 18080
rect 5215 18040 5264 18068
rect 5215 18037 5227 18040
rect 5169 18031 5227 18037
rect 5258 18028 5264 18040
rect 5316 18028 5322 18080
rect 11885 18071 11943 18077
rect 11885 18037 11897 18071
rect 11931 18068 11943 18071
rect 12434 18068 12440 18080
rect 11931 18040 12440 18068
rect 11931 18037 11943 18040
rect 11885 18031 11943 18037
rect 12434 18028 12440 18040
rect 12492 18028 12498 18080
rect 12621 18071 12679 18077
rect 12621 18037 12633 18071
rect 12667 18068 12679 18071
rect 12710 18068 12716 18080
rect 12667 18040 12716 18068
rect 12667 18037 12679 18040
rect 12621 18031 12679 18037
rect 12710 18028 12716 18040
rect 12768 18028 12774 18080
rect 12805 18071 12863 18077
rect 12805 18037 12817 18071
rect 12851 18068 12863 18071
rect 12986 18068 12992 18080
rect 12851 18040 12992 18068
rect 12851 18037 12863 18040
rect 12805 18031 12863 18037
rect 12986 18028 12992 18040
rect 13044 18028 13050 18080
rect 17218 18028 17224 18080
rect 17276 18028 17282 18080
rect 17678 18028 17684 18080
rect 17736 18028 17742 18080
rect 19150 18028 19156 18080
rect 19208 18068 19214 18080
rect 20898 18068 20904 18080
rect 19208 18040 20904 18068
rect 19208 18028 19214 18040
rect 20898 18028 20904 18040
rect 20956 18068 20962 18080
rect 23382 18068 23388 18080
rect 20956 18040 23388 18068
rect 20956 18028 20962 18040
rect 23382 18028 23388 18040
rect 23440 18028 23446 18080
rect 1104 17978 25208 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 25208 17978
rect 1104 17904 25208 17926
rect 12066 17824 12072 17876
rect 12124 17864 12130 17876
rect 13170 17864 13176 17876
rect 12124 17836 13176 17864
rect 12124 17824 12130 17836
rect 13170 17824 13176 17836
rect 13228 17824 13234 17876
rect 13630 17824 13636 17876
rect 13688 17864 13694 17876
rect 13909 17867 13967 17873
rect 13909 17864 13921 17867
rect 13688 17836 13921 17864
rect 13688 17824 13694 17836
rect 13909 17833 13921 17836
rect 13955 17833 13967 17867
rect 13909 17827 13967 17833
rect 14734 17824 14740 17876
rect 14792 17864 14798 17876
rect 15562 17864 15568 17876
rect 14792 17836 15568 17864
rect 14792 17824 14798 17836
rect 15562 17824 15568 17836
rect 15620 17824 15626 17876
rect 16850 17824 16856 17876
rect 16908 17824 16914 17876
rect 18785 17867 18843 17873
rect 18785 17833 18797 17867
rect 18831 17864 18843 17867
rect 18874 17864 18880 17876
rect 18831 17836 18880 17864
rect 18831 17833 18843 17836
rect 18785 17827 18843 17833
rect 18874 17824 18880 17836
rect 18932 17824 18938 17876
rect 18966 17824 18972 17876
rect 19024 17824 19030 17876
rect 20806 17824 20812 17876
rect 20864 17864 20870 17876
rect 20993 17867 21051 17873
rect 20993 17864 21005 17867
rect 20864 17836 21005 17864
rect 20864 17824 20870 17836
rect 20993 17833 21005 17836
rect 21039 17833 21051 17867
rect 20993 17827 21051 17833
rect 16669 17799 16727 17805
rect 16669 17765 16681 17799
rect 16715 17796 16727 17799
rect 17034 17796 17040 17808
rect 16715 17768 17040 17796
rect 16715 17765 16727 17768
rect 16669 17759 16727 17765
rect 17034 17756 17040 17768
rect 17092 17796 17098 17808
rect 17402 17796 17408 17808
rect 17092 17768 17408 17796
rect 17092 17756 17098 17768
rect 17402 17756 17408 17768
rect 17460 17756 17466 17808
rect 1394 17688 1400 17740
rect 1452 17728 1458 17740
rect 2682 17728 2688 17740
rect 1452 17700 2688 17728
rect 1452 17688 1458 17700
rect 2682 17688 2688 17700
rect 2740 17688 2746 17740
rect 10594 17688 10600 17740
rect 10652 17688 10658 17740
rect 12161 17731 12219 17737
rect 12161 17697 12173 17731
rect 12207 17728 12219 17731
rect 13906 17728 13912 17740
rect 12207 17700 13912 17728
rect 12207 17697 12219 17700
rect 12161 17691 12219 17697
rect 13906 17688 13912 17700
rect 13964 17728 13970 17740
rect 16298 17728 16304 17740
rect 13964 17700 16304 17728
rect 13964 17688 13970 17700
rect 16298 17688 16304 17700
rect 16356 17688 16362 17740
rect 18414 17688 18420 17740
rect 18472 17728 18478 17740
rect 19245 17731 19303 17737
rect 19245 17728 19257 17731
rect 18472 17700 19257 17728
rect 18472 17688 18478 17700
rect 19245 17697 19257 17700
rect 19291 17728 19303 17731
rect 21634 17728 21640 17740
rect 19291 17700 21640 17728
rect 19291 17697 19303 17700
rect 19245 17691 19303 17697
rect 21634 17688 21640 17700
rect 21692 17728 21698 17740
rect 22002 17728 22008 17740
rect 21692 17700 22008 17728
rect 21692 17688 21698 17700
rect 22002 17688 22008 17700
rect 22060 17688 22066 17740
rect 1765 17663 1823 17669
rect 1765 17629 1777 17663
rect 1811 17660 1823 17663
rect 1854 17660 1860 17672
rect 1811 17632 1860 17660
rect 1811 17629 1823 17632
rect 1765 17623 1823 17629
rect 1854 17620 1860 17632
rect 1912 17620 1918 17672
rect 3191 17663 3249 17669
rect 3191 17629 3203 17663
rect 3237 17660 3249 17663
rect 3789 17663 3847 17669
rect 3789 17660 3801 17663
rect 3237 17632 3801 17660
rect 3237 17629 3249 17632
rect 3191 17623 3249 17629
rect 3789 17629 3801 17632
rect 3835 17629 3847 17663
rect 3789 17623 3847 17629
rect 9582 17620 9588 17672
rect 9640 17660 9646 17672
rect 10321 17663 10379 17669
rect 10321 17660 10333 17663
rect 9640 17632 10333 17660
rect 9640 17620 9646 17632
rect 10321 17629 10333 17632
rect 10367 17629 10379 17663
rect 10321 17623 10379 17629
rect 17218 17620 17224 17672
rect 17276 17620 17282 17672
rect 17954 17620 17960 17672
rect 18012 17660 18018 17672
rect 18601 17663 18659 17669
rect 18601 17660 18613 17663
rect 18012 17632 18613 17660
rect 18012 17620 18018 17632
rect 18601 17629 18613 17632
rect 18647 17660 18659 17663
rect 18877 17663 18935 17669
rect 18877 17660 18889 17663
rect 18647 17632 18889 17660
rect 18647 17629 18659 17632
rect 18601 17623 18659 17629
rect 18877 17629 18889 17632
rect 18923 17629 18935 17663
rect 18877 17623 18935 17629
rect 19058 17620 19064 17672
rect 19116 17620 19122 17672
rect 3326 17592 3332 17604
rect 2806 17564 3332 17592
rect 3326 17552 3332 17564
rect 3384 17552 3390 17604
rect 11330 17552 11336 17604
rect 11388 17552 11394 17604
rect 12437 17595 12495 17601
rect 12437 17561 12449 17595
rect 12483 17592 12495 17595
rect 12710 17592 12716 17604
rect 12483 17564 12716 17592
rect 12483 17561 12495 17564
rect 12437 17555 12495 17561
rect 12710 17552 12716 17564
rect 12768 17552 12774 17604
rect 13998 17592 14004 17604
rect 13662 17564 14004 17592
rect 13998 17552 14004 17564
rect 14056 17592 14062 17604
rect 14734 17592 14740 17604
rect 14056 17564 14740 17592
rect 14056 17552 14062 17564
rect 14734 17552 14740 17564
rect 14792 17552 14798 17604
rect 15562 17552 15568 17604
rect 15620 17592 15626 17604
rect 16025 17595 16083 17601
rect 15620 17564 15700 17592
rect 15620 17552 15626 17564
rect 4154 17484 4160 17536
rect 4212 17524 4218 17536
rect 4433 17527 4491 17533
rect 4433 17524 4445 17527
rect 4212 17496 4445 17524
rect 4212 17484 4218 17496
rect 4433 17493 4445 17496
rect 4479 17493 4491 17527
rect 4433 17487 4491 17493
rect 14553 17527 14611 17533
rect 14553 17493 14565 17527
rect 14599 17524 14611 17527
rect 15194 17524 15200 17536
rect 14599 17496 15200 17524
rect 14599 17493 14611 17496
rect 14553 17487 14611 17493
rect 15194 17484 15200 17496
rect 15252 17484 15258 17536
rect 15672 17524 15700 17564
rect 16025 17561 16037 17595
rect 16071 17592 16083 17595
rect 16114 17592 16120 17604
rect 16071 17564 16120 17592
rect 16071 17561 16083 17564
rect 16025 17555 16083 17561
rect 16114 17552 16120 17564
rect 16172 17552 16178 17604
rect 16574 17592 16580 17604
rect 16224 17564 16580 17592
rect 16224 17524 16252 17564
rect 16574 17552 16580 17564
rect 16632 17552 16638 17604
rect 17236 17592 17264 17620
rect 18417 17595 18475 17601
rect 18417 17592 18429 17595
rect 17236 17564 18429 17592
rect 18417 17561 18429 17564
rect 18463 17561 18475 17595
rect 18417 17555 18475 17561
rect 15672 17496 16252 17524
rect 16390 17484 16396 17536
rect 16448 17524 16454 17536
rect 16853 17527 16911 17533
rect 16853 17524 16865 17527
rect 16448 17496 16865 17524
rect 16448 17484 16454 17496
rect 16853 17493 16865 17496
rect 16899 17524 16911 17527
rect 18322 17524 18328 17536
rect 16899 17496 18328 17524
rect 16899 17493 16911 17496
rect 16853 17487 16911 17493
rect 18322 17484 18328 17496
rect 18380 17484 18386 17536
rect 18432 17524 18460 17555
rect 19076 17524 19104 17620
rect 19518 17552 19524 17604
rect 19576 17552 19582 17604
rect 20070 17552 20076 17604
rect 20128 17552 20134 17604
rect 18432 17496 19104 17524
rect 1104 17434 25208 17456
rect 1104 17382 4874 17434
rect 4926 17382 4938 17434
rect 4990 17382 5002 17434
rect 5054 17382 5066 17434
rect 5118 17382 5130 17434
rect 5182 17382 25208 17434
rect 1104 17360 25208 17382
rect 2225 17323 2283 17329
rect 2225 17289 2237 17323
rect 2271 17320 2283 17323
rect 2866 17320 2872 17332
rect 2271 17292 2872 17320
rect 2271 17289 2283 17292
rect 2225 17283 2283 17289
rect 2866 17280 2872 17292
rect 2924 17280 2930 17332
rect 3418 17320 3424 17332
rect 3068 17292 3424 17320
rect 2731 17255 2789 17261
rect 2731 17221 2743 17255
rect 2777 17252 2789 17255
rect 3068 17252 3096 17292
rect 3418 17280 3424 17292
rect 3476 17280 3482 17332
rect 11146 17280 11152 17332
rect 11204 17320 11210 17332
rect 11333 17323 11391 17329
rect 11333 17320 11345 17323
rect 11204 17292 11345 17320
rect 11204 17280 11210 17292
rect 11333 17289 11345 17292
rect 11379 17289 11391 17323
rect 11333 17283 11391 17289
rect 15825 17323 15883 17329
rect 15825 17289 15837 17323
rect 15871 17320 15883 17323
rect 17678 17320 17684 17332
rect 15871 17292 17684 17320
rect 15871 17289 15883 17292
rect 15825 17283 15883 17289
rect 17678 17280 17684 17292
rect 17736 17280 17742 17332
rect 18046 17280 18052 17332
rect 18104 17320 18110 17332
rect 18509 17323 18567 17329
rect 18509 17320 18521 17323
rect 18104 17292 18521 17320
rect 18104 17280 18110 17292
rect 18509 17289 18521 17292
rect 18555 17289 18567 17323
rect 18509 17283 18567 17289
rect 18693 17323 18751 17329
rect 18693 17289 18705 17323
rect 18739 17320 18751 17323
rect 19150 17320 19156 17332
rect 18739 17292 19156 17320
rect 18739 17289 18751 17292
rect 18693 17283 18751 17289
rect 2777 17224 3096 17252
rect 2777 17221 2789 17224
rect 2731 17215 2789 17221
rect 3326 17212 3332 17264
rect 3384 17212 3390 17264
rect 9858 17212 9864 17264
rect 9916 17212 9922 17264
rect 15930 17212 15936 17264
rect 15988 17252 15994 17264
rect 16025 17255 16083 17261
rect 16025 17252 16037 17255
rect 15988 17224 16037 17252
rect 15988 17212 15994 17224
rect 16025 17221 16037 17224
rect 16071 17252 16083 17255
rect 16390 17252 16396 17264
rect 16071 17224 16396 17252
rect 16071 17221 16083 17224
rect 16025 17215 16083 17221
rect 16390 17212 16396 17224
rect 16448 17212 16454 17264
rect 17034 17212 17040 17264
rect 17092 17212 17098 17264
rect 17494 17212 17500 17264
rect 17552 17212 17558 17264
rect 18322 17212 18328 17264
rect 18380 17252 18386 17264
rect 18708 17252 18736 17283
rect 19150 17280 19156 17292
rect 19208 17280 19214 17332
rect 18380 17224 18736 17252
rect 18380 17212 18386 17224
rect 4154 17144 4160 17196
rect 4212 17144 4218 17196
rect 4525 17187 4583 17193
rect 4525 17153 4537 17187
rect 4571 17184 4583 17187
rect 4614 17184 4620 17196
rect 4571 17156 4620 17184
rect 4571 17153 4583 17156
rect 4525 17147 4583 17153
rect 4614 17144 4620 17156
rect 4672 17144 4678 17196
rect 8662 17144 8668 17196
rect 8720 17184 8726 17196
rect 9582 17184 9588 17196
rect 8720 17156 9588 17184
rect 8720 17144 8726 17156
rect 9582 17144 9588 17156
rect 9640 17144 9646 17196
rect 11330 17184 11336 17196
rect 10994 17156 11336 17184
rect 11330 17144 11336 17156
rect 11388 17144 11394 17196
rect 16298 17144 16304 17196
rect 16356 17184 16362 17196
rect 16761 17187 16819 17193
rect 16761 17184 16773 17187
rect 16356 17156 16773 17184
rect 16356 17144 16362 17156
rect 16761 17153 16773 17156
rect 16807 17153 16819 17187
rect 16761 17147 16819 17153
rect 18877 17187 18935 17193
rect 18877 17153 18889 17187
rect 18923 17184 18935 17187
rect 19426 17184 19432 17196
rect 18923 17156 19432 17184
rect 18923 17153 18935 17156
rect 18877 17147 18935 17153
rect 19426 17144 19432 17156
rect 19484 17144 19490 17196
rect 1854 17076 1860 17128
rect 1912 17116 1918 17128
rect 2317 17119 2375 17125
rect 2317 17116 2329 17119
rect 1912 17088 2329 17116
rect 1912 17076 1918 17088
rect 2317 17085 2329 17088
rect 2363 17085 2375 17119
rect 2317 17079 2375 17085
rect 2501 17119 2559 17125
rect 2501 17085 2513 17119
rect 2547 17116 2559 17119
rect 2958 17116 2964 17128
rect 2547 17088 2964 17116
rect 2547 17085 2559 17088
rect 2501 17079 2559 17085
rect 2958 17076 2964 17088
rect 3016 17116 3022 17128
rect 3418 17116 3424 17128
rect 3016 17088 3424 17116
rect 3016 17076 3022 17088
rect 3418 17076 3424 17088
rect 3476 17076 3482 17128
rect 16574 17076 16580 17128
rect 16632 17116 16638 17128
rect 17494 17116 17500 17128
rect 16632 17088 17500 17116
rect 16632 17076 16638 17088
rect 17494 17076 17500 17088
rect 17552 17076 17558 17128
rect 15657 17051 15715 17057
rect 15657 17017 15669 17051
rect 15703 17048 15715 17051
rect 16114 17048 16120 17060
rect 15703 17020 16120 17048
rect 15703 17017 15715 17020
rect 15657 17011 15715 17017
rect 16114 17008 16120 17020
rect 16172 17008 16178 17060
rect 1762 16940 1768 16992
rect 1820 16980 1826 16992
rect 1857 16983 1915 16989
rect 1857 16980 1869 16983
rect 1820 16952 1869 16980
rect 1820 16940 1826 16952
rect 1857 16949 1869 16952
rect 1903 16949 1915 16983
rect 1857 16943 1915 16949
rect 15841 16983 15899 16989
rect 15841 16949 15853 16983
rect 15887 16980 15899 16983
rect 16206 16980 16212 16992
rect 15887 16952 16212 16980
rect 15887 16949 15899 16952
rect 15841 16943 15899 16949
rect 16206 16940 16212 16952
rect 16264 16940 16270 16992
rect 1104 16890 25208 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 25208 16890
rect 1104 16816 25208 16838
rect 2866 16736 2872 16788
rect 2924 16776 2930 16788
rect 3191 16779 3249 16785
rect 3191 16776 3203 16779
rect 2924 16748 3203 16776
rect 2924 16736 2930 16748
rect 3191 16745 3203 16748
rect 3237 16745 3249 16779
rect 3191 16739 3249 16745
rect 8846 16736 8852 16788
rect 8904 16776 8910 16788
rect 9217 16779 9275 16785
rect 9217 16776 9229 16779
rect 8904 16748 9229 16776
rect 8904 16736 8910 16748
rect 9217 16745 9229 16748
rect 9263 16776 9275 16779
rect 10042 16776 10048 16788
rect 9263 16748 10048 16776
rect 9263 16745 9275 16748
rect 9217 16739 9275 16745
rect 10042 16736 10048 16748
rect 10100 16736 10106 16788
rect 21082 16668 21088 16720
rect 21140 16708 21146 16720
rect 22281 16711 22339 16717
rect 22281 16708 22293 16711
rect 21140 16680 22293 16708
rect 21140 16668 21146 16680
rect 22281 16677 22293 16680
rect 22327 16677 22339 16711
rect 22281 16671 22339 16677
rect 1394 16600 1400 16652
rect 1452 16600 1458 16652
rect 1762 16600 1768 16652
rect 1820 16600 1826 16652
rect 4614 16600 4620 16652
rect 4672 16640 4678 16652
rect 5353 16643 5411 16649
rect 5353 16640 5365 16643
rect 4672 16612 5365 16640
rect 4672 16600 4678 16612
rect 5353 16609 5365 16612
rect 5399 16609 5411 16643
rect 5353 16603 5411 16609
rect 6914 16600 6920 16652
rect 6972 16640 6978 16652
rect 7147 16643 7205 16649
rect 7147 16640 7159 16643
rect 6972 16612 7159 16640
rect 6972 16600 6978 16612
rect 7147 16609 7159 16612
rect 7193 16640 7205 16643
rect 8113 16643 8171 16649
rect 8113 16640 8125 16643
rect 7193 16612 8125 16640
rect 7193 16609 7205 16612
rect 7147 16603 7205 16609
rect 8113 16609 8125 16612
rect 8159 16609 8171 16643
rect 8113 16603 8171 16609
rect 8202 16600 8208 16652
rect 8260 16600 8266 16652
rect 22189 16643 22247 16649
rect 22189 16609 22201 16643
rect 22235 16640 22247 16643
rect 22373 16643 22431 16649
rect 22235 16612 22324 16640
rect 22235 16609 22247 16612
rect 22189 16603 22247 16609
rect 22296 16584 22324 16612
rect 22373 16609 22385 16643
rect 22419 16640 22431 16643
rect 22922 16640 22928 16652
rect 22419 16612 22928 16640
rect 22419 16609 22431 16612
rect 22373 16603 22431 16609
rect 22922 16600 22928 16612
rect 22980 16600 22986 16652
rect 5718 16532 5724 16584
rect 5776 16532 5782 16584
rect 22278 16532 22284 16584
rect 22336 16532 22342 16584
rect 22465 16575 22523 16581
rect 22465 16541 22477 16575
rect 22511 16541 22523 16575
rect 22465 16535 22523 16541
rect 3326 16504 3332 16516
rect 2806 16476 3332 16504
rect 3326 16464 3332 16476
rect 3384 16464 3390 16516
rect 6086 16464 6092 16516
rect 6144 16464 6150 16516
rect 9306 16464 9312 16516
rect 9364 16464 9370 16516
rect 20070 16464 20076 16516
rect 20128 16504 20134 16516
rect 21634 16504 21640 16516
rect 20128 16476 21640 16504
rect 20128 16464 20134 16476
rect 21634 16464 21640 16476
rect 21692 16504 21698 16516
rect 21692 16476 22094 16504
rect 21692 16464 21698 16476
rect 7653 16439 7711 16445
rect 7653 16405 7665 16439
rect 7699 16436 7711 16439
rect 7834 16436 7840 16448
rect 7699 16408 7840 16436
rect 7699 16405 7711 16408
rect 7653 16399 7711 16405
rect 7834 16396 7840 16408
rect 7892 16396 7898 16448
rect 8021 16439 8079 16445
rect 8021 16405 8033 16439
rect 8067 16436 8079 16439
rect 9030 16436 9036 16448
rect 8067 16408 9036 16436
rect 8067 16405 8079 16408
rect 8021 16399 8079 16405
rect 9030 16396 9036 16408
rect 9088 16396 9094 16448
rect 22066 16436 22094 16476
rect 22186 16464 22192 16516
rect 22244 16504 22250 16516
rect 22480 16504 22508 16535
rect 22244 16476 22508 16504
rect 22244 16464 22250 16476
rect 23198 16436 23204 16448
rect 22066 16408 23204 16436
rect 23198 16396 23204 16408
rect 23256 16396 23262 16448
rect 1104 16346 25208 16368
rect 1104 16294 4874 16346
rect 4926 16294 4938 16346
rect 4990 16294 5002 16346
rect 5054 16294 5066 16346
rect 5118 16294 5130 16346
rect 5182 16294 25208 16346
rect 1104 16272 25208 16294
rect 5718 16192 5724 16244
rect 5776 16232 5782 16244
rect 6365 16235 6423 16241
rect 6365 16232 6377 16235
rect 5776 16204 6377 16232
rect 5776 16192 5782 16204
rect 6365 16201 6377 16204
rect 6411 16201 6423 16235
rect 6365 16195 6423 16201
rect 6733 16235 6791 16241
rect 6733 16201 6745 16235
rect 6779 16232 6791 16235
rect 6914 16232 6920 16244
rect 6779 16204 6920 16232
rect 6779 16201 6791 16204
rect 6733 16195 6791 16201
rect 6914 16192 6920 16204
rect 6972 16192 6978 16244
rect 8662 16232 8668 16244
rect 7484 16204 8668 16232
rect 2777 16167 2835 16173
rect 2777 16133 2789 16167
rect 2823 16164 2835 16167
rect 2866 16164 2872 16176
rect 2823 16136 2872 16164
rect 2823 16133 2835 16136
rect 2777 16127 2835 16133
rect 2866 16124 2872 16136
rect 2924 16124 2930 16176
rect 5813 16099 5871 16105
rect 5813 16065 5825 16099
rect 5859 16096 5871 16099
rect 6822 16096 6828 16108
rect 5859 16068 6828 16096
rect 5859 16065 5871 16068
rect 5813 16059 5871 16065
rect 6822 16056 6828 16068
rect 6880 16056 6886 16108
rect 7484 16105 7512 16204
rect 8662 16192 8668 16204
rect 8720 16192 8726 16244
rect 13909 16235 13967 16241
rect 13909 16201 13921 16235
rect 13955 16232 13967 16235
rect 14277 16235 14335 16241
rect 13955 16204 14228 16232
rect 13955 16201 13967 16204
rect 13909 16195 13967 16201
rect 8846 16124 8852 16176
rect 8904 16124 8910 16176
rect 9030 16124 9036 16176
rect 9088 16164 9094 16176
rect 9263 16167 9321 16173
rect 9263 16164 9275 16167
rect 9088 16136 9275 16164
rect 9088 16124 9094 16136
rect 9263 16133 9275 16136
rect 9309 16164 9321 16167
rect 10505 16167 10563 16173
rect 10505 16164 10517 16167
rect 9309 16136 10517 16164
rect 9309 16133 9321 16136
rect 9263 16127 9321 16133
rect 10505 16133 10517 16136
rect 10551 16164 10563 16167
rect 11974 16164 11980 16176
rect 10551 16136 11980 16164
rect 10551 16133 10563 16136
rect 10505 16127 10563 16133
rect 11974 16124 11980 16136
rect 12032 16124 12038 16176
rect 7469 16099 7527 16105
rect 7469 16065 7481 16099
rect 7515 16065 7527 16099
rect 7469 16059 7527 16065
rect 7834 16056 7840 16108
rect 7892 16056 7898 16108
rect 10413 16099 10471 16105
rect 10413 16065 10425 16099
rect 10459 16096 10471 16099
rect 12250 16096 12256 16108
rect 10459 16068 12256 16096
rect 10459 16065 10471 16068
rect 10413 16059 10471 16065
rect 12250 16056 12256 16068
rect 12308 16056 12314 16108
rect 13541 16099 13599 16105
rect 13541 16065 13553 16099
rect 13587 16065 13599 16099
rect 13541 16059 13599 16065
rect 2774 15988 2780 16040
rect 2832 16028 2838 16040
rect 2869 16031 2927 16037
rect 2869 16028 2881 16031
rect 2832 16000 2881 16028
rect 2832 15988 2838 16000
rect 2869 15997 2881 16000
rect 2915 15997 2927 16031
rect 2869 15991 2927 15997
rect 2958 15988 2964 16040
rect 3016 16028 3022 16040
rect 3142 16028 3148 16040
rect 3016 16000 3148 16028
rect 3016 15988 3022 16000
rect 3142 15988 3148 16000
rect 3200 15988 3206 16040
rect 5902 15988 5908 16040
rect 5960 15988 5966 16040
rect 5994 15988 6000 16040
rect 6052 16028 6058 16040
rect 6917 16031 6975 16037
rect 6917 16028 6929 16031
rect 6052 16000 6929 16028
rect 6052 15988 6058 16000
rect 6917 15997 6929 16000
rect 6963 15997 6975 16031
rect 6917 15991 6975 15997
rect 10594 15988 10600 16040
rect 10652 15988 10658 16040
rect 13556 15960 13584 16059
rect 13722 16056 13728 16108
rect 13780 16096 13786 16108
rect 14001 16099 14059 16105
rect 14001 16096 14013 16099
rect 13780 16068 14013 16096
rect 13780 16056 13786 16068
rect 14001 16065 14013 16068
rect 14047 16065 14059 16099
rect 14001 16059 14059 16065
rect 13633 16031 13691 16037
rect 13633 15997 13645 16031
rect 13679 16028 13691 16031
rect 14090 16028 14096 16040
rect 13679 16000 14096 16028
rect 13679 15997 13691 16000
rect 13633 15991 13691 15997
rect 14090 15988 14096 16000
rect 14148 15988 14154 16040
rect 14200 15960 14228 16204
rect 14277 16201 14289 16235
rect 14323 16232 14335 16235
rect 14323 16204 15056 16232
rect 14323 16201 14335 16204
rect 14277 16195 14335 16201
rect 15028 16105 15056 16204
rect 20070 16164 20076 16176
rect 19918 16136 20076 16164
rect 20070 16124 20076 16136
rect 20128 16124 20134 16176
rect 20916 16136 21956 16164
rect 15013 16099 15071 16105
rect 15013 16065 15025 16099
rect 15059 16096 15071 16099
rect 15470 16096 15476 16108
rect 15059 16068 15476 16096
rect 15059 16065 15071 16068
rect 15013 16059 15071 16065
rect 15470 16056 15476 16068
rect 15528 16056 15534 16108
rect 15654 16056 15660 16108
rect 15712 16056 15718 16108
rect 18414 16056 18420 16108
rect 18472 16056 18478 16108
rect 20916 16105 20944 16136
rect 21192 16105 21220 16136
rect 20717 16099 20775 16105
rect 20717 16065 20729 16099
rect 20763 16065 20775 16099
rect 20717 16059 20775 16065
rect 20901 16099 20959 16105
rect 20901 16065 20913 16099
rect 20947 16065 20959 16099
rect 20901 16059 20959 16065
rect 20993 16099 21051 16105
rect 20993 16065 21005 16099
rect 21039 16065 21051 16099
rect 20993 16059 21051 16065
rect 21177 16099 21235 16105
rect 21177 16065 21189 16099
rect 21223 16065 21235 16099
rect 21177 16059 21235 16065
rect 14274 15988 14280 16040
rect 14332 15988 14338 16040
rect 14734 15988 14740 16040
rect 14792 15988 14798 16040
rect 14826 15988 14832 16040
rect 14884 15988 14890 16040
rect 14921 16031 14979 16037
rect 14921 15997 14933 16031
rect 14967 15997 14979 16031
rect 14921 15991 14979 15997
rect 14936 15960 14964 15991
rect 15378 15988 15384 16040
rect 15436 16028 15442 16040
rect 15565 16031 15623 16037
rect 15565 16028 15577 16031
rect 15436 16000 15577 16028
rect 15436 15988 15442 16000
rect 15565 15997 15577 16000
rect 15611 15997 15623 16031
rect 15565 15991 15623 15997
rect 18693 16031 18751 16037
rect 18693 15997 18705 16031
rect 18739 16028 18751 16031
rect 19886 16028 19892 16040
rect 18739 16000 19892 16028
rect 18739 15997 18751 16000
rect 18693 15991 18751 15997
rect 19886 15988 19892 16000
rect 19944 15988 19950 16040
rect 20165 16031 20223 16037
rect 20165 15997 20177 16031
rect 20211 16028 20223 16031
rect 20732 16028 20760 16059
rect 20211 16000 20760 16028
rect 20211 15997 20223 16000
rect 20165 15991 20223 15997
rect 20806 15988 20812 16040
rect 20864 16028 20870 16040
rect 21008 16028 21036 16059
rect 21358 16056 21364 16108
rect 21416 16056 21422 16108
rect 20864 16000 21036 16028
rect 21637 16031 21695 16037
rect 20864 15988 20870 16000
rect 21637 15997 21649 16031
rect 21683 16028 21695 16031
rect 21821 16031 21879 16037
rect 21821 16028 21833 16031
rect 21683 16000 21833 16028
rect 21683 15997 21695 16000
rect 21637 15991 21695 15997
rect 21821 15997 21833 16000
rect 21867 15997 21879 16031
rect 21928 16028 21956 16136
rect 23198 16124 23204 16176
rect 23256 16164 23262 16176
rect 23382 16164 23388 16176
rect 23256 16136 23388 16164
rect 23256 16124 23262 16136
rect 23382 16124 23388 16136
rect 23440 16164 23446 16176
rect 23440 16136 23598 16164
rect 23440 16124 23446 16136
rect 22094 16056 22100 16108
rect 22152 16096 22158 16108
rect 22833 16099 22891 16105
rect 22833 16096 22845 16099
rect 22152 16068 22845 16096
rect 22152 16056 22158 16068
rect 22833 16065 22845 16068
rect 22879 16065 22891 16099
rect 22833 16059 22891 16065
rect 22373 16031 22431 16037
rect 22373 16028 22385 16031
rect 21928 16000 22385 16028
rect 21821 15991 21879 15997
rect 22373 15997 22385 16000
rect 22419 16028 22431 16031
rect 22646 16028 22652 16040
rect 22419 16000 22652 16028
rect 22419 15997 22431 16000
rect 22373 15991 22431 15997
rect 22646 15988 22652 16000
rect 22704 15988 22710 16040
rect 23106 15988 23112 16040
rect 23164 15988 23170 16040
rect 13556 15932 14136 15960
rect 14200 15932 14964 15960
rect 14108 15904 14136 15932
rect 2038 15852 2044 15904
rect 2096 15892 2102 15904
rect 2409 15895 2467 15901
rect 2409 15892 2421 15895
rect 2096 15864 2421 15892
rect 2096 15852 2102 15864
rect 2409 15861 2421 15864
rect 2455 15861 2467 15895
rect 2409 15855 2467 15861
rect 5350 15852 5356 15904
rect 5408 15892 5414 15904
rect 5445 15895 5503 15901
rect 5445 15892 5457 15895
rect 5408 15864 5457 15892
rect 5408 15852 5414 15864
rect 5445 15861 5457 15864
rect 5491 15861 5503 15895
rect 5445 15855 5503 15861
rect 10045 15895 10103 15901
rect 10045 15861 10057 15895
rect 10091 15892 10103 15895
rect 10134 15892 10140 15904
rect 10091 15864 10140 15892
rect 10091 15861 10103 15864
rect 10045 15855 10103 15861
rect 10134 15852 10140 15864
rect 10192 15852 10198 15904
rect 12802 15852 12808 15904
rect 12860 15892 12866 15904
rect 13541 15895 13599 15901
rect 13541 15892 13553 15895
rect 12860 15864 13553 15892
rect 12860 15852 12866 15864
rect 13541 15861 13553 15864
rect 13587 15892 13599 15895
rect 13722 15892 13728 15904
rect 13587 15864 13728 15892
rect 13587 15861 13599 15864
rect 13541 15855 13599 15861
rect 13722 15852 13728 15864
rect 13780 15852 13786 15904
rect 14090 15852 14096 15904
rect 14148 15852 14154 15904
rect 14936 15892 14964 15932
rect 15197 15963 15255 15969
rect 15197 15929 15209 15963
rect 15243 15960 15255 15963
rect 16022 15960 16028 15972
rect 15243 15932 16028 15960
rect 15243 15929 15255 15932
rect 15197 15923 15255 15929
rect 16022 15920 16028 15932
rect 16080 15920 16086 15972
rect 20346 15920 20352 15972
rect 20404 15960 20410 15972
rect 20993 15963 21051 15969
rect 20993 15960 21005 15963
rect 20404 15932 21005 15960
rect 20404 15920 20410 15932
rect 20993 15929 21005 15932
rect 21039 15929 21051 15963
rect 20993 15923 21051 15929
rect 21453 15963 21511 15969
rect 21453 15929 21465 15963
rect 21499 15960 21511 15963
rect 22278 15960 22284 15972
rect 21499 15932 22284 15960
rect 21499 15929 21511 15932
rect 21453 15923 21511 15929
rect 22278 15920 22284 15932
rect 22336 15920 22342 15972
rect 15562 15892 15568 15904
rect 14936 15864 15568 15892
rect 15562 15852 15568 15864
rect 15620 15852 15626 15904
rect 15933 15895 15991 15901
rect 15933 15861 15945 15895
rect 15979 15892 15991 15895
rect 17770 15892 17776 15904
rect 15979 15864 17776 15892
rect 15979 15861 15991 15864
rect 15933 15855 15991 15861
rect 17770 15852 17776 15864
rect 17828 15852 17834 15904
rect 20622 15852 20628 15904
rect 20680 15892 20686 15904
rect 20901 15895 20959 15901
rect 20901 15892 20913 15895
rect 20680 15864 20913 15892
rect 20680 15852 20686 15864
rect 20901 15861 20913 15864
rect 20947 15861 20959 15895
rect 20901 15855 20959 15861
rect 21174 15852 21180 15904
rect 21232 15892 21238 15904
rect 21361 15895 21419 15901
rect 21361 15892 21373 15895
rect 21232 15864 21373 15892
rect 21232 15852 21238 15864
rect 21361 15861 21373 15864
rect 21407 15861 21419 15895
rect 21361 15855 21419 15861
rect 22002 15852 22008 15904
rect 22060 15892 22066 15904
rect 23198 15892 23204 15904
rect 22060 15864 23204 15892
rect 22060 15852 22066 15864
rect 23198 15852 23204 15864
rect 23256 15852 23262 15904
rect 23290 15852 23296 15904
rect 23348 15892 23354 15904
rect 24581 15895 24639 15901
rect 24581 15892 24593 15895
rect 23348 15864 24593 15892
rect 23348 15852 23354 15864
rect 24581 15861 24593 15864
rect 24627 15861 24639 15895
rect 24581 15855 24639 15861
rect 1104 15802 25208 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 25208 15802
rect 1104 15728 25208 15750
rect 6086 15648 6092 15700
rect 6144 15688 6150 15700
rect 7101 15691 7159 15697
rect 7101 15688 7113 15691
rect 6144 15660 7113 15688
rect 6144 15648 6150 15660
rect 7101 15657 7113 15660
rect 7147 15657 7159 15691
rect 7101 15651 7159 15657
rect 7742 15648 7748 15700
rect 7800 15688 7806 15700
rect 8202 15688 8208 15700
rect 7800 15660 8208 15688
rect 7800 15648 7806 15660
rect 8202 15648 8208 15660
rect 8260 15688 8266 15700
rect 10594 15688 10600 15700
rect 8260 15660 8340 15688
rect 8260 15648 8266 15660
rect 1394 15580 1400 15632
rect 1452 15620 1458 15632
rect 4706 15620 4712 15632
rect 1452 15592 1716 15620
rect 1452 15580 1458 15592
rect 1688 15561 1716 15592
rect 4448 15592 4712 15620
rect 1673 15555 1731 15561
rect 1673 15521 1685 15555
rect 1719 15552 1731 15555
rect 2590 15552 2596 15564
rect 1719 15524 2596 15552
rect 1719 15521 1731 15524
rect 1673 15515 1731 15521
rect 2590 15512 2596 15524
rect 2648 15512 2654 15564
rect 4448 15561 4476 15592
rect 4706 15580 4712 15592
rect 4764 15580 4770 15632
rect 4433 15555 4491 15561
rect 4433 15521 4445 15555
rect 4479 15521 4491 15555
rect 4433 15515 4491 15521
rect 4614 15512 4620 15564
rect 4672 15552 4678 15564
rect 4985 15555 5043 15561
rect 4985 15552 4997 15555
rect 4672 15524 4997 15552
rect 4672 15512 4678 15524
rect 4985 15521 4997 15524
rect 5031 15521 5043 15555
rect 4985 15515 5043 15521
rect 5350 15512 5356 15564
rect 5408 15512 5414 15564
rect 6822 15561 6828 15564
rect 6779 15555 6828 15561
rect 6779 15552 6791 15555
rect 6735 15524 6791 15552
rect 6779 15521 6791 15524
rect 6825 15521 6828 15555
rect 6779 15515 6828 15521
rect 6822 15512 6828 15515
rect 6880 15552 6886 15564
rect 8312 15561 8340 15660
rect 9140 15660 10600 15688
rect 9140 15561 9168 15660
rect 10594 15648 10600 15660
rect 10652 15648 10658 15700
rect 13173 15691 13231 15697
rect 13173 15657 13185 15691
rect 13219 15688 13231 15691
rect 14826 15688 14832 15700
rect 13219 15660 14832 15688
rect 13219 15657 13231 15660
rect 13173 15651 13231 15657
rect 14826 15648 14832 15660
rect 14884 15688 14890 15700
rect 14884 15660 15884 15688
rect 14884 15648 14890 15660
rect 12434 15580 12440 15632
rect 12492 15620 12498 15632
rect 13722 15620 13728 15632
rect 12492 15592 13728 15620
rect 12492 15580 12498 15592
rect 13722 15580 13728 15592
rect 13780 15580 13786 15632
rect 14090 15580 14096 15632
rect 14148 15580 14154 15632
rect 15378 15580 15384 15632
rect 15436 15580 15442 15632
rect 15746 15580 15752 15632
rect 15804 15580 15810 15632
rect 8113 15555 8171 15561
rect 8113 15552 8125 15555
rect 6880 15524 8125 15552
rect 6880 15512 6886 15524
rect 8113 15521 8125 15524
rect 8159 15521 8171 15555
rect 8113 15515 8171 15521
rect 8297 15555 8355 15561
rect 8297 15521 8309 15555
rect 8343 15521 8355 15555
rect 8297 15515 8355 15521
rect 9125 15555 9183 15561
rect 9125 15521 9137 15555
rect 9171 15521 9183 15555
rect 9125 15515 9183 15521
rect 9582 15512 9588 15564
rect 9640 15552 9646 15564
rect 9769 15555 9827 15561
rect 9769 15552 9781 15555
rect 9640 15524 9781 15552
rect 9640 15512 9646 15524
rect 9769 15521 9781 15524
rect 9815 15521 9827 15555
rect 9769 15515 9827 15521
rect 10134 15512 10140 15564
rect 10192 15512 10198 15564
rect 10244 15524 11008 15552
rect 1394 15444 1400 15496
rect 1452 15444 1458 15496
rect 2038 15444 2044 15496
rect 2096 15444 2102 15496
rect 2866 15444 2872 15496
rect 2924 15484 2930 15496
rect 3467 15487 3525 15493
rect 3467 15484 3479 15487
rect 2924 15456 3479 15484
rect 2924 15444 2930 15456
rect 3467 15453 3479 15456
rect 3513 15484 3525 15487
rect 4249 15487 4307 15493
rect 4249 15484 4261 15487
rect 3513 15456 4261 15484
rect 3513 15453 3525 15456
rect 3467 15447 3525 15453
rect 4249 15453 4261 15456
rect 4295 15453 4307 15487
rect 4249 15447 4307 15453
rect 7009 15487 7067 15493
rect 7009 15453 7021 15487
rect 7055 15484 7067 15487
rect 8846 15484 8852 15496
rect 7055 15456 8852 15484
rect 7055 15453 7067 15456
rect 7009 15447 7067 15453
rect 8846 15444 8852 15456
rect 8904 15444 8910 15496
rect 9306 15444 9312 15496
rect 9364 15484 9370 15496
rect 10244 15484 10272 15524
rect 10980 15496 11008 15524
rect 12250 15512 12256 15564
rect 12308 15552 12314 15564
rect 13265 15555 13323 15561
rect 13265 15552 13277 15555
rect 12308 15524 13277 15552
rect 12308 15512 12314 15524
rect 13265 15521 13277 15524
rect 13311 15521 13323 15555
rect 13265 15515 13323 15521
rect 13541 15555 13599 15561
rect 13541 15521 13553 15555
rect 13587 15552 13599 15555
rect 14108 15552 14136 15580
rect 14737 15555 14795 15561
rect 13587 15524 14596 15552
rect 13587 15521 13599 15524
rect 13541 15515 13599 15521
rect 9364 15456 10272 15484
rect 9364 15444 9370 15456
rect 10962 15444 10968 15496
rect 11020 15484 11026 15496
rect 11793 15487 11851 15493
rect 11793 15484 11805 15487
rect 11020 15456 11805 15484
rect 11020 15444 11026 15456
rect 11793 15453 11805 15456
rect 11839 15453 11851 15487
rect 11793 15447 11851 15453
rect 12894 15444 12900 15496
rect 12952 15444 12958 15496
rect 13280 15484 13308 15515
rect 13633 15487 13691 15493
rect 13633 15484 13645 15487
rect 13280 15456 13645 15484
rect 13633 15453 13645 15456
rect 13679 15453 13691 15487
rect 13633 15447 13691 15453
rect 13722 15444 13728 15496
rect 13780 15493 13786 15496
rect 13780 15447 13788 15493
rect 13780 15444 13786 15447
rect 14090 15444 14096 15496
rect 14148 15444 14154 15496
rect 14568 15493 14596 15524
rect 14737 15521 14749 15555
rect 14783 15552 14795 15555
rect 14921 15555 14979 15561
rect 14921 15552 14933 15555
rect 14783 15524 14933 15552
rect 14783 15521 14795 15524
rect 14737 15515 14795 15521
rect 14921 15521 14933 15524
rect 14967 15521 14979 15555
rect 15764 15552 15792 15580
rect 14921 15515 14979 15521
rect 15028 15524 15792 15552
rect 15028 15493 15056 15524
rect 15856 15496 15884 15660
rect 19794 15648 19800 15700
rect 19852 15648 19858 15700
rect 21358 15648 21364 15700
rect 21416 15688 21422 15700
rect 22925 15691 22983 15697
rect 21416 15660 22784 15688
rect 21416 15648 21422 15660
rect 19705 15623 19763 15629
rect 19705 15589 19717 15623
rect 19751 15620 19763 15623
rect 20346 15620 20352 15632
rect 19751 15592 20352 15620
rect 19751 15589 19763 15592
rect 19705 15583 19763 15589
rect 20346 15580 20352 15592
rect 20404 15580 20410 15632
rect 22646 15580 22652 15632
rect 22704 15580 22710 15632
rect 15933 15555 15991 15561
rect 15933 15521 15945 15555
rect 15979 15552 15991 15555
rect 16574 15552 16580 15564
rect 15979 15524 16580 15552
rect 15979 15521 15991 15524
rect 15933 15515 15991 15521
rect 16574 15512 16580 15524
rect 16632 15512 16638 15564
rect 20714 15552 20720 15564
rect 18248 15524 20720 15552
rect 14277 15487 14335 15493
rect 14277 15453 14289 15487
rect 14323 15453 14335 15487
rect 14277 15447 14335 15453
rect 14553 15487 14611 15493
rect 14553 15453 14565 15487
rect 14599 15453 14611 15487
rect 14553 15447 14611 15453
rect 15013 15487 15071 15493
rect 15013 15453 15025 15487
rect 15059 15453 15071 15487
rect 15013 15447 15071 15453
rect 3326 15416 3332 15428
rect 3082 15388 3332 15416
rect 3326 15376 3332 15388
rect 3384 15416 3390 15428
rect 3970 15416 3976 15428
rect 3384 15388 3976 15416
rect 3384 15376 3390 15388
rect 3970 15376 3976 15388
rect 4028 15376 4034 15428
rect 6086 15376 6092 15428
rect 6144 15376 6150 15428
rect 11330 15416 11336 15428
rect 9324 15388 9904 15416
rect 11178 15388 11336 15416
rect 1581 15351 1639 15357
rect 1581 15317 1593 15351
rect 1627 15348 1639 15351
rect 2958 15348 2964 15360
rect 1627 15320 2964 15348
rect 1627 15317 1639 15320
rect 1581 15311 1639 15317
rect 2958 15308 2964 15320
rect 3016 15308 3022 15360
rect 3602 15308 3608 15360
rect 3660 15348 3666 15360
rect 3789 15351 3847 15357
rect 3789 15348 3801 15351
rect 3660 15320 3801 15348
rect 3660 15308 3666 15320
rect 3789 15317 3801 15320
rect 3835 15317 3847 15351
rect 3789 15311 3847 15317
rect 4157 15351 4215 15357
rect 4157 15317 4169 15351
rect 4203 15348 4215 15351
rect 4430 15348 4436 15360
rect 4203 15320 4436 15348
rect 4203 15317 4215 15320
rect 4157 15311 4215 15317
rect 4430 15308 4436 15320
rect 4488 15308 4494 15360
rect 7653 15351 7711 15357
rect 7653 15317 7665 15351
rect 7699 15348 7711 15351
rect 7834 15348 7840 15360
rect 7699 15320 7840 15348
rect 7699 15317 7711 15320
rect 7653 15311 7711 15317
rect 7834 15308 7840 15320
rect 7892 15308 7898 15360
rect 8021 15351 8079 15357
rect 8021 15317 8033 15351
rect 8067 15348 8079 15351
rect 9214 15348 9220 15360
rect 8067 15320 9220 15348
rect 8067 15317 8079 15320
rect 8021 15311 8079 15317
rect 9214 15308 9220 15320
rect 9272 15308 9278 15360
rect 9324 15357 9352 15388
rect 9309 15351 9367 15357
rect 9309 15317 9321 15351
rect 9355 15317 9367 15351
rect 9309 15311 9367 15317
rect 9674 15308 9680 15360
rect 9732 15308 9738 15360
rect 9876 15348 9904 15388
rect 10686 15348 10692 15360
rect 9876 15320 10692 15348
rect 10686 15308 10692 15320
rect 10744 15308 10750 15360
rect 10778 15308 10784 15360
rect 10836 15348 10842 15360
rect 11256 15348 11284 15388
rect 11330 15376 11336 15388
rect 11388 15416 11394 15428
rect 11977 15419 12035 15425
rect 11977 15416 11989 15419
rect 11388 15388 11989 15416
rect 11388 15376 11394 15388
rect 11977 15385 11989 15388
rect 12023 15385 12035 15419
rect 11977 15379 12035 15385
rect 13004 15388 13308 15416
rect 10836 15320 11284 15348
rect 11563 15351 11621 15357
rect 10836 15308 10842 15320
rect 11563 15317 11575 15351
rect 11609 15348 11621 15351
rect 12250 15348 12256 15360
rect 11609 15320 12256 15348
rect 11609 15317 11621 15320
rect 11563 15311 11621 15317
rect 12250 15308 12256 15320
rect 12308 15308 12314 15360
rect 12526 15308 12532 15360
rect 12584 15348 12590 15360
rect 13004 15357 13032 15388
rect 12989 15351 13047 15357
rect 12989 15348 13001 15351
rect 12584 15320 13001 15348
rect 12584 15308 12590 15320
rect 12989 15317 13001 15320
rect 13035 15317 13047 15351
rect 12989 15311 13047 15317
rect 13081 15351 13139 15357
rect 13081 15317 13093 15351
rect 13127 15348 13139 15351
rect 13170 15348 13176 15360
rect 13127 15320 13176 15348
rect 13127 15317 13139 15320
rect 13081 15311 13139 15317
rect 13170 15308 13176 15320
rect 13228 15308 13234 15360
rect 13280 15348 13308 15388
rect 13354 15376 13360 15428
rect 13412 15376 13418 15428
rect 13541 15419 13599 15425
rect 13541 15385 13553 15419
rect 13587 15385 13599 15419
rect 13541 15379 13599 15385
rect 13446 15348 13452 15360
rect 13280 15320 13452 15348
rect 13446 15308 13452 15320
rect 13504 15348 13510 15360
rect 13556 15348 13584 15379
rect 13814 15376 13820 15428
rect 13872 15416 13878 15428
rect 14292 15416 14320 15447
rect 15470 15444 15476 15496
rect 15528 15444 15534 15496
rect 15562 15444 15568 15496
rect 15620 15444 15626 15496
rect 15749 15487 15807 15493
rect 15749 15453 15761 15487
rect 15795 15484 15807 15487
rect 15838 15484 15844 15496
rect 15795 15456 15844 15484
rect 15795 15453 15807 15456
rect 15749 15447 15807 15453
rect 15838 15444 15844 15456
rect 15896 15444 15902 15496
rect 16298 15444 16304 15496
rect 16356 15444 16362 15496
rect 18248 15493 18276 15524
rect 20714 15512 20720 15524
rect 20772 15512 20778 15564
rect 20898 15512 20904 15564
rect 20956 15552 20962 15564
rect 21818 15552 21824 15564
rect 20956 15524 21824 15552
rect 20956 15512 20962 15524
rect 21818 15512 21824 15524
rect 21876 15512 21882 15564
rect 22756 15552 22784 15660
rect 22925 15657 22937 15691
rect 22971 15688 22983 15691
rect 23106 15688 23112 15700
rect 22971 15660 23112 15688
rect 22971 15657 22983 15660
rect 22925 15651 22983 15657
rect 23106 15648 23112 15660
rect 23164 15648 23170 15700
rect 23382 15648 23388 15700
rect 23440 15688 23446 15700
rect 24581 15691 24639 15697
rect 24581 15688 24593 15691
rect 23440 15660 24593 15688
rect 23440 15648 23446 15660
rect 24581 15657 24593 15660
rect 24627 15657 24639 15691
rect 24581 15651 24639 15657
rect 23198 15580 23204 15632
rect 23256 15620 23262 15632
rect 24029 15623 24087 15629
rect 24029 15620 24041 15623
rect 23256 15592 24041 15620
rect 23256 15580 23262 15592
rect 24029 15589 24041 15592
rect 24075 15589 24087 15623
rect 24029 15583 24087 15589
rect 23477 15555 23535 15561
rect 23477 15552 23489 15555
rect 22756 15524 23489 15552
rect 23477 15521 23489 15524
rect 23523 15521 23535 15555
rect 23477 15515 23535 15521
rect 20346 15493 20352 15496
rect 18233 15487 18291 15493
rect 18233 15453 18245 15487
rect 18279 15453 18291 15487
rect 18233 15447 18291 15453
rect 20165 15487 20223 15493
rect 20165 15453 20177 15487
rect 20211 15453 20223 15487
rect 20165 15447 20223 15453
rect 20323 15487 20352 15493
rect 20323 15453 20335 15487
rect 20323 15447 20352 15453
rect 17494 15416 17500 15428
rect 13872 15388 14320 15416
rect 17342 15388 17500 15416
rect 13872 15376 13878 15388
rect 17494 15376 17500 15388
rect 17552 15416 17558 15428
rect 17865 15419 17923 15425
rect 17865 15416 17877 15419
rect 17552 15388 17877 15416
rect 17552 15376 17558 15388
rect 17865 15385 17877 15388
rect 17911 15385 17923 15419
rect 17865 15379 17923 15385
rect 19334 15376 19340 15428
rect 19392 15416 19398 15428
rect 20180 15416 20208 15447
rect 20346 15444 20352 15447
rect 20404 15444 20410 15496
rect 20622 15444 20628 15496
rect 20680 15444 20686 15496
rect 23290 15444 23296 15496
rect 23348 15484 23354 15496
rect 23385 15487 23443 15493
rect 23385 15484 23397 15487
rect 23348 15456 23397 15484
rect 23348 15444 23354 15456
rect 23385 15453 23397 15456
rect 23431 15453 23443 15487
rect 23385 15447 23443 15453
rect 19392 15388 20208 15416
rect 20441 15419 20499 15425
rect 19392 15376 19398 15388
rect 20441 15385 20453 15419
rect 20487 15385 20499 15419
rect 20441 15379 20499 15385
rect 20533 15419 20591 15425
rect 20533 15385 20545 15419
rect 20579 15416 20591 15419
rect 21082 15416 21088 15428
rect 20579 15388 21088 15416
rect 20579 15385 20591 15388
rect 20533 15379 20591 15385
rect 13504 15320 13584 15348
rect 13504 15308 13510 15320
rect 14734 15308 14740 15360
rect 14792 15348 14798 15360
rect 16206 15348 16212 15360
rect 14792 15320 16212 15348
rect 14792 15308 14798 15320
rect 16206 15308 16212 15320
rect 16264 15308 16270 15360
rect 17218 15308 17224 15360
rect 17276 15348 17282 15360
rect 17727 15351 17785 15357
rect 17727 15348 17739 15351
rect 17276 15320 17739 15348
rect 17276 15308 17282 15320
rect 17727 15317 17739 15320
rect 17773 15317 17785 15351
rect 20456 15348 20484 15379
rect 21082 15376 21088 15388
rect 21140 15376 21146 15428
rect 21174 15376 21180 15428
rect 21232 15376 21238 15428
rect 21634 15376 21640 15428
rect 21692 15376 21698 15428
rect 22462 15376 22468 15428
rect 22520 15416 22526 15428
rect 23753 15419 23811 15425
rect 23753 15416 23765 15419
rect 22520 15388 23765 15416
rect 22520 15376 22526 15388
rect 23753 15385 23765 15388
rect 23799 15385 23811 15419
rect 23753 15379 23811 15385
rect 24486 15376 24492 15428
rect 24544 15376 24550 15428
rect 20714 15348 20720 15360
rect 20456 15320 20720 15348
rect 17727 15311 17785 15317
rect 20714 15308 20720 15320
rect 20772 15308 20778 15360
rect 20809 15351 20867 15357
rect 20809 15317 20821 15351
rect 20855 15348 20867 15351
rect 20990 15348 20996 15360
rect 20855 15320 20996 15348
rect 20855 15317 20867 15320
rect 20809 15311 20867 15317
rect 20990 15308 20996 15320
rect 21048 15348 21054 15360
rect 21358 15348 21364 15360
rect 21048 15320 21364 15348
rect 21048 15308 21054 15320
rect 21358 15308 21364 15320
rect 21416 15308 21422 15360
rect 23290 15308 23296 15360
rect 23348 15308 23354 15360
rect 24213 15351 24271 15357
rect 24213 15317 24225 15351
rect 24259 15348 24271 15351
rect 24302 15348 24308 15360
rect 24259 15320 24308 15348
rect 24259 15317 24271 15320
rect 24213 15311 24271 15317
rect 24302 15308 24308 15320
rect 24360 15308 24366 15360
rect 1104 15258 25208 15280
rect 1104 15206 4874 15258
rect 4926 15206 4938 15258
rect 4990 15206 5002 15258
rect 5054 15206 5066 15258
rect 5118 15206 5130 15258
rect 5182 15206 25208 15258
rect 1104 15184 25208 15206
rect 106 15104 112 15156
rect 164 15144 170 15156
rect 15565 15147 15623 15153
rect 164 15116 12940 15144
rect 164 15104 170 15116
rect 2590 15036 2596 15088
rect 2648 15076 2654 15088
rect 2648 15048 3280 15076
rect 2648 15036 2654 15048
rect 2774 14968 2780 15020
rect 2832 14968 2838 15020
rect 2866 14968 2872 15020
rect 2924 14968 2930 15020
rect 3252 15017 3280 15048
rect 3970 15036 3976 15088
rect 4028 15036 4034 15088
rect 5994 15036 6000 15088
rect 6052 15076 6058 15088
rect 6822 15076 6828 15088
rect 6052 15048 6828 15076
rect 6052 15036 6058 15048
rect 6822 15036 6828 15048
rect 6880 15036 6886 15088
rect 8846 15036 8852 15088
rect 8904 15036 8910 15088
rect 10778 15036 10784 15088
rect 10836 15036 10842 15088
rect 12526 15076 12532 15088
rect 11532 15048 12532 15076
rect 3237 15011 3295 15017
rect 3237 14977 3249 15011
rect 3283 14977 3295 15011
rect 3237 14971 3295 14977
rect 3602 14968 3608 15020
rect 3660 14968 3666 15020
rect 6638 14968 6644 15020
rect 6696 15008 6702 15020
rect 6733 15011 6791 15017
rect 6733 15008 6745 15011
rect 6696 14980 6745 15008
rect 6696 14968 6702 14980
rect 6733 14977 6745 14980
rect 6779 14977 6791 15011
rect 6840 15008 6868 15036
rect 11532 15020 11560 15048
rect 12526 15036 12532 15048
rect 12584 15036 12590 15088
rect 12802 15036 12808 15088
rect 12860 15036 12866 15088
rect 12912 15085 12940 15116
rect 15565 15113 15577 15147
rect 15611 15144 15623 15147
rect 15654 15144 15660 15156
rect 15611 15116 15660 15144
rect 15611 15113 15623 15116
rect 15565 15107 15623 15113
rect 15654 15104 15660 15116
rect 15712 15104 15718 15156
rect 15749 15147 15807 15153
rect 15749 15113 15761 15147
rect 15795 15144 15807 15147
rect 16298 15144 16304 15156
rect 15795 15116 16304 15144
rect 15795 15113 15807 15116
rect 15749 15107 15807 15113
rect 16298 15104 16304 15116
rect 16356 15104 16362 15156
rect 18874 15144 18880 15156
rect 16776 15116 18880 15144
rect 16776 15088 16804 15116
rect 18874 15104 18880 15116
rect 18932 15104 18938 15156
rect 22465 15147 22523 15153
rect 22465 15144 22477 15147
rect 22066 15116 22477 15144
rect 12897 15079 12955 15085
rect 12897 15045 12909 15079
rect 12943 15045 12955 15079
rect 12897 15039 12955 15045
rect 14645 15079 14703 15085
rect 14645 15045 14657 15079
rect 14691 15076 14703 15079
rect 16758 15076 16764 15088
rect 14691 15048 16764 15076
rect 14691 15045 14703 15048
rect 14645 15039 14703 15045
rect 7469 15011 7527 15017
rect 6840 14980 6960 15008
rect 6733 14971 6791 14977
rect 3053 14943 3111 14949
rect 3053 14909 3065 14943
rect 3099 14940 3111 14943
rect 3142 14940 3148 14952
rect 3099 14912 3148 14940
rect 3099 14909 3111 14912
rect 3053 14903 3111 14909
rect 3142 14900 3148 14912
rect 3200 14900 3206 14952
rect 6546 14900 6552 14952
rect 6604 14940 6610 14952
rect 6932 14949 6960 14980
rect 7469 14977 7481 15011
rect 7515 15008 7527 15011
rect 7515 14980 7972 15008
rect 7515 14977 7527 14980
rect 7469 14971 7527 14977
rect 6825 14943 6883 14949
rect 6825 14940 6837 14943
rect 6604 14912 6837 14940
rect 6604 14900 6610 14912
rect 6825 14909 6837 14912
rect 6871 14909 6883 14943
rect 6825 14903 6883 14909
rect 6917 14943 6975 14949
rect 6917 14909 6929 14943
rect 6963 14909 6975 14943
rect 6917 14903 6975 14909
rect 7834 14900 7840 14952
rect 7892 14900 7898 14952
rect 7944 14940 7972 14980
rect 9674 14968 9680 15020
rect 9732 15008 9738 15020
rect 9769 15011 9827 15017
rect 9769 15008 9781 15011
rect 9732 14980 9781 15008
rect 9732 14968 9738 14980
rect 9769 14977 9781 14980
rect 9815 14977 9827 15011
rect 9769 14971 9827 14977
rect 10686 14968 10692 15020
rect 10744 15008 10750 15020
rect 11195 15011 11253 15017
rect 11195 15008 11207 15011
rect 10744 14980 11207 15008
rect 10744 14968 10750 14980
rect 11195 14977 11207 14980
rect 11241 15008 11253 15011
rect 11514 15008 11520 15020
rect 11241 14980 11520 15008
rect 11241 14977 11253 14980
rect 11195 14971 11253 14977
rect 11514 14968 11520 14980
rect 11572 14968 11578 15020
rect 12250 14968 12256 15020
rect 12308 14968 12314 15020
rect 12434 14968 12440 15020
rect 12492 14968 12498 15020
rect 12621 15011 12679 15017
rect 12621 14977 12633 15011
rect 12667 15008 12679 15011
rect 12986 15008 12992 15020
rect 12667 14980 12992 15008
rect 12667 14977 12679 14980
rect 12621 14971 12679 14977
rect 12986 14968 12992 14980
rect 13044 15008 13050 15020
rect 13354 15008 13360 15020
rect 13044 14980 13360 15008
rect 13044 14968 13050 14980
rect 13354 14968 13360 14980
rect 13412 14968 13418 15020
rect 8662 14940 8668 14952
rect 7944 14912 8668 14940
rect 8662 14900 8668 14912
rect 8720 14940 8726 14952
rect 9401 14943 9459 14949
rect 9401 14940 9413 14943
rect 8720 14912 9413 14940
rect 8720 14900 8726 14912
rect 9401 14909 9413 14912
rect 9447 14909 9459 14943
rect 9401 14903 9459 14909
rect 11698 14900 11704 14952
rect 11756 14900 11762 14952
rect 14660 14940 14688 15039
rect 16758 15036 16764 15048
rect 16816 15036 16822 15088
rect 18506 15076 18512 15088
rect 18354 15048 18512 15076
rect 18506 15036 18512 15048
rect 18564 15076 18570 15088
rect 18564 15048 20010 15076
rect 18564 15036 18570 15048
rect 20806 15036 20812 15088
rect 20864 15076 20870 15088
rect 22066 15076 22094 15116
rect 22465 15113 22477 15116
rect 22511 15113 22523 15147
rect 22465 15107 22523 15113
rect 20864 15048 22094 15076
rect 20864 15036 20870 15048
rect 22186 15036 22192 15088
rect 22244 15036 22250 15088
rect 23198 15076 23204 15088
rect 22664 15048 23204 15076
rect 14918 14968 14924 15020
rect 14976 14968 14982 15020
rect 15197 15011 15255 15017
rect 15197 14977 15209 15011
rect 15243 15008 15255 15011
rect 15286 15008 15292 15020
rect 15243 14980 15292 15008
rect 15243 14977 15255 14980
rect 15197 14971 15255 14977
rect 15286 14968 15292 14980
rect 15344 14968 15350 15020
rect 15381 15011 15439 15017
rect 15381 14977 15393 15011
rect 15427 15008 15439 15011
rect 15470 15008 15476 15020
rect 15427 14980 15476 15008
rect 15427 14977 15439 14980
rect 15381 14971 15439 14977
rect 15470 14968 15476 14980
rect 15528 14968 15534 15020
rect 15657 15011 15715 15017
rect 15657 14977 15669 15011
rect 15703 14977 15715 15011
rect 15657 14971 15715 14977
rect 11808 14912 14688 14940
rect 14936 14940 14964 14968
rect 15672 14940 15700 14971
rect 15746 14968 15752 15020
rect 15804 15008 15810 15020
rect 15933 15011 15991 15017
rect 15933 15008 15945 15011
rect 15804 14980 15945 15008
rect 15804 14968 15810 14980
rect 15933 14977 15945 14980
rect 15979 14977 15991 15011
rect 15933 14971 15991 14977
rect 16022 14968 16028 15020
rect 16080 14968 16086 15020
rect 16206 14968 16212 15020
rect 16264 15008 16270 15020
rect 16301 15011 16359 15017
rect 16301 15008 16313 15011
rect 16264 14980 16313 15008
rect 16264 14968 16270 14980
rect 16301 14977 16313 14980
rect 16347 14977 16359 15011
rect 16301 14971 16359 14977
rect 16393 15011 16451 15017
rect 16393 14977 16405 15011
rect 16439 15008 16451 15011
rect 17218 15008 17224 15020
rect 16439 14980 17224 15008
rect 16439 14977 16451 14980
rect 16393 14971 16451 14977
rect 17218 14968 17224 14980
rect 17276 14968 17282 15020
rect 21453 15011 21511 15017
rect 21453 14977 21465 15011
rect 21499 14977 21511 15011
rect 21453 14971 21511 14977
rect 21637 15011 21695 15017
rect 21637 14977 21649 15011
rect 21683 15008 21695 15011
rect 22097 15011 22155 15017
rect 22097 15008 22109 15011
rect 21683 14980 22109 15008
rect 21683 14977 21695 14980
rect 21637 14971 21695 14977
rect 22097 14977 22109 14980
rect 22143 15008 22155 15011
rect 22204 15008 22232 15036
rect 22143 14980 22232 15008
rect 22281 15011 22339 15017
rect 22143 14977 22155 14980
rect 22097 14971 22155 14977
rect 22281 14977 22293 15011
rect 22327 15008 22339 15011
rect 22554 15008 22560 15020
rect 22327 14980 22560 15008
rect 22327 14977 22339 14980
rect 22281 14971 22339 14977
rect 14936 14912 15700 14940
rect 4430 14832 4436 14884
rect 4488 14872 4494 14884
rect 5031 14875 5089 14881
rect 5031 14872 5043 14875
rect 4488 14844 5043 14872
rect 4488 14832 4494 14844
rect 5031 14841 5043 14844
rect 5077 14872 5089 14875
rect 5077 14844 6592 14872
rect 5077 14841 5089 14844
rect 5031 14835 5089 14841
rect 1762 14764 1768 14816
rect 1820 14804 1826 14816
rect 2409 14807 2467 14813
rect 2409 14804 2421 14807
rect 1820 14776 2421 14804
rect 1820 14764 1826 14776
rect 2409 14773 2421 14776
rect 2455 14773 2467 14807
rect 2409 14767 2467 14773
rect 4706 14764 4712 14816
rect 4764 14804 4770 14816
rect 5350 14804 5356 14816
rect 4764 14776 5356 14804
rect 4764 14764 4770 14776
rect 5350 14764 5356 14776
rect 5408 14764 5414 14816
rect 6365 14807 6423 14813
rect 6365 14773 6377 14807
rect 6411 14804 6423 14807
rect 6454 14804 6460 14816
rect 6411 14776 6460 14804
rect 6411 14773 6423 14776
rect 6365 14767 6423 14773
rect 6454 14764 6460 14776
rect 6512 14764 6518 14816
rect 6564 14804 6592 14844
rect 8938 14832 8944 14884
rect 8996 14872 9002 14884
rect 11808 14872 11836 14912
rect 16574 14900 16580 14952
rect 16632 14940 16638 14952
rect 16945 14943 17003 14949
rect 16945 14940 16957 14943
rect 16632 14912 16957 14940
rect 16632 14900 16638 14912
rect 16945 14909 16957 14912
rect 16991 14909 17003 14943
rect 16945 14903 17003 14909
rect 17310 14900 17316 14952
rect 17368 14900 17374 14952
rect 19245 14943 19303 14949
rect 19245 14909 19257 14943
rect 19291 14909 19303 14943
rect 19245 14903 19303 14909
rect 8996 14844 9444 14872
rect 8996 14832 9002 14844
rect 7650 14804 7656 14816
rect 6564 14776 7656 14804
rect 7650 14764 7656 14776
rect 7708 14764 7714 14816
rect 9214 14764 9220 14816
rect 9272 14813 9278 14816
rect 9272 14807 9321 14813
rect 9272 14773 9275 14807
rect 9309 14773 9321 14807
rect 9416 14804 9444 14844
rect 11072 14844 11836 14872
rect 11072 14804 11100 14844
rect 12066 14832 12072 14884
rect 12124 14832 12130 14884
rect 9416 14776 11100 14804
rect 12161 14807 12219 14813
rect 9272 14767 9321 14773
rect 12161 14773 12173 14807
rect 12207 14804 12219 14807
rect 12434 14804 12440 14816
rect 12207 14776 12440 14804
rect 12207 14773 12219 14776
rect 12161 14767 12219 14773
rect 9272 14764 9278 14767
rect 12434 14764 12440 14776
rect 12492 14764 12498 14816
rect 12618 14764 12624 14816
rect 12676 14804 12682 14816
rect 13170 14804 13176 14816
rect 12676 14776 13176 14804
rect 12676 14764 12682 14776
rect 13170 14764 13176 14776
rect 13228 14764 13234 14816
rect 13262 14764 13268 14816
rect 13320 14804 13326 14816
rect 14737 14807 14795 14813
rect 14737 14804 14749 14807
rect 13320 14776 14749 14804
rect 13320 14764 13326 14776
rect 14737 14773 14749 14776
rect 14783 14773 14795 14807
rect 14737 14767 14795 14773
rect 18046 14764 18052 14816
rect 18104 14804 18110 14816
rect 18739 14807 18797 14813
rect 18739 14804 18751 14807
rect 18104 14776 18751 14804
rect 18104 14764 18110 14776
rect 18739 14773 18751 14776
rect 18785 14773 18797 14807
rect 19260 14804 19288 14903
rect 19518 14900 19524 14952
rect 19576 14900 19582 14952
rect 21266 14900 21272 14952
rect 21324 14900 21330 14952
rect 21468 14940 21496 14971
rect 22186 14940 22192 14952
rect 21468 14912 22192 14940
rect 22186 14900 22192 14912
rect 22244 14940 22250 14952
rect 22296 14940 22324 14971
rect 22554 14968 22560 14980
rect 22612 14968 22618 15020
rect 22664 15017 22692 15048
rect 23198 15036 23204 15048
rect 23256 15036 23262 15088
rect 24302 15036 24308 15088
rect 24360 15076 24366 15088
rect 24581 15079 24639 15085
rect 24581 15076 24593 15079
rect 24360 15048 24593 15076
rect 24360 15036 24366 15048
rect 24581 15045 24593 15048
rect 24627 15045 24639 15079
rect 24581 15039 24639 15045
rect 22649 15011 22707 15017
rect 22649 14977 22661 15011
rect 22695 14977 22707 15011
rect 22649 14971 22707 14977
rect 22922 14968 22928 15020
rect 22980 14968 22986 15020
rect 23474 14968 23480 15020
rect 23532 14968 23538 15020
rect 22244 14912 22324 14940
rect 22741 14943 22799 14949
rect 22244 14900 22250 14912
rect 22741 14909 22753 14943
rect 22787 14909 22799 14943
rect 22741 14903 22799 14909
rect 21284 14872 21312 14900
rect 22554 14872 22560 14884
rect 21284 14844 22560 14872
rect 22554 14832 22560 14844
rect 22612 14872 22618 14884
rect 22756 14872 22784 14903
rect 24854 14900 24860 14952
rect 24912 14900 24918 14952
rect 22612 14844 22784 14872
rect 22612 14832 22618 14844
rect 20898 14804 20904 14816
rect 19260 14776 20904 14804
rect 18739 14767 18797 14773
rect 20898 14764 20904 14776
rect 20956 14764 20962 14816
rect 21637 14807 21695 14813
rect 21637 14773 21649 14807
rect 21683 14804 21695 14807
rect 21726 14804 21732 14816
rect 21683 14776 21732 14804
rect 21683 14773 21695 14776
rect 21637 14767 21695 14773
rect 21726 14764 21732 14776
rect 21784 14764 21790 14816
rect 21910 14764 21916 14816
rect 21968 14764 21974 14816
rect 22278 14764 22284 14816
rect 22336 14804 22342 14816
rect 22649 14807 22707 14813
rect 22649 14804 22661 14807
rect 22336 14776 22661 14804
rect 22336 14764 22342 14776
rect 22649 14773 22661 14776
rect 22695 14804 22707 14807
rect 23109 14807 23167 14813
rect 23109 14804 23121 14807
rect 22695 14776 23121 14804
rect 22695 14773 22707 14776
rect 22649 14767 22707 14773
rect 23109 14773 23121 14776
rect 23155 14773 23167 14807
rect 23109 14767 23167 14773
rect 1104 14714 25208 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 25208 14714
rect 1104 14640 25208 14662
rect 2774 14560 2780 14612
rect 2832 14600 2838 14612
rect 3234 14609 3240 14612
rect 3191 14603 3240 14609
rect 3191 14600 3203 14603
rect 2832 14572 3203 14600
rect 2832 14560 2838 14572
rect 3191 14569 3203 14572
rect 3237 14569 3240 14603
rect 3191 14563 3240 14569
rect 3234 14560 3240 14563
rect 3292 14560 3298 14612
rect 5031 14603 5089 14609
rect 5031 14569 5043 14603
rect 5077 14600 5089 14603
rect 5902 14600 5908 14612
rect 5077 14572 5908 14600
rect 5077 14569 5089 14572
rect 5031 14563 5089 14569
rect 5902 14560 5908 14572
rect 5960 14600 5966 14612
rect 6638 14600 6644 14612
rect 5960 14572 6644 14600
rect 5960 14560 5966 14572
rect 6638 14560 6644 14572
rect 6696 14560 6702 14612
rect 12342 14600 12348 14612
rect 11440 14572 12348 14600
rect 6822 14492 6828 14544
rect 6880 14532 6886 14544
rect 7745 14535 7803 14541
rect 7745 14532 7757 14535
rect 6880 14504 7757 14532
rect 6880 14492 6886 14504
rect 7745 14501 7757 14504
rect 7791 14501 7803 14535
rect 7745 14495 7803 14501
rect 1762 14424 1768 14476
rect 1820 14424 1826 14476
rect 3142 14424 3148 14476
rect 3200 14464 3206 14476
rect 4709 14467 4767 14473
rect 4709 14464 4721 14467
rect 3200 14436 4721 14464
rect 3200 14424 3206 14436
rect 4709 14433 4721 14436
rect 4755 14464 4767 14467
rect 5994 14464 6000 14476
rect 4755 14436 6000 14464
rect 4755 14433 4767 14436
rect 4709 14427 4767 14433
rect 5994 14424 6000 14436
rect 6052 14424 6058 14476
rect 6454 14424 6460 14476
rect 6512 14424 6518 14476
rect 6914 14424 6920 14476
rect 6972 14464 6978 14476
rect 7469 14467 7527 14473
rect 7469 14464 7481 14467
rect 6972 14436 7481 14464
rect 6972 14424 6978 14436
rect 7469 14433 7481 14436
rect 7515 14433 7527 14467
rect 7469 14427 7527 14433
rect 1397 14399 1455 14405
rect 1397 14365 1409 14399
rect 1443 14396 1455 14399
rect 1670 14396 1676 14408
rect 1443 14368 1676 14396
rect 1443 14365 1455 14368
rect 1397 14359 1455 14365
rect 1670 14356 1676 14368
rect 1728 14356 1734 14408
rect 3326 14396 3332 14408
rect 2792 14368 3332 14396
rect 2792 14314 2820 14368
rect 3326 14356 3332 14368
rect 3384 14396 3390 14408
rect 5626 14396 5632 14408
rect 3384 14368 5632 14396
rect 3384 14356 3390 14368
rect 5626 14356 5632 14368
rect 5684 14356 5690 14408
rect 6546 14356 6552 14408
rect 6604 14396 6610 14408
rect 6604 14368 6776 14396
rect 6604 14356 6610 14368
rect 6086 14288 6092 14340
rect 6144 14288 6150 14340
rect 6748 14328 6776 14368
rect 6822 14356 6828 14408
rect 6880 14396 6886 14408
rect 8110 14396 8116 14408
rect 6880 14368 8116 14396
rect 6880 14356 6886 14368
rect 8110 14356 8116 14368
rect 8168 14396 8174 14408
rect 9217 14399 9275 14405
rect 9217 14396 9229 14399
rect 8168 14368 9229 14396
rect 8168 14356 8174 14368
rect 9217 14365 9229 14368
rect 9263 14365 9275 14399
rect 9217 14359 9275 14365
rect 9585 14399 9643 14405
rect 9585 14365 9597 14399
rect 9631 14396 9643 14399
rect 9674 14396 9680 14408
rect 9631 14368 9680 14396
rect 9631 14365 9643 14368
rect 9585 14359 9643 14365
rect 9674 14356 9680 14368
rect 9732 14356 9738 14408
rect 11440 14340 11468 14572
rect 12342 14560 12348 14572
rect 12400 14560 12406 14612
rect 13814 14560 13820 14612
rect 13872 14600 13878 14612
rect 14277 14603 14335 14609
rect 14277 14600 14289 14603
rect 13872 14572 14289 14600
rect 13872 14560 13878 14572
rect 14277 14569 14289 14572
rect 14323 14569 14335 14603
rect 14277 14563 14335 14569
rect 14461 14603 14519 14609
rect 14461 14569 14473 14603
rect 14507 14600 14519 14603
rect 14918 14600 14924 14612
rect 14507 14572 14924 14600
rect 14507 14569 14519 14572
rect 14461 14563 14519 14569
rect 14918 14560 14924 14572
rect 14976 14560 14982 14612
rect 15473 14603 15531 14609
rect 15473 14569 15485 14603
rect 15519 14600 15531 14603
rect 15838 14600 15844 14612
rect 15519 14572 15844 14600
rect 15519 14569 15531 14572
rect 15473 14563 15531 14569
rect 15838 14560 15844 14572
rect 15896 14560 15902 14612
rect 17310 14560 17316 14612
rect 17368 14560 17374 14612
rect 19518 14560 19524 14612
rect 19576 14600 19582 14612
rect 20441 14603 20499 14609
rect 20441 14600 20453 14603
rect 19576 14572 20453 14600
rect 19576 14560 19582 14572
rect 20441 14569 20453 14572
rect 20487 14569 20499 14603
rect 20441 14563 20499 14569
rect 21358 14560 21364 14612
rect 21416 14600 21422 14612
rect 21729 14603 21787 14609
rect 21729 14600 21741 14603
rect 21416 14572 21741 14600
rect 21416 14560 21422 14572
rect 21729 14569 21741 14572
rect 21775 14600 21787 14603
rect 22002 14600 22008 14612
rect 21775 14572 22008 14600
rect 21775 14569 21787 14572
rect 21729 14563 21787 14569
rect 22002 14560 22008 14572
rect 22060 14560 22066 14612
rect 22370 14560 22376 14612
rect 22428 14600 22434 14612
rect 22741 14603 22799 14609
rect 22741 14600 22753 14603
rect 22428 14572 22753 14600
rect 22428 14560 22434 14572
rect 22741 14569 22753 14572
rect 22787 14569 22799 14603
rect 22741 14563 22799 14569
rect 22925 14603 22983 14609
rect 22925 14569 22937 14603
rect 22971 14569 22983 14603
rect 22925 14563 22983 14569
rect 12066 14492 12072 14544
rect 12124 14492 12130 14544
rect 14090 14492 14096 14544
rect 14148 14532 14154 14544
rect 14829 14535 14887 14541
rect 14829 14532 14841 14535
rect 14148 14504 14841 14532
rect 14148 14492 14154 14504
rect 14829 14501 14841 14504
rect 14875 14501 14887 14535
rect 21082 14532 21088 14544
rect 14829 14495 14887 14501
rect 15304 14504 17908 14532
rect 12434 14424 12440 14476
rect 12492 14424 12498 14476
rect 12897 14467 12955 14473
rect 12897 14464 12909 14467
rect 12636 14436 12909 14464
rect 11514 14356 11520 14408
rect 11572 14356 11578 14408
rect 11606 14356 11612 14408
rect 11664 14396 11670 14408
rect 11885 14399 11943 14405
rect 11885 14396 11897 14399
rect 11664 14368 11897 14396
rect 11664 14356 11670 14368
rect 11885 14365 11897 14368
rect 11931 14365 11943 14399
rect 11885 14359 11943 14365
rect 12345 14399 12403 14405
rect 12345 14365 12357 14399
rect 12391 14365 12403 14399
rect 12345 14359 12403 14365
rect 7285 14331 7343 14337
rect 7285 14328 7297 14331
rect 6748 14300 7297 14328
rect 7285 14297 7297 14300
rect 7331 14297 7343 14331
rect 7285 14291 7343 14297
rect 7929 14331 7987 14337
rect 7929 14297 7941 14331
rect 7975 14328 7987 14331
rect 9306 14328 9312 14340
rect 7975 14300 9312 14328
rect 7975 14297 7987 14300
rect 7929 14291 7987 14297
rect 9306 14288 9312 14300
rect 9364 14288 9370 14340
rect 10134 14288 10140 14340
rect 10192 14288 10198 14340
rect 11422 14288 11428 14340
rect 11480 14328 11486 14340
rect 11701 14331 11759 14337
rect 11701 14328 11713 14331
rect 11480 14300 11713 14328
rect 11480 14288 11486 14300
rect 11701 14297 11713 14300
rect 11747 14297 11759 14331
rect 11701 14291 11759 14297
rect 11790 14288 11796 14340
rect 11848 14328 11854 14340
rect 12250 14328 12256 14340
rect 11848 14300 12256 14328
rect 11848 14288 11854 14300
rect 12250 14288 12256 14300
rect 12308 14288 12314 14340
rect 12360 14328 12388 14359
rect 12636 14328 12664 14436
rect 12897 14433 12909 14436
rect 12943 14433 12955 14467
rect 12897 14427 12955 14433
rect 14182 14424 14188 14476
rect 14240 14464 14246 14476
rect 15197 14467 15255 14473
rect 15197 14464 15209 14467
rect 14240 14436 15209 14464
rect 14240 14424 14246 14436
rect 15197 14433 15209 14436
rect 15243 14433 15255 14467
rect 15197 14427 15255 14433
rect 12805 14399 12863 14405
rect 12805 14365 12817 14399
rect 12851 14365 12863 14399
rect 12805 14359 12863 14365
rect 12360 14300 12664 14328
rect 12820 14272 12848 14359
rect 12986 14356 12992 14408
rect 13044 14356 13050 14408
rect 13078 14356 13084 14408
rect 13136 14356 13142 14408
rect 13170 14356 13176 14408
rect 13228 14396 13234 14408
rect 13354 14396 13360 14408
rect 13228 14368 13360 14396
rect 13228 14356 13234 14368
rect 13354 14356 13360 14368
rect 13412 14356 13418 14408
rect 13446 14356 13452 14408
rect 13504 14356 13510 14408
rect 15013 14399 15071 14405
rect 15013 14396 15025 14399
rect 13547 14368 15025 14396
rect 13004 14328 13032 14356
rect 13265 14331 13323 14337
rect 13265 14328 13277 14331
rect 13004 14300 13277 14328
rect 13265 14297 13277 14300
rect 13311 14297 13323 14331
rect 13265 14291 13323 14297
rect 4157 14263 4215 14269
rect 4157 14229 4169 14263
rect 4203 14260 4215 14263
rect 4430 14260 4436 14272
rect 4203 14232 4436 14260
rect 4203 14229 4215 14232
rect 4157 14223 4215 14229
rect 4430 14220 4436 14232
rect 4488 14220 4494 14272
rect 4522 14220 4528 14272
rect 4580 14220 4586 14272
rect 4617 14263 4675 14269
rect 4617 14229 4629 14263
rect 4663 14260 4675 14263
rect 4706 14260 4712 14272
rect 4663 14232 4712 14260
rect 4663 14229 4675 14232
rect 4617 14223 4675 14229
rect 4706 14220 4712 14232
rect 4764 14220 4770 14272
rect 5534 14220 5540 14272
rect 5592 14260 5598 14272
rect 6917 14263 6975 14269
rect 6917 14260 6929 14263
rect 5592 14232 6929 14260
rect 5592 14220 5598 14232
rect 6917 14229 6929 14232
rect 6963 14229 6975 14263
rect 6917 14223 6975 14229
rect 7374 14220 7380 14272
rect 7432 14220 7438 14272
rect 10410 14220 10416 14272
rect 10468 14260 10474 14272
rect 11011 14263 11069 14269
rect 11011 14260 11023 14263
rect 10468 14232 11023 14260
rect 10468 14220 10474 14232
rect 11011 14229 11023 14232
rect 11057 14260 11069 14263
rect 12618 14260 12624 14272
rect 11057 14232 12624 14260
rect 11057 14229 11069 14232
rect 11011 14223 11069 14229
rect 12618 14220 12624 14232
rect 12676 14220 12682 14272
rect 12710 14220 12716 14272
rect 12768 14220 12774 14272
rect 12802 14220 12808 14272
rect 12860 14260 12866 14272
rect 13547 14260 13575 14368
rect 15013 14365 15025 14368
rect 15059 14365 15071 14399
rect 15013 14359 15071 14365
rect 15304 14340 15332 14504
rect 17770 14424 17776 14476
rect 17828 14424 17834 14476
rect 17880 14473 17908 14504
rect 20916 14504 21088 14532
rect 20916 14473 20944 14504
rect 21082 14492 21088 14504
rect 21140 14532 21146 14544
rect 21266 14532 21272 14544
rect 21140 14504 21272 14532
rect 21140 14492 21146 14504
rect 21266 14492 21272 14504
rect 21324 14492 21330 14544
rect 22940 14532 22968 14563
rect 23290 14560 23296 14612
rect 23348 14560 23354 14612
rect 22940 14504 23428 14532
rect 17865 14467 17923 14473
rect 17865 14433 17877 14467
rect 17911 14433 17923 14467
rect 17865 14427 17923 14433
rect 20901 14467 20959 14473
rect 20901 14433 20913 14467
rect 20947 14433 20959 14467
rect 20901 14427 20959 14433
rect 20990 14424 20996 14476
rect 21048 14424 21054 14476
rect 23400 14408 23428 14504
rect 17681 14399 17739 14405
rect 17681 14365 17693 14399
rect 17727 14396 17739 14399
rect 18046 14396 18052 14408
rect 17727 14368 18052 14396
rect 17727 14365 17739 14368
rect 17681 14359 17739 14365
rect 18046 14356 18052 14368
rect 18104 14356 18110 14408
rect 20809 14399 20867 14405
rect 20809 14365 20821 14399
rect 20855 14396 20867 14399
rect 21634 14396 21640 14408
rect 20855 14368 21640 14396
rect 20855 14365 20867 14368
rect 20809 14359 20867 14365
rect 21634 14356 21640 14368
rect 21692 14356 21698 14408
rect 21726 14356 21732 14408
rect 21784 14356 21790 14408
rect 21910 14356 21916 14408
rect 21968 14356 21974 14408
rect 22186 14356 22192 14408
rect 22244 14356 22250 14408
rect 22278 14356 22284 14408
rect 22336 14396 22342 14408
rect 22373 14399 22431 14405
rect 22373 14396 22385 14399
rect 22336 14368 22385 14396
rect 22336 14356 22342 14368
rect 22373 14365 22385 14368
rect 22419 14365 22431 14399
rect 23014 14396 23020 14408
rect 22924 14371 23020 14396
rect 22373 14359 22431 14365
rect 22879 14368 23020 14371
rect 22879 14365 22952 14368
rect 13722 14288 13728 14340
rect 13780 14328 13786 14340
rect 14090 14328 14096 14340
rect 13780 14300 14096 14328
rect 13780 14288 13786 14300
rect 14090 14288 14096 14300
rect 14148 14288 14154 14340
rect 14200 14300 14964 14328
rect 12860 14232 13575 14260
rect 13633 14263 13691 14269
rect 12860 14220 12866 14232
rect 13633 14229 13645 14263
rect 13679 14260 13691 14263
rect 14200 14260 14228 14300
rect 13679 14232 14228 14260
rect 13679 14229 13691 14232
rect 13633 14223 13691 14229
rect 14274 14220 14280 14272
rect 14332 14269 14338 14272
rect 14332 14263 14351 14269
rect 14339 14229 14351 14263
rect 14936 14260 14964 14300
rect 15286 14288 15292 14340
rect 15344 14288 15350 14340
rect 20990 14288 20996 14340
rect 21048 14328 21054 14340
rect 22005 14331 22063 14337
rect 22005 14328 22017 14331
rect 21048 14300 22017 14328
rect 21048 14288 21054 14300
rect 22005 14297 22017 14300
rect 22051 14297 22063 14331
rect 22879 14331 22891 14365
rect 22925 14334 22952 14365
rect 23014 14356 23020 14368
rect 23072 14396 23078 14408
rect 23201 14399 23259 14405
rect 23201 14396 23213 14399
rect 23072 14368 23213 14396
rect 23072 14356 23078 14368
rect 23201 14365 23213 14368
rect 23247 14365 23259 14399
rect 23201 14359 23259 14365
rect 23382 14356 23388 14408
rect 23440 14356 23446 14408
rect 22925 14331 22937 14334
rect 22879 14325 22937 14331
rect 22005 14291 22063 14297
rect 23106 14288 23112 14340
rect 23164 14288 23170 14340
rect 15489 14263 15547 14269
rect 15489 14260 15501 14263
rect 14936 14232 15501 14260
rect 14332 14223 14351 14229
rect 15489 14229 15501 14232
rect 15535 14229 15547 14263
rect 15489 14223 15547 14229
rect 15657 14263 15715 14269
rect 15657 14229 15669 14263
rect 15703 14260 15715 14263
rect 15746 14260 15752 14272
rect 15703 14232 15752 14260
rect 15703 14229 15715 14232
rect 15657 14223 15715 14229
rect 14332 14220 14338 14223
rect 15746 14220 15752 14232
rect 15804 14220 15810 14272
rect 1104 14170 25208 14192
rect 1104 14118 4874 14170
rect 4926 14118 4938 14170
rect 4990 14118 5002 14170
rect 5054 14118 5066 14170
rect 5118 14118 5130 14170
rect 5182 14118 25208 14170
rect 1104 14096 25208 14118
rect 1581 14059 1639 14065
rect 1581 14025 1593 14059
rect 1627 14056 1639 14059
rect 1762 14056 1768 14068
rect 1627 14028 1768 14056
rect 1627 14025 1639 14028
rect 1581 14019 1639 14025
rect 1762 14016 1768 14028
rect 1820 14016 1826 14068
rect 4522 14016 4528 14068
rect 4580 14056 4586 14068
rect 5859 14059 5917 14065
rect 5859 14056 5871 14059
rect 4580 14028 5871 14056
rect 4580 14016 4586 14028
rect 5859 14025 5871 14028
rect 5905 14056 5917 14059
rect 6825 14059 6883 14065
rect 6825 14056 6837 14059
rect 5905 14028 6837 14056
rect 5905 14025 5917 14028
rect 5859 14019 5917 14025
rect 6825 14025 6837 14028
rect 6871 14056 6883 14059
rect 7374 14056 7380 14068
rect 6871 14028 7380 14056
rect 6871 14025 6883 14028
rect 6825 14019 6883 14025
rect 7374 14016 7380 14028
rect 7432 14016 7438 14068
rect 8202 14016 8208 14068
rect 8260 14056 8266 14068
rect 8260 14028 8800 14056
rect 8260 14016 8266 14028
rect 3326 13948 3332 14000
rect 3384 13948 3390 14000
rect 842 13880 848 13932
rect 900 13920 906 13932
rect 1397 13923 1455 13929
rect 1397 13920 1409 13923
rect 900 13892 1409 13920
rect 900 13880 906 13892
rect 1397 13889 1409 13892
rect 1443 13889 1455 13923
rect 1397 13883 1455 13889
rect 1670 13880 1676 13932
rect 1728 13920 1734 13932
rect 1949 13923 2007 13929
rect 1949 13920 1961 13923
rect 1728 13892 1961 13920
rect 1728 13880 1734 13892
rect 1949 13889 1961 13892
rect 1995 13920 2007 13923
rect 3743 13923 3801 13929
rect 1995 13892 2452 13920
rect 1995 13889 2007 13892
rect 1949 13883 2007 13889
rect 2314 13812 2320 13864
rect 2372 13812 2378 13864
rect 2424 13852 2452 13892
rect 3743 13889 3755 13923
rect 3789 13920 3801 13923
rect 3789 13892 4200 13920
rect 3789 13889 3801 13892
rect 3743 13883 3801 13889
rect 4065 13855 4123 13861
rect 4065 13852 4077 13855
rect 2424 13824 4077 13852
rect 4065 13821 4077 13824
rect 4111 13821 4123 13855
rect 4172 13852 4200 13892
rect 4430 13880 4436 13932
rect 4488 13880 4494 13932
rect 5460 13920 5488 13974
rect 6638 13948 6644 14000
rect 6696 13988 6702 14000
rect 7653 13991 7711 13997
rect 7653 13988 7665 13991
rect 6696 13960 7665 13988
rect 6696 13948 6702 13960
rect 7653 13957 7665 13960
rect 7699 13957 7711 13991
rect 8772 13988 8800 14028
rect 9674 14016 9680 14068
rect 9732 14056 9738 14068
rect 10045 14059 10103 14065
rect 10045 14056 10057 14059
rect 9732 14028 10057 14056
rect 9732 14016 9738 14028
rect 10045 14025 10057 14028
rect 10091 14025 10103 14059
rect 10045 14019 10103 14025
rect 10410 14016 10416 14068
rect 10468 14016 10474 14068
rect 12986 14056 12992 14068
rect 12268 14028 12992 14056
rect 8772 13960 8878 13988
rect 7653 13951 7711 13957
rect 12066 13948 12072 14000
rect 12124 13988 12130 14000
rect 12124 13960 12204 13988
rect 12124 13948 12130 13960
rect 5626 13920 5632 13932
rect 5460 13892 5632 13920
rect 5626 13880 5632 13892
rect 5684 13920 5690 13932
rect 6733 13923 6791 13929
rect 5684 13892 6684 13920
rect 5684 13880 5690 13892
rect 6656 13864 6684 13892
rect 6733 13889 6745 13923
rect 6779 13920 6791 13923
rect 7466 13920 7472 13932
rect 6779 13892 7472 13920
rect 6779 13889 6791 13892
rect 6733 13883 6791 13889
rect 7466 13880 7472 13892
rect 7524 13880 7530 13932
rect 7561 13923 7619 13929
rect 7561 13889 7573 13923
rect 7607 13920 7619 13923
rect 7607 13892 8064 13920
rect 7607 13889 7619 13892
rect 7561 13883 7619 13889
rect 4706 13852 4712 13864
rect 4172 13824 4712 13852
rect 4065 13815 4123 13821
rect 4080 13716 4108 13815
rect 4706 13812 4712 13824
rect 4764 13812 4770 13864
rect 6638 13812 6644 13864
rect 6696 13812 6702 13864
rect 7009 13855 7067 13861
rect 7009 13821 7021 13855
rect 7055 13852 7067 13855
rect 7742 13852 7748 13864
rect 7055 13824 7748 13852
rect 7055 13821 7067 13824
rect 7009 13815 7067 13821
rect 5350 13744 5356 13796
rect 5408 13784 5414 13796
rect 6914 13784 6920 13796
rect 5408 13756 6920 13784
rect 5408 13744 5414 13756
rect 6914 13744 6920 13756
rect 6972 13784 6978 13796
rect 7024 13784 7052 13815
rect 7742 13812 7748 13824
rect 7800 13812 7806 13864
rect 8036 13852 8064 13892
rect 8110 13880 8116 13932
rect 8168 13880 8174 13932
rect 11698 13880 11704 13932
rect 11756 13920 11762 13932
rect 12176 13929 12204 13960
rect 11885 13923 11943 13929
rect 11885 13920 11897 13923
rect 11756 13892 11897 13920
rect 11756 13880 11762 13892
rect 11885 13889 11897 13892
rect 11931 13889 11943 13923
rect 11885 13883 11943 13889
rect 12161 13923 12219 13929
rect 12161 13889 12173 13923
rect 12207 13889 12219 13923
rect 12161 13883 12219 13889
rect 8386 13852 8392 13864
rect 8036 13824 8392 13852
rect 8386 13812 8392 13824
rect 8444 13812 8450 13864
rect 8478 13812 8484 13864
rect 8536 13812 8542 13864
rect 10502 13852 10508 13864
rect 9692 13824 10508 13852
rect 6972 13756 7052 13784
rect 6972 13744 6978 13756
rect 4890 13716 4896 13728
rect 4080 13688 4896 13716
rect 4890 13676 4896 13688
rect 4948 13676 4954 13728
rect 6365 13719 6423 13725
rect 6365 13685 6377 13719
rect 6411 13716 6423 13719
rect 6730 13716 6736 13728
rect 6411 13688 6736 13716
rect 6411 13685 6423 13688
rect 6365 13679 6423 13685
rect 6730 13676 6736 13688
rect 6788 13676 6794 13728
rect 7190 13676 7196 13728
rect 7248 13676 7254 13728
rect 7466 13676 7472 13728
rect 7524 13716 7530 13728
rect 9692 13716 9720 13824
rect 10502 13812 10508 13824
rect 10560 13812 10566 13864
rect 10689 13855 10747 13861
rect 10689 13821 10701 13855
rect 10735 13821 10747 13855
rect 10689 13815 10747 13821
rect 11977 13855 12035 13861
rect 11977 13821 11989 13855
rect 12023 13821 12035 13855
rect 11977 13815 12035 13821
rect 10594 13744 10600 13796
rect 10652 13784 10658 13796
rect 10704 13784 10732 13815
rect 10652 13756 10732 13784
rect 10652 13744 10658 13756
rect 11330 13744 11336 13796
rect 11388 13784 11394 13796
rect 11992 13784 12020 13815
rect 12066 13812 12072 13864
rect 12124 13852 12130 13864
rect 12268 13852 12296 14028
rect 12986 14016 12992 14028
rect 13044 14016 13050 14068
rect 13718 14059 13776 14065
rect 13718 14025 13730 14059
rect 13764 14056 13776 14059
rect 15470 14056 15476 14068
rect 13764 14028 15476 14056
rect 13764 14025 13776 14028
rect 13718 14019 13776 14025
rect 15470 14016 15476 14028
rect 15528 14016 15534 14068
rect 17497 14059 17555 14065
rect 17497 14025 17509 14059
rect 17543 14056 17555 14059
rect 18690 14056 18696 14068
rect 17543 14028 18696 14056
rect 17543 14025 17555 14028
rect 17497 14019 17555 14025
rect 18690 14016 18696 14028
rect 18748 14016 18754 14068
rect 21450 14016 21456 14068
rect 21508 14056 21514 14068
rect 22833 14059 22891 14065
rect 22833 14056 22845 14059
rect 21508 14028 22845 14056
rect 21508 14016 21514 14028
rect 22833 14025 22845 14028
rect 22879 14025 22891 14059
rect 22833 14019 22891 14025
rect 22922 14016 22928 14068
rect 22980 14056 22986 14068
rect 23474 14056 23480 14068
rect 22980 14028 23480 14056
rect 22980 14016 22986 14028
rect 23474 14016 23480 14028
rect 23532 14016 23538 14068
rect 12710 13948 12716 14000
rect 12768 13988 12774 14000
rect 13817 13991 13875 13997
rect 13817 13988 13829 13991
rect 12768 13960 13829 13988
rect 12768 13948 12774 13960
rect 13817 13957 13829 13960
rect 13863 13988 13875 13991
rect 14274 13988 14280 14000
rect 13863 13960 14280 13988
rect 13863 13957 13875 13960
rect 13817 13951 13875 13957
rect 14274 13948 14280 13960
rect 14332 13948 14338 14000
rect 20990 13948 20996 14000
rect 21048 13988 21054 14000
rect 23382 13988 23388 14000
rect 21048 13960 22508 13988
rect 21048 13948 21054 13960
rect 12621 13923 12679 13929
rect 12621 13920 12633 13923
rect 12360 13892 12633 13920
rect 12360 13861 12388 13892
rect 12621 13889 12633 13892
rect 12667 13889 12679 13923
rect 13532 13913 13590 13919
rect 13532 13910 13544 13913
rect 12621 13883 12679 13889
rect 13464 13882 13544 13910
rect 12124 13824 12296 13852
rect 12345 13855 12403 13861
rect 12124 13812 12130 13824
rect 12345 13821 12357 13855
rect 12391 13821 12403 13855
rect 12345 13815 12403 13821
rect 12713 13855 12771 13861
rect 12713 13821 12725 13855
rect 12759 13852 12771 13855
rect 13262 13852 13268 13864
rect 12759 13824 13268 13852
rect 12759 13821 12771 13824
rect 12713 13815 12771 13821
rect 13262 13812 13268 13824
rect 13320 13812 13326 13864
rect 12802 13784 12808 13796
rect 11388 13756 12808 13784
rect 11388 13744 11394 13756
rect 12802 13744 12808 13756
rect 12860 13744 12866 13796
rect 12989 13787 13047 13793
rect 12989 13753 13001 13787
rect 13035 13784 13047 13787
rect 13354 13784 13360 13796
rect 13035 13756 13360 13784
rect 13035 13753 13047 13756
rect 12989 13747 13047 13753
rect 13354 13744 13360 13756
rect 13412 13744 13418 13796
rect 13464 13784 13492 13882
rect 13532 13879 13544 13882
rect 13578 13879 13590 13913
rect 13630 13880 13636 13932
rect 13688 13880 13694 13932
rect 17034 13880 17040 13932
rect 17092 13920 17098 13932
rect 17313 13923 17371 13929
rect 17313 13920 17325 13923
rect 17092 13892 17325 13920
rect 17092 13880 17098 13892
rect 17313 13889 17325 13892
rect 17359 13889 17371 13923
rect 17313 13883 17371 13889
rect 17494 13880 17500 13932
rect 17552 13880 17558 13932
rect 21910 13880 21916 13932
rect 21968 13920 21974 13932
rect 22005 13923 22063 13929
rect 22005 13920 22017 13923
rect 21968 13892 22017 13920
rect 21968 13880 21974 13892
rect 22005 13889 22017 13892
rect 22051 13889 22063 13923
rect 22005 13883 22063 13889
rect 22186 13880 22192 13932
rect 22244 13880 22250 13932
rect 22480 13929 22508 13960
rect 22572 13960 23388 13988
rect 22572 13929 22600 13960
rect 23382 13948 23388 13960
rect 23440 13948 23446 14000
rect 22465 13923 22523 13929
rect 22465 13889 22477 13923
rect 22511 13889 22523 13923
rect 22465 13883 22523 13889
rect 22557 13923 22615 13929
rect 22557 13889 22569 13923
rect 22603 13889 22615 13923
rect 22557 13883 22615 13889
rect 22646 13880 22652 13932
rect 22704 13920 22710 13932
rect 23109 13923 23167 13929
rect 23109 13920 23121 13923
rect 22704 13892 23121 13920
rect 22704 13880 22710 13892
rect 23109 13889 23121 13892
rect 23155 13920 23167 13923
rect 23290 13920 23296 13932
rect 23155 13892 23296 13920
rect 23155 13889 23167 13892
rect 23109 13883 23167 13889
rect 23290 13880 23296 13892
rect 23348 13880 23354 13932
rect 13532 13873 13590 13879
rect 17862 13812 17868 13864
rect 17920 13812 17926 13864
rect 22738 13812 22744 13864
rect 22796 13812 22802 13864
rect 22833 13855 22891 13861
rect 22833 13821 22845 13855
rect 22879 13852 22891 13855
rect 22922 13852 22928 13864
rect 22879 13824 22928 13852
rect 22879 13821 22891 13824
rect 22833 13815 22891 13821
rect 22922 13812 22928 13824
rect 22980 13852 22986 13864
rect 23658 13852 23664 13864
rect 22980 13824 23664 13852
rect 22980 13812 22986 13824
rect 23658 13812 23664 13824
rect 23716 13812 23722 13864
rect 13814 13784 13820 13796
rect 13464 13756 13820 13784
rect 13814 13744 13820 13756
rect 13872 13744 13878 13796
rect 18046 13744 18052 13796
rect 18104 13784 18110 13796
rect 18141 13787 18199 13793
rect 18141 13784 18153 13787
rect 18104 13756 18153 13784
rect 18104 13744 18110 13756
rect 18141 13753 18153 13756
rect 18187 13753 18199 13787
rect 18141 13747 18199 13753
rect 22462 13744 22468 13796
rect 22520 13784 22526 13796
rect 23017 13787 23075 13793
rect 23017 13784 23029 13787
rect 22520 13756 23029 13784
rect 22520 13744 22526 13756
rect 23017 13753 23029 13756
rect 23063 13753 23075 13787
rect 23017 13747 23075 13753
rect 7524 13688 9720 13716
rect 7524 13676 7530 13688
rect 9858 13676 9864 13728
rect 9916 13725 9922 13728
rect 9916 13719 9965 13725
rect 9916 13685 9919 13719
rect 9953 13716 9965 13719
rect 11348 13716 11376 13744
rect 9953 13688 11376 13716
rect 9953 13685 9965 13688
rect 9916 13679 9965 13685
rect 9916 13676 9922 13679
rect 18322 13676 18328 13728
rect 18380 13676 18386 13728
rect 22189 13719 22247 13725
rect 22189 13685 22201 13719
rect 22235 13716 22247 13719
rect 22278 13716 22284 13728
rect 22235 13688 22284 13716
rect 22235 13685 22247 13688
rect 22189 13679 22247 13685
rect 22278 13676 22284 13688
rect 22336 13676 22342 13728
rect 22373 13719 22431 13725
rect 22373 13685 22385 13719
rect 22419 13716 22431 13719
rect 22554 13716 22560 13728
rect 22419 13688 22560 13716
rect 22419 13685 22431 13688
rect 22373 13679 22431 13685
rect 22554 13676 22560 13688
rect 22612 13676 22618 13728
rect 22649 13719 22707 13725
rect 22649 13685 22661 13719
rect 22695 13716 22707 13719
rect 22830 13716 22836 13728
rect 22695 13688 22836 13716
rect 22695 13685 22707 13688
rect 22649 13679 22707 13685
rect 22830 13676 22836 13688
rect 22888 13676 22894 13728
rect 1104 13626 25208 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 25208 13626
rect 1104 13552 25208 13574
rect 2314 13472 2320 13524
rect 2372 13512 2378 13524
rect 2777 13515 2835 13521
rect 2777 13512 2789 13515
rect 2372 13484 2789 13512
rect 2372 13472 2378 13484
rect 2777 13481 2789 13484
rect 2823 13481 2835 13515
rect 2777 13475 2835 13481
rect 8478 13472 8484 13524
rect 8536 13512 8542 13524
rect 8941 13515 8999 13521
rect 8941 13512 8953 13515
rect 8536 13484 8953 13512
rect 8536 13472 8542 13484
rect 8941 13481 8953 13484
rect 8987 13481 8999 13515
rect 8941 13475 8999 13481
rect 11698 13472 11704 13524
rect 11756 13512 11762 13524
rect 12069 13515 12127 13521
rect 12069 13512 12081 13515
rect 11756 13484 12081 13512
rect 11756 13472 11762 13484
rect 12069 13481 12081 13484
rect 12115 13481 12127 13515
rect 12069 13475 12127 13481
rect 14090 13472 14096 13524
rect 14148 13512 14154 13524
rect 14277 13515 14335 13521
rect 14277 13512 14289 13515
rect 14148 13484 14289 13512
rect 14148 13472 14154 13484
rect 14277 13481 14289 13484
rect 14323 13481 14335 13515
rect 14277 13475 14335 13481
rect 16298 13472 16304 13524
rect 16356 13512 16362 13524
rect 18506 13512 18512 13524
rect 16356 13484 18512 13512
rect 16356 13472 16362 13484
rect 18506 13472 18512 13484
rect 18564 13472 18570 13524
rect 21821 13515 21879 13521
rect 21821 13481 21833 13515
rect 21867 13512 21879 13515
rect 21910 13512 21916 13524
rect 21867 13484 21916 13512
rect 21867 13481 21879 13484
rect 21821 13475 21879 13481
rect 21910 13472 21916 13484
rect 21968 13472 21974 13524
rect 22278 13472 22284 13524
rect 22336 13512 22342 13524
rect 22373 13515 22431 13521
rect 22373 13512 22385 13515
rect 22336 13484 22385 13512
rect 22336 13472 22342 13484
rect 22373 13481 22385 13484
rect 22419 13481 22431 13515
rect 22373 13475 22431 13481
rect 22462 13472 22468 13524
rect 22520 13512 22526 13524
rect 22557 13515 22615 13521
rect 22557 13512 22569 13515
rect 22520 13484 22569 13512
rect 22520 13472 22526 13484
rect 22557 13481 22569 13484
rect 22603 13481 22615 13515
rect 22557 13475 22615 13481
rect 22925 13515 22983 13521
rect 22925 13481 22937 13515
rect 22971 13512 22983 13515
rect 23014 13512 23020 13524
rect 22971 13484 23020 13512
rect 22971 13481 22983 13484
rect 22925 13475 22983 13481
rect 3142 13404 3148 13456
rect 3200 13444 3206 13456
rect 3200 13416 3372 13444
rect 3200 13404 3206 13416
rect 3234 13336 3240 13388
rect 3292 13336 3298 13388
rect 3344 13385 3372 13416
rect 8386 13404 8392 13456
rect 8444 13444 8450 13456
rect 8619 13447 8677 13453
rect 8619 13444 8631 13447
rect 8444 13416 8631 13444
rect 8444 13404 8450 13416
rect 8619 13413 8631 13416
rect 8665 13444 8677 13447
rect 11517 13447 11575 13453
rect 8665 13416 9444 13444
rect 8665 13413 8677 13416
rect 8619 13407 8677 13413
rect 9416 13388 9444 13416
rect 11517 13413 11529 13447
rect 11563 13444 11575 13447
rect 11790 13444 11796 13456
rect 11563 13416 11796 13444
rect 11563 13413 11575 13416
rect 11517 13407 11575 13413
rect 11790 13404 11796 13416
rect 11848 13404 11854 13456
rect 17402 13404 17408 13456
rect 17460 13404 17466 13456
rect 17770 13404 17776 13456
rect 17828 13444 17834 13456
rect 17828 13416 18828 13444
rect 17828 13404 17834 13416
rect 3329 13379 3387 13385
rect 3329 13345 3341 13379
rect 3375 13345 3387 13379
rect 3329 13339 3387 13345
rect 4614 13336 4620 13388
rect 4672 13376 4678 13388
rect 4890 13376 4896 13388
rect 4672 13348 4896 13376
rect 4672 13336 4678 13348
rect 4890 13336 4896 13348
rect 4948 13336 4954 13388
rect 5261 13379 5319 13385
rect 5261 13345 5273 13379
rect 5307 13376 5319 13379
rect 5534 13376 5540 13388
rect 5307 13348 5540 13376
rect 5307 13345 5319 13348
rect 5261 13339 5319 13345
rect 5534 13336 5540 13348
rect 5592 13336 5598 13388
rect 6822 13336 6828 13388
rect 6880 13336 6886 13388
rect 7190 13336 7196 13388
rect 7248 13336 7254 13388
rect 9398 13336 9404 13388
rect 9456 13336 9462 13388
rect 9585 13379 9643 13385
rect 9585 13345 9597 13379
rect 9631 13376 9643 13379
rect 9766 13376 9772 13388
rect 9631 13348 9772 13376
rect 9631 13345 9643 13348
rect 9585 13339 9643 13345
rect 9766 13336 9772 13348
rect 9824 13376 9830 13388
rect 10594 13376 10600 13388
rect 9824 13348 10600 13376
rect 9824 13336 9830 13348
rect 10594 13336 10600 13348
rect 10652 13336 10658 13388
rect 17420 13376 17448 13404
rect 17957 13379 18015 13385
rect 17957 13376 17969 13379
rect 16224 13348 17264 13376
rect 17420 13348 17969 13376
rect 16224 13320 16252 13348
rect 3145 13311 3203 13317
rect 3145 13277 3157 13311
rect 3191 13308 3203 13311
rect 4706 13308 4712 13320
rect 3191 13280 4712 13308
rect 3191 13277 3203 13280
rect 3145 13271 3203 13277
rect 4706 13268 4712 13280
rect 4764 13268 4770 13320
rect 6638 13308 6644 13320
rect 6288 13280 6644 13308
rect 6288 13226 6316 13280
rect 6638 13268 6644 13280
rect 6696 13268 6702 13320
rect 11422 13268 11428 13320
rect 11480 13308 11486 13320
rect 11793 13311 11851 13317
rect 11793 13308 11805 13311
rect 11480 13280 11805 13308
rect 11480 13268 11486 13280
rect 11793 13277 11805 13280
rect 11839 13277 11851 13311
rect 15286 13308 15292 13320
rect 11793 13271 11851 13277
rect 14384 13280 15292 13308
rect 8202 13200 8208 13252
rect 8260 13200 8266 13252
rect 11514 13200 11520 13252
rect 11572 13240 11578 13252
rect 11885 13243 11943 13249
rect 11885 13240 11897 13243
rect 11572 13212 11897 13240
rect 11572 13200 11578 13212
rect 11885 13209 11897 13212
rect 11931 13209 11943 13243
rect 11885 13203 11943 13209
rect 13078 13200 13084 13252
rect 13136 13240 13142 13252
rect 14093 13243 14151 13249
rect 14093 13240 14105 13243
rect 13136 13212 14105 13240
rect 13136 13200 13142 13212
rect 14093 13209 14105 13212
rect 14139 13209 14151 13243
rect 14093 13203 14151 13209
rect 14298 13243 14356 13249
rect 14298 13209 14310 13243
rect 14344 13240 14356 13243
rect 14384 13240 14412 13280
rect 15286 13268 15292 13280
rect 15344 13268 15350 13320
rect 15746 13268 15752 13320
rect 15804 13268 15810 13320
rect 16022 13268 16028 13320
rect 16080 13308 16086 13320
rect 16206 13308 16212 13320
rect 16080 13280 16212 13308
rect 16080 13268 16086 13280
rect 16206 13268 16212 13280
rect 16264 13268 16270 13320
rect 16758 13268 16764 13320
rect 16816 13268 16822 13320
rect 17129 13311 17187 13317
rect 17129 13277 17141 13311
rect 17175 13277 17187 13311
rect 17236 13308 17264 13348
rect 17957 13345 17969 13348
rect 18003 13345 18015 13379
rect 17957 13339 18015 13345
rect 17405 13311 17463 13317
rect 17405 13308 17417 13311
rect 17236 13280 17417 13308
rect 17129 13271 17187 13277
rect 17405 13277 17417 13280
rect 17451 13277 17463 13311
rect 17405 13271 17463 13277
rect 17144 13240 17172 13271
rect 17678 13268 17684 13320
rect 17736 13268 17742 13320
rect 17770 13268 17776 13320
rect 17828 13268 17834 13320
rect 17865 13311 17923 13317
rect 17865 13277 17877 13311
rect 17911 13277 17923 13311
rect 17972 13308 18000 13339
rect 18046 13336 18052 13388
rect 18104 13376 18110 13388
rect 18693 13379 18751 13385
rect 18693 13376 18705 13379
rect 18104 13348 18705 13376
rect 18104 13336 18110 13348
rect 18693 13345 18705 13348
rect 18739 13345 18751 13379
rect 18693 13339 18751 13345
rect 18233 13311 18291 13317
rect 18233 13308 18245 13311
rect 17972 13280 18245 13308
rect 17865 13271 17923 13277
rect 18233 13277 18245 13280
rect 18279 13277 18291 13311
rect 18233 13271 18291 13277
rect 18509 13311 18567 13317
rect 18509 13277 18521 13311
rect 18555 13308 18567 13311
rect 18800 13308 18828 13416
rect 21266 13404 21272 13456
rect 21324 13404 21330 13456
rect 22005 13447 22063 13453
rect 22005 13413 22017 13447
rect 22051 13444 22063 13447
rect 22094 13444 22100 13456
rect 22051 13416 22100 13444
rect 22051 13413 22063 13416
rect 22005 13407 22063 13413
rect 22094 13404 22100 13416
rect 22152 13404 22158 13456
rect 22572 13444 22600 13475
rect 23014 13472 23020 13484
rect 23072 13472 23078 13524
rect 23109 13515 23167 13521
rect 23109 13481 23121 13515
rect 23155 13512 23167 13515
rect 23198 13512 23204 13524
rect 23155 13484 23204 13512
rect 23155 13481 23167 13484
rect 23109 13475 23167 13481
rect 23198 13472 23204 13484
rect 23256 13472 23262 13524
rect 23658 13472 23664 13524
rect 23716 13472 23722 13524
rect 22572 13416 22968 13444
rect 22841 13321 22899 13327
rect 18555 13280 18828 13308
rect 18555 13277 18567 13280
rect 18509 13271 18567 13277
rect 14344 13212 14412 13240
rect 14476 13212 17172 13240
rect 14344 13209 14356 13212
rect 14298 13203 14356 13209
rect 6546 13132 6552 13184
rect 6604 13172 6610 13184
rect 6687 13175 6745 13181
rect 6687 13172 6699 13175
rect 6604 13144 6699 13172
rect 6604 13132 6610 13144
rect 6687 13141 6699 13144
rect 6733 13141 6745 13175
rect 6687 13135 6745 13141
rect 9309 13175 9367 13181
rect 9309 13141 9321 13175
rect 9355 13172 9367 13175
rect 9858 13172 9864 13184
rect 9355 13144 9864 13172
rect 9355 13141 9367 13144
rect 9309 13135 9367 13141
rect 9858 13132 9864 13144
rect 9916 13132 9922 13184
rect 11606 13132 11612 13184
rect 11664 13172 11670 13184
rect 14476 13181 14504 13212
rect 17218 13200 17224 13252
rect 17276 13240 17282 13252
rect 17586 13240 17592 13252
rect 17276 13212 17592 13240
rect 17276 13200 17282 13212
rect 17586 13200 17592 13212
rect 17644 13240 17650 13252
rect 17788 13240 17816 13268
rect 17644 13212 17816 13240
rect 17880 13240 17908 13271
rect 20990 13268 20996 13320
rect 21048 13268 21054 13320
rect 21082 13268 21088 13320
rect 21140 13268 21146 13320
rect 21269 13311 21327 13317
rect 21269 13277 21281 13311
rect 21315 13308 21327 13311
rect 21450 13308 21456 13320
rect 21315 13280 21456 13308
rect 21315 13277 21327 13280
rect 21269 13271 21327 13277
rect 21450 13268 21456 13280
rect 21508 13268 21514 13320
rect 21542 13268 21548 13320
rect 21600 13268 21606 13320
rect 21729 13311 21787 13317
rect 21729 13277 21741 13311
rect 21775 13308 21787 13311
rect 22002 13308 22008 13320
rect 21775 13280 22008 13308
rect 21775 13277 21787 13280
rect 21729 13271 21787 13277
rect 22002 13268 22008 13280
rect 22060 13308 22066 13320
rect 22281 13311 22339 13317
rect 22281 13308 22293 13311
rect 22060 13280 22293 13308
rect 22060 13268 22066 13280
rect 22281 13277 22293 13280
rect 22327 13308 22339 13311
rect 22370 13308 22376 13320
rect 22327 13280 22376 13308
rect 22327 13277 22339 13280
rect 22281 13271 22339 13277
rect 22370 13268 22376 13280
rect 22428 13268 22434 13320
rect 22841 13287 22853 13321
rect 22887 13318 22899 13321
rect 22940 13318 22968 13416
rect 23106 13336 23112 13388
rect 23164 13376 23170 13388
rect 23385 13379 23443 13385
rect 23385 13376 23397 13379
rect 23164 13348 23397 13376
rect 23164 13336 23170 13348
rect 23385 13345 23397 13348
rect 23431 13376 23443 13379
rect 24486 13376 24492 13388
rect 23431 13348 24492 13376
rect 23431 13345 23443 13348
rect 23385 13339 23443 13345
rect 22887 13290 22968 13318
rect 23017 13311 23075 13317
rect 22887 13287 22899 13290
rect 22841 13281 22899 13287
rect 23017 13277 23029 13311
rect 23063 13308 23075 13311
rect 23198 13308 23204 13320
rect 23063 13280 23204 13308
rect 23063 13277 23075 13280
rect 23017 13271 23075 13277
rect 23198 13268 23204 13280
rect 23256 13268 23262 13320
rect 23290 13268 23296 13320
rect 23348 13268 23354 13320
rect 23474 13268 23480 13320
rect 23532 13308 23538 13320
rect 23860 13317 23888 13348
rect 24486 13336 24492 13348
rect 24544 13336 24550 13388
rect 23661 13311 23719 13317
rect 23661 13308 23673 13311
rect 23532 13280 23673 13308
rect 23532 13268 23538 13280
rect 23661 13277 23673 13280
rect 23707 13277 23719 13311
rect 23661 13271 23719 13277
rect 23845 13311 23903 13317
rect 23845 13277 23857 13311
rect 23891 13277 23903 13311
rect 23845 13271 23903 13277
rect 23937 13311 23995 13317
rect 23937 13277 23949 13311
rect 23983 13277 23995 13311
rect 23937 13271 23995 13277
rect 22541 13243 22599 13249
rect 22541 13240 22553 13243
rect 17880 13212 18368 13240
rect 17644 13200 17650 13212
rect 11701 13175 11759 13181
rect 11701 13172 11713 13175
rect 11664 13144 11713 13172
rect 11664 13132 11670 13144
rect 11701 13141 11713 13144
rect 11747 13141 11759 13175
rect 11701 13135 11759 13141
rect 14461 13175 14519 13181
rect 14461 13141 14473 13175
rect 14507 13141 14519 13175
rect 14461 13135 14519 13141
rect 15010 13132 15016 13184
rect 15068 13172 15074 13184
rect 15565 13175 15623 13181
rect 15565 13172 15577 13175
rect 15068 13144 15577 13172
rect 15068 13132 15074 13144
rect 15565 13141 15577 13144
rect 15611 13141 15623 13175
rect 15565 13135 15623 13141
rect 15933 13175 15991 13181
rect 15933 13141 15945 13175
rect 15979 13172 15991 13175
rect 16209 13175 16267 13181
rect 16209 13172 16221 13175
rect 15979 13144 16221 13172
rect 15979 13141 15991 13144
rect 15933 13135 15991 13141
rect 16209 13141 16221 13144
rect 16255 13141 16267 13175
rect 16209 13135 16267 13141
rect 16942 13132 16948 13184
rect 17000 13132 17006 13184
rect 17034 13132 17040 13184
rect 17092 13172 17098 13184
rect 17313 13175 17371 13181
rect 17313 13172 17325 13175
rect 17092 13144 17325 13172
rect 17092 13132 17098 13144
rect 17313 13141 17325 13144
rect 17359 13141 17371 13175
rect 17313 13135 17371 13141
rect 18138 13132 18144 13184
rect 18196 13132 18202 13184
rect 18340 13181 18368 13212
rect 22480 13212 22553 13240
rect 18325 13175 18383 13181
rect 18325 13141 18337 13175
rect 18371 13172 18383 13175
rect 18414 13172 18420 13184
rect 18371 13144 18420 13172
rect 18371 13141 18383 13144
rect 18325 13135 18383 13141
rect 18414 13132 18420 13144
rect 18472 13132 18478 13184
rect 20622 13132 20628 13184
rect 20680 13172 20686 13184
rect 21174 13172 21180 13184
rect 20680 13144 21180 13172
rect 20680 13132 20686 13144
rect 21174 13132 21180 13144
rect 21232 13172 21238 13184
rect 21361 13175 21419 13181
rect 21361 13172 21373 13175
rect 21232 13144 21373 13172
rect 21232 13132 21238 13144
rect 21361 13141 21373 13144
rect 21407 13141 21419 13175
rect 21361 13135 21419 13141
rect 22094 13132 22100 13184
rect 22152 13172 22158 13184
rect 22480 13172 22508 13212
rect 22541 13209 22553 13212
rect 22587 13209 22599 13243
rect 22541 13203 22599 13209
rect 22646 13200 22652 13252
rect 22704 13249 22710 13252
rect 22704 13243 22753 13249
rect 22704 13209 22707 13243
rect 22741 13209 22753 13243
rect 23308 13240 23336 13268
rect 23566 13240 23572 13252
rect 23308 13212 23572 13240
rect 22704 13203 22753 13209
rect 22704 13200 22710 13203
rect 23566 13200 23572 13212
rect 23624 13240 23630 13252
rect 23952 13240 23980 13271
rect 24026 13268 24032 13320
rect 24084 13308 24090 13320
rect 24121 13311 24179 13317
rect 24121 13308 24133 13311
rect 24084 13280 24133 13308
rect 24084 13268 24090 13280
rect 24121 13277 24133 13280
rect 24167 13277 24179 13311
rect 24121 13271 24179 13277
rect 24578 13268 24584 13320
rect 24636 13268 24642 13320
rect 23624 13212 23980 13240
rect 23624 13200 23630 13212
rect 22152 13144 22508 13172
rect 24029 13175 24087 13181
rect 22152 13132 22158 13144
rect 24029 13141 24041 13175
rect 24075 13172 24087 13175
rect 24302 13172 24308 13184
rect 24075 13144 24308 13172
rect 24075 13141 24087 13144
rect 24029 13135 24087 13141
rect 24302 13132 24308 13144
rect 24360 13132 24366 13184
rect 24762 13132 24768 13184
rect 24820 13132 24826 13184
rect 1104 13082 25208 13104
rect 1104 13030 4874 13082
rect 4926 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 25208 13082
rect 1104 13008 25208 13030
rect 3234 12928 3240 12980
rect 3292 12968 3298 12980
rect 3697 12971 3755 12977
rect 3697 12968 3709 12971
rect 3292 12940 3709 12968
rect 3292 12928 3298 12940
rect 3697 12937 3709 12940
rect 3743 12937 3755 12971
rect 3697 12931 3755 12937
rect 5169 12971 5227 12977
rect 5169 12937 5181 12971
rect 5215 12968 5227 12971
rect 6638 12968 6644 12980
rect 5215 12940 6644 12968
rect 5215 12937 5227 12940
rect 5169 12931 5227 12937
rect 6638 12928 6644 12940
rect 6696 12928 6702 12980
rect 7466 12928 7472 12980
rect 7524 12968 7530 12980
rect 8159 12971 8217 12977
rect 8159 12968 8171 12971
rect 7524 12940 8171 12968
rect 7524 12928 7530 12940
rect 8159 12937 8171 12940
rect 8205 12937 8217 12971
rect 8159 12931 8217 12937
rect 16758 12928 16764 12980
rect 16816 12968 16822 12980
rect 16816 12940 17632 12968
rect 16816 12928 16822 12940
rect 4614 12860 4620 12912
rect 4672 12900 4678 12912
rect 4672 12872 6408 12900
rect 4672 12860 4678 12872
rect 3789 12835 3847 12841
rect 3789 12801 3801 12835
rect 3835 12832 3847 12835
rect 6270 12832 6276 12844
rect 3835 12804 6276 12832
rect 3835 12801 3847 12804
rect 3789 12795 3847 12801
rect 6270 12792 6276 12804
rect 6328 12792 6334 12844
rect 6380 12841 6408 12872
rect 7098 12860 7104 12912
rect 7156 12860 7162 12912
rect 16298 12900 16304 12912
rect 16054 12872 16304 12900
rect 16298 12860 16304 12872
rect 16356 12860 16362 12912
rect 17126 12860 17132 12912
rect 17184 12900 17190 12912
rect 17494 12900 17500 12912
rect 17184 12872 17500 12900
rect 17184 12860 17190 12872
rect 17494 12860 17500 12872
rect 17552 12860 17558 12912
rect 17604 12909 17632 12940
rect 18690 12928 18696 12980
rect 18748 12968 18754 12980
rect 18748 12940 19656 12968
rect 18748 12928 18754 12940
rect 17589 12903 17647 12909
rect 17589 12869 17601 12903
rect 17635 12869 17647 12903
rect 17589 12863 17647 12869
rect 6365 12835 6423 12841
rect 6365 12801 6377 12835
rect 6411 12801 6423 12835
rect 6365 12795 6423 12801
rect 6730 12792 6736 12844
rect 6788 12792 6794 12844
rect 9493 12835 9551 12841
rect 9493 12801 9505 12835
rect 9539 12832 9551 12835
rect 10686 12832 10692 12844
rect 9539 12804 10692 12832
rect 9539 12801 9551 12804
rect 9493 12795 9551 12801
rect 10686 12792 10692 12804
rect 10744 12832 10750 12844
rect 12066 12832 12072 12844
rect 10744 12804 12072 12832
rect 10744 12792 10750 12804
rect 12066 12792 12072 12804
rect 12124 12792 12130 12844
rect 12253 12835 12311 12841
rect 12253 12801 12265 12835
rect 12299 12832 12311 12835
rect 13814 12832 13820 12844
rect 12299 12804 13820 12832
rect 12299 12801 12311 12804
rect 12253 12795 12311 12801
rect 13814 12792 13820 12804
rect 13872 12792 13878 12844
rect 15010 12792 15016 12844
rect 15068 12792 15074 12844
rect 16439 12835 16497 12841
rect 16439 12801 16451 12835
rect 16485 12832 16497 12835
rect 16669 12835 16727 12841
rect 16669 12832 16681 12835
rect 16485 12804 16681 12832
rect 16485 12801 16497 12804
rect 16439 12795 16497 12801
rect 16669 12801 16681 12804
rect 16715 12832 16727 12835
rect 16758 12832 16764 12844
rect 16715 12804 16764 12832
rect 16715 12801 16727 12804
rect 16669 12795 16727 12801
rect 16758 12792 16764 12804
rect 16816 12792 16822 12844
rect 16853 12835 16911 12841
rect 16853 12801 16865 12835
rect 16899 12801 16911 12835
rect 16853 12795 16911 12801
rect 16945 12835 17003 12841
rect 16945 12801 16957 12835
rect 16991 12832 17003 12835
rect 17034 12832 17040 12844
rect 16991 12804 17040 12832
rect 16991 12801 17003 12804
rect 16945 12795 17003 12801
rect 3605 12767 3663 12773
rect 3605 12733 3617 12767
rect 3651 12733 3663 12767
rect 3605 12727 3663 12733
rect 2314 12656 2320 12708
rect 2372 12696 2378 12708
rect 3620 12696 3648 12727
rect 4706 12724 4712 12776
rect 4764 12764 4770 12776
rect 5261 12767 5319 12773
rect 5261 12764 5273 12767
rect 4764 12736 5273 12764
rect 4764 12724 4770 12736
rect 5261 12733 5273 12736
rect 5307 12733 5319 12767
rect 5261 12727 5319 12733
rect 5350 12724 5356 12776
rect 5408 12764 5414 12776
rect 5408 12736 5488 12764
rect 5408 12724 5414 12736
rect 5460 12696 5488 12736
rect 9582 12724 9588 12776
rect 9640 12724 9646 12776
rect 9766 12724 9772 12776
rect 9824 12724 9830 12776
rect 14642 12724 14648 12776
rect 14700 12724 14706 12776
rect 16868 12764 16896 12795
rect 17034 12792 17040 12804
rect 17092 12792 17098 12844
rect 17218 12792 17224 12844
rect 17276 12792 17282 12844
rect 17313 12835 17371 12841
rect 17313 12801 17325 12835
rect 17359 12832 17371 12835
rect 17604 12832 17632 12863
rect 17678 12860 17684 12912
rect 17736 12900 17742 12912
rect 19628 12909 19656 12940
rect 21358 12928 21364 12980
rect 21416 12928 21422 12980
rect 21450 12928 21456 12980
rect 21508 12968 21514 12980
rect 21545 12971 21603 12977
rect 21545 12968 21557 12971
rect 21508 12940 21557 12968
rect 21508 12928 21514 12940
rect 21545 12937 21557 12940
rect 21591 12937 21603 12971
rect 21545 12931 21603 12937
rect 21634 12928 21640 12980
rect 21692 12968 21698 12980
rect 21821 12971 21879 12977
rect 21821 12968 21833 12971
rect 21692 12940 21833 12968
rect 21692 12928 21698 12940
rect 21821 12937 21833 12940
rect 21867 12937 21879 12971
rect 21821 12931 21879 12937
rect 21928 12940 22140 12968
rect 19521 12903 19579 12909
rect 19521 12900 19533 12903
rect 17736 12872 18276 12900
rect 17736 12860 17742 12872
rect 18248 12841 18276 12872
rect 18616 12872 19533 12900
rect 17359 12804 17632 12832
rect 17773 12835 17831 12841
rect 17359 12801 17371 12804
rect 17313 12795 17371 12801
rect 17773 12801 17785 12835
rect 17819 12801 17831 12835
rect 17773 12795 17831 12801
rect 18233 12835 18291 12841
rect 18233 12801 18245 12835
rect 18279 12801 18291 12835
rect 18233 12795 18291 12801
rect 17236 12764 17264 12792
rect 17788 12764 17816 12795
rect 16868 12736 17816 12764
rect 18322 12724 18328 12776
rect 18380 12724 18386 12776
rect 18616 12773 18644 12872
rect 19521 12869 19533 12872
rect 19567 12869 19579 12903
rect 19521 12863 19579 12869
rect 19613 12903 19671 12909
rect 19613 12869 19625 12903
rect 19659 12869 19671 12903
rect 21928 12900 21956 12940
rect 19613 12863 19671 12869
rect 21192 12872 21956 12900
rect 22112 12900 22140 12940
rect 22462 12928 22468 12980
rect 22520 12928 22526 12980
rect 24121 12971 24179 12977
rect 24121 12968 24133 12971
rect 22756 12940 24133 12968
rect 22649 12903 22707 12909
rect 22649 12900 22661 12903
rect 22112 12872 22661 12900
rect 18690 12792 18696 12844
rect 18748 12832 18754 12844
rect 18877 12835 18935 12841
rect 18877 12832 18889 12835
rect 18748 12804 18889 12832
rect 18748 12792 18754 12804
rect 18877 12801 18889 12804
rect 18923 12801 18935 12835
rect 18877 12795 18935 12801
rect 19337 12835 19395 12841
rect 19337 12801 19349 12835
rect 19383 12801 19395 12835
rect 19337 12795 19395 12801
rect 18601 12767 18659 12773
rect 18601 12733 18613 12767
rect 18647 12733 18659 12767
rect 18601 12727 18659 12733
rect 18782 12724 18788 12776
rect 18840 12724 18846 12776
rect 19352 12764 19380 12795
rect 19702 12792 19708 12844
rect 19760 12792 19766 12844
rect 21192 12841 21220 12872
rect 22649 12869 22661 12872
rect 22695 12869 22707 12903
rect 22649 12863 22707 12869
rect 21177 12835 21235 12841
rect 21177 12801 21189 12835
rect 21223 12801 21235 12835
rect 21637 12835 21695 12841
rect 21637 12832 21649 12835
rect 21177 12795 21235 12801
rect 21376 12804 21649 12832
rect 20898 12764 20904 12776
rect 19352 12736 20904 12764
rect 20898 12724 20904 12736
rect 20956 12724 20962 12776
rect 21082 12724 21088 12776
rect 21140 12764 21146 12776
rect 21269 12767 21327 12773
rect 21269 12764 21281 12767
rect 21140 12736 21281 12764
rect 21140 12724 21146 12736
rect 21269 12733 21281 12736
rect 21315 12733 21327 12767
rect 21269 12727 21327 12733
rect 2372 12668 5488 12696
rect 16761 12699 16819 12705
rect 2372 12656 2378 12668
rect 16761 12665 16773 12699
rect 16807 12696 16819 12699
rect 18230 12696 18236 12708
rect 16807 12668 18236 12696
rect 16807 12665 16819 12668
rect 16761 12659 16819 12665
rect 18230 12656 18236 12668
rect 18288 12656 18294 12708
rect 19245 12699 19303 12705
rect 19245 12665 19257 12699
rect 19291 12696 19303 12699
rect 21376 12696 21404 12804
rect 21637 12801 21649 12804
rect 21683 12801 21695 12835
rect 21637 12795 21695 12801
rect 22554 12792 22560 12844
rect 22612 12830 22618 12844
rect 22756 12832 22784 12940
rect 24121 12937 24133 12940
rect 24167 12937 24179 12971
rect 24121 12931 24179 12937
rect 23474 12860 23480 12912
rect 23532 12900 23538 12912
rect 23569 12903 23627 12909
rect 23569 12900 23581 12903
rect 23532 12872 23581 12900
rect 23532 12860 23538 12872
rect 23569 12869 23581 12872
rect 23615 12900 23627 12903
rect 24026 12900 24032 12912
rect 23615 12872 24032 12900
rect 23615 12869 23627 12872
rect 23569 12863 23627 12869
rect 24026 12860 24032 12872
rect 24084 12860 24090 12912
rect 24397 12903 24455 12909
rect 24397 12900 24409 12903
rect 24228 12872 24409 12900
rect 22664 12830 22784 12832
rect 22612 12804 22784 12830
rect 22612 12802 22692 12804
rect 22612 12792 22618 12802
rect 22830 12792 22836 12844
rect 22888 12832 22894 12844
rect 23014 12832 23020 12844
rect 22888 12804 23020 12832
rect 22888 12792 22894 12804
rect 23014 12792 23020 12804
rect 23072 12792 23078 12844
rect 23106 12792 23112 12844
rect 23164 12792 23170 12844
rect 23293 12835 23351 12841
rect 23293 12801 23305 12835
rect 23339 12801 23351 12835
rect 23293 12795 23351 12801
rect 21910 12724 21916 12776
rect 21968 12764 21974 12776
rect 22097 12767 22155 12773
rect 22097 12764 22109 12767
rect 21968 12736 22109 12764
rect 21968 12724 21974 12736
rect 22097 12733 22109 12736
rect 22143 12733 22155 12767
rect 23308 12764 23336 12795
rect 23382 12792 23388 12844
rect 23440 12832 23446 12844
rect 24228 12841 24256 12872
rect 24397 12869 24409 12872
rect 24443 12869 24455 12903
rect 24397 12863 24455 12869
rect 24213 12835 24271 12841
rect 24213 12832 24225 12835
rect 23440 12804 24225 12832
rect 23440 12792 23446 12804
rect 24213 12801 24225 12804
rect 24259 12801 24271 12835
rect 24213 12795 24271 12801
rect 24302 12792 24308 12844
rect 24360 12792 24366 12844
rect 24486 12792 24492 12844
rect 24544 12792 24550 12844
rect 24320 12764 24348 12792
rect 23308 12736 24348 12764
rect 22097 12727 22155 12733
rect 19291 12668 21404 12696
rect 22189 12699 22247 12705
rect 19291 12665 19303 12668
rect 19245 12659 19303 12665
rect 22189 12665 22201 12699
rect 22235 12696 22247 12699
rect 22370 12696 22376 12708
rect 22235 12668 22376 12696
rect 22235 12665 22247 12668
rect 22189 12659 22247 12665
rect 22370 12656 22376 12668
rect 22428 12696 22434 12708
rect 22925 12699 22983 12705
rect 22925 12696 22937 12699
rect 22428 12668 22937 12696
rect 22428 12656 22434 12668
rect 22925 12665 22937 12668
rect 22971 12665 22983 12699
rect 22925 12659 22983 12665
rect 23937 12699 23995 12705
rect 23937 12665 23949 12699
rect 23983 12696 23995 12699
rect 24504 12696 24532 12792
rect 23983 12668 24532 12696
rect 23983 12665 23995 12668
rect 23937 12659 23995 12665
rect 4062 12588 4068 12640
rect 4120 12628 4126 12640
rect 4157 12631 4215 12637
rect 4157 12628 4169 12631
rect 4120 12600 4169 12628
rect 4120 12588 4126 12600
rect 4157 12597 4169 12600
rect 4203 12597 4215 12631
rect 4157 12591 4215 12597
rect 4798 12588 4804 12640
rect 4856 12588 4862 12640
rect 9122 12588 9128 12640
rect 9180 12588 9186 12640
rect 12158 12588 12164 12640
rect 12216 12588 12222 12640
rect 17402 12588 17408 12640
rect 17460 12628 17466 12640
rect 17497 12631 17555 12637
rect 17497 12628 17509 12631
rect 17460 12600 17509 12628
rect 17460 12588 17466 12600
rect 17497 12597 17509 12600
rect 17543 12597 17555 12631
rect 17497 12591 17555 12597
rect 17957 12631 18015 12637
rect 17957 12597 17969 12631
rect 18003 12628 18015 12631
rect 18414 12628 18420 12640
rect 18003 12600 18420 12628
rect 18003 12597 18015 12600
rect 17957 12591 18015 12597
rect 18414 12588 18420 12600
rect 18472 12588 18478 12640
rect 19889 12631 19947 12637
rect 19889 12597 19901 12631
rect 19935 12628 19947 12631
rect 19978 12628 19984 12640
rect 19935 12600 19984 12628
rect 19935 12597 19947 12600
rect 19889 12591 19947 12597
rect 19978 12588 19984 12600
rect 20036 12588 20042 12640
rect 20990 12588 20996 12640
rect 21048 12588 21054 12640
rect 21174 12588 21180 12640
rect 21232 12628 21238 12640
rect 22281 12631 22339 12637
rect 22281 12628 22293 12631
rect 21232 12600 22293 12628
rect 21232 12588 21238 12600
rect 22281 12597 22293 12600
rect 22327 12597 22339 12631
rect 22281 12591 22339 12597
rect 22462 12588 22468 12640
rect 22520 12628 22526 12640
rect 22830 12628 22836 12640
rect 22520 12600 22836 12628
rect 22520 12588 22526 12600
rect 22830 12588 22836 12600
rect 22888 12588 22894 12640
rect 23382 12588 23388 12640
rect 23440 12588 23446 12640
rect 23566 12588 23572 12640
rect 23624 12588 23630 12640
rect 1104 12538 25208 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 25208 12538
rect 1104 12464 25208 12486
rect 6638 12384 6644 12436
rect 6696 12424 6702 12436
rect 9582 12424 9588 12436
rect 6696 12396 9588 12424
rect 6696 12384 6702 12396
rect 9582 12384 9588 12396
rect 9640 12384 9646 12436
rect 10686 12384 10692 12436
rect 10744 12433 10750 12436
rect 10744 12427 10793 12433
rect 10744 12393 10747 12427
rect 10781 12393 10793 12427
rect 10744 12387 10793 12393
rect 16623 12427 16681 12433
rect 16623 12393 16635 12427
rect 16669 12424 16681 12427
rect 17034 12424 17040 12436
rect 16669 12396 17040 12424
rect 16669 12393 16681 12396
rect 16623 12387 16681 12393
rect 10744 12384 10750 12387
rect 17034 12384 17040 12396
rect 17092 12384 17098 12436
rect 17405 12427 17463 12433
rect 17405 12393 17417 12427
rect 17451 12424 17463 12427
rect 17494 12424 17500 12436
rect 17451 12396 17500 12424
rect 17451 12393 17463 12396
rect 17405 12387 17463 12393
rect 17494 12384 17500 12396
rect 17552 12384 17558 12436
rect 17589 12427 17647 12433
rect 17589 12393 17601 12427
rect 17635 12424 17647 12427
rect 17862 12424 17868 12436
rect 17635 12396 17868 12424
rect 17635 12393 17647 12396
rect 17589 12387 17647 12393
rect 17862 12384 17868 12396
rect 17920 12384 17926 12436
rect 18325 12427 18383 12433
rect 18325 12393 18337 12427
rect 18371 12424 18383 12427
rect 18782 12424 18788 12436
rect 18371 12396 18788 12424
rect 18371 12393 18383 12396
rect 18325 12387 18383 12393
rect 18782 12384 18788 12396
rect 18840 12384 18846 12436
rect 19429 12427 19487 12433
rect 19429 12393 19441 12427
rect 19475 12424 19487 12427
rect 22094 12424 22100 12436
rect 19475 12396 22100 12424
rect 19475 12393 19487 12396
rect 19429 12387 19487 12393
rect 22094 12384 22100 12396
rect 22152 12384 22158 12436
rect 22370 12384 22376 12436
rect 22428 12384 22434 12436
rect 22462 12384 22468 12436
rect 22520 12424 22526 12436
rect 22722 12427 22780 12433
rect 22722 12424 22734 12427
rect 22520 12396 22734 12424
rect 22520 12384 22526 12396
rect 22722 12393 22734 12396
rect 22768 12393 22780 12427
rect 22722 12387 22780 12393
rect 24026 12384 24032 12436
rect 24084 12424 24090 12436
rect 24213 12427 24271 12433
rect 24213 12424 24225 12427
rect 24084 12396 24225 12424
rect 24084 12384 24090 12396
rect 24213 12393 24225 12396
rect 24259 12393 24271 12427
rect 24213 12387 24271 12393
rect 11701 12359 11759 12365
rect 11701 12325 11713 12359
rect 11747 12356 11759 12359
rect 12342 12356 12348 12368
rect 11747 12328 12348 12356
rect 11747 12325 11759 12328
rect 11701 12319 11759 12325
rect 12342 12316 12348 12328
rect 12400 12356 12406 12368
rect 13081 12359 13139 12365
rect 13081 12356 13093 12359
rect 12400 12328 13093 12356
rect 12400 12316 12406 12328
rect 13081 12325 13093 12328
rect 13127 12325 13139 12359
rect 17052 12356 17080 12384
rect 17773 12359 17831 12365
rect 17773 12356 17785 12359
rect 17052 12328 17785 12356
rect 13081 12319 13139 12325
rect 17773 12325 17785 12328
rect 17819 12325 17831 12359
rect 17773 12319 17831 12325
rect 18141 12359 18199 12365
rect 18141 12325 18153 12359
rect 18187 12356 18199 12359
rect 19702 12356 19708 12368
rect 18187 12328 19708 12356
rect 18187 12325 18199 12328
rect 18141 12319 18199 12325
rect 19702 12316 19708 12328
rect 19760 12316 19766 12368
rect 21450 12356 21456 12368
rect 20180 12328 21456 12356
rect 1397 12291 1455 12297
rect 1397 12257 1409 12291
rect 1443 12288 1455 12291
rect 3789 12291 3847 12297
rect 3789 12288 3801 12291
rect 1443 12260 3801 12288
rect 1443 12257 1455 12260
rect 1397 12251 1455 12257
rect 3789 12257 3801 12260
rect 3835 12288 3847 12291
rect 4614 12288 4620 12300
rect 3835 12260 4620 12288
rect 3835 12257 3847 12260
rect 3789 12251 3847 12257
rect 4614 12248 4620 12260
rect 4672 12248 4678 12300
rect 9122 12248 9128 12300
rect 9180 12288 9186 12300
rect 9309 12291 9367 12297
rect 9309 12288 9321 12291
rect 9180 12260 9321 12288
rect 9180 12248 9186 12260
rect 9309 12257 9321 12260
rect 9355 12257 9367 12291
rect 9309 12251 9367 12257
rect 11149 12291 11207 12297
rect 11149 12257 11161 12291
rect 11195 12288 11207 12291
rect 11606 12288 11612 12300
rect 11195 12260 11612 12288
rect 11195 12257 11207 12260
rect 11149 12251 11207 12257
rect 3418 12180 3424 12232
rect 3476 12180 3482 12232
rect 4154 12180 4160 12232
rect 4212 12180 4218 12232
rect 6822 12180 6828 12232
rect 6880 12220 6886 12232
rect 8941 12223 8999 12229
rect 8941 12220 8953 12223
rect 6880 12192 8953 12220
rect 6880 12180 6886 12192
rect 8941 12189 8953 12192
rect 8987 12220 8999 12223
rect 9214 12220 9220 12232
rect 8987 12192 9220 12220
rect 8987 12189 8999 12192
rect 8941 12183 8999 12189
rect 9214 12180 9220 12192
rect 9272 12180 9278 12232
rect 1670 12112 1676 12164
rect 1728 12112 1734 12164
rect 5718 12152 5724 12164
rect 2898 12124 3924 12152
rect 5198 12124 5724 12152
rect 3142 12044 3148 12096
rect 3200 12044 3206 12096
rect 3326 12044 3332 12096
rect 3384 12044 3390 12096
rect 3896 12084 3924 12124
rect 5276 12084 5304 12124
rect 5718 12112 5724 12124
rect 5776 12152 5782 12164
rect 7098 12152 7104 12164
rect 5776 12124 7104 12152
rect 5776 12112 5782 12124
rect 7098 12112 7104 12124
rect 7156 12112 7162 12164
rect 9674 12112 9680 12164
rect 9732 12112 9738 12164
rect 3896 12056 5304 12084
rect 5583 12087 5641 12093
rect 5583 12053 5595 12087
rect 5629 12084 5641 12087
rect 6270 12084 6276 12096
rect 5629 12056 6276 12084
rect 5629 12053 5641 12056
rect 5583 12047 5641 12053
rect 6270 12044 6276 12056
rect 6328 12044 6334 12096
rect 8662 12044 8668 12096
rect 8720 12084 8726 12096
rect 11164 12084 11192 12251
rect 11606 12248 11612 12260
rect 11664 12248 11670 12300
rect 12250 12248 12256 12300
rect 12308 12248 12314 12300
rect 15197 12291 15255 12297
rect 15197 12257 15209 12291
rect 15243 12288 15255 12291
rect 16942 12288 16948 12300
rect 15243 12260 16948 12288
rect 15243 12257 15255 12260
rect 15197 12251 15255 12257
rect 16942 12248 16948 12260
rect 17000 12248 17006 12300
rect 17494 12248 17500 12300
rect 17552 12288 17558 12300
rect 19797 12291 19855 12297
rect 19797 12288 19809 12291
rect 17552 12260 18368 12288
rect 17552 12248 17558 12260
rect 11330 12180 11336 12232
rect 11388 12180 11394 12232
rect 11422 12180 11428 12232
rect 11480 12180 11486 12232
rect 11514 12180 11520 12232
rect 11572 12180 11578 12232
rect 12158 12220 12164 12232
rect 12119 12192 12164 12220
rect 12158 12180 12164 12192
rect 12216 12220 12222 12232
rect 12621 12223 12679 12229
rect 12621 12220 12633 12223
rect 12216 12192 12633 12220
rect 12216 12180 12222 12192
rect 12621 12189 12633 12192
rect 12667 12189 12679 12223
rect 12621 12183 12679 12189
rect 12802 12180 12808 12232
rect 12860 12180 12866 12232
rect 13354 12180 13360 12232
rect 13412 12180 13418 12232
rect 14826 12180 14832 12232
rect 14884 12180 14890 12232
rect 17586 12220 17592 12232
rect 17236 12192 17592 12220
rect 11348 12152 11376 12180
rect 12066 12152 12072 12164
rect 11348 12124 12072 12152
rect 12066 12112 12072 12124
rect 12124 12112 12130 12164
rect 13170 12152 13176 12164
rect 12544 12124 13176 12152
rect 12544 12093 12572 12124
rect 13170 12112 13176 12124
rect 13228 12152 13234 12164
rect 13541 12155 13599 12161
rect 13541 12152 13553 12155
rect 13228 12124 13553 12152
rect 13228 12112 13234 12124
rect 13541 12121 13553 12124
rect 13587 12121 13599 12155
rect 16390 12152 16396 12164
rect 16238 12124 16396 12152
rect 13541 12115 13599 12121
rect 16390 12112 16396 12124
rect 16448 12112 16454 12164
rect 17236 12161 17264 12192
rect 17586 12180 17592 12192
rect 17644 12180 17650 12232
rect 17681 12223 17739 12229
rect 17681 12189 17693 12223
rect 17727 12189 17739 12223
rect 17681 12183 17739 12189
rect 17957 12223 18015 12229
rect 17957 12189 17969 12223
rect 18003 12189 18015 12223
rect 17957 12183 18015 12189
rect 17221 12155 17279 12161
rect 17221 12121 17233 12155
rect 17267 12121 17279 12155
rect 17221 12115 17279 12121
rect 17402 12112 17408 12164
rect 17460 12161 17466 12164
rect 17460 12155 17479 12161
rect 17467 12121 17479 12155
rect 17460 12115 17479 12121
rect 17460 12112 17466 12115
rect 17696 12096 17724 12183
rect 8720 12056 11192 12084
rect 12529 12087 12587 12093
rect 8720 12044 8726 12056
rect 12529 12053 12541 12087
rect 12575 12053 12587 12087
rect 12529 12047 12587 12053
rect 12710 12044 12716 12096
rect 12768 12084 12774 12096
rect 12897 12087 12955 12093
rect 12897 12084 12909 12087
rect 12768 12056 12909 12084
rect 12768 12044 12774 12056
rect 12897 12053 12909 12056
rect 12943 12053 12955 12087
rect 12897 12047 12955 12053
rect 13725 12087 13783 12093
rect 13725 12053 13737 12087
rect 13771 12084 13783 12087
rect 13906 12084 13912 12096
rect 13771 12056 13912 12084
rect 13771 12053 13783 12056
rect 13725 12047 13783 12053
rect 13906 12044 13912 12056
rect 13964 12044 13970 12096
rect 17126 12044 17132 12096
rect 17184 12084 17190 12096
rect 17678 12084 17684 12096
rect 17184 12056 17684 12084
rect 17184 12044 17190 12056
rect 17678 12044 17684 12056
rect 17736 12044 17742 12096
rect 17972 12084 18000 12183
rect 18230 12180 18236 12232
rect 18288 12180 18294 12232
rect 18340 12220 18368 12260
rect 18524 12260 19809 12288
rect 18524 12232 18552 12260
rect 19797 12257 19809 12260
rect 19843 12257 19855 12291
rect 19797 12251 19855 12257
rect 18414 12220 18420 12232
rect 18340 12192 18420 12220
rect 18414 12180 18420 12192
rect 18472 12180 18478 12232
rect 18506 12180 18512 12232
rect 18564 12180 18570 12232
rect 18693 12223 18751 12229
rect 18693 12189 18705 12223
rect 18739 12220 18751 12223
rect 18782 12220 18788 12232
rect 18739 12192 18788 12220
rect 18739 12189 18751 12192
rect 18693 12183 18751 12189
rect 18782 12180 18788 12192
rect 18840 12180 18846 12232
rect 18877 12223 18935 12229
rect 18877 12189 18889 12223
rect 18923 12220 18935 12223
rect 19058 12220 19064 12232
rect 18923 12192 19064 12220
rect 18923 12189 18935 12192
rect 18877 12183 18935 12189
rect 19058 12180 19064 12192
rect 19116 12180 19122 12232
rect 19610 12180 19616 12232
rect 19668 12180 19674 12232
rect 19886 12180 19892 12232
rect 19944 12180 19950 12232
rect 20180 12229 20208 12328
rect 21450 12316 21456 12328
rect 21508 12356 21514 12368
rect 21545 12359 21603 12365
rect 21545 12356 21557 12359
rect 21508 12328 21557 12356
rect 21508 12316 21514 12328
rect 21545 12325 21557 12328
rect 21591 12325 21603 12359
rect 22186 12356 22192 12368
rect 21545 12319 21603 12325
rect 21744 12328 22192 12356
rect 20714 12248 20720 12300
rect 20772 12288 20778 12300
rect 20993 12291 21051 12297
rect 20993 12288 21005 12291
rect 20772 12260 21005 12288
rect 20772 12248 20778 12260
rect 20993 12257 21005 12260
rect 21039 12257 21051 12291
rect 20993 12251 21051 12257
rect 21082 12248 21088 12300
rect 21140 12288 21146 12300
rect 21634 12288 21640 12300
rect 21140 12260 21640 12288
rect 21140 12248 21146 12260
rect 19981 12223 20039 12229
rect 19981 12189 19993 12223
rect 20027 12189 20039 12223
rect 19981 12183 20039 12189
rect 20165 12223 20223 12229
rect 20165 12189 20177 12223
rect 20211 12189 20223 12223
rect 20165 12183 20223 12189
rect 18601 12155 18659 12161
rect 18601 12121 18613 12155
rect 18647 12152 18659 12155
rect 19996 12152 20024 12183
rect 20622 12180 20628 12232
rect 20680 12180 20686 12232
rect 20898 12180 20904 12232
rect 20956 12180 20962 12232
rect 21376 12229 21404 12260
rect 21634 12248 21640 12260
rect 21692 12248 21698 12300
rect 21177 12223 21235 12229
rect 21177 12189 21189 12223
rect 21223 12220 21235 12223
rect 21361 12223 21419 12229
rect 21223 12192 21312 12220
rect 21223 12189 21235 12192
rect 21177 12183 21235 12189
rect 20070 12152 20076 12164
rect 18647 12124 20076 12152
rect 18647 12121 18659 12124
rect 18601 12115 18659 12121
rect 20070 12112 20076 12124
rect 20128 12112 20134 12164
rect 21284 12152 21312 12192
rect 21361 12189 21373 12223
rect 21407 12189 21419 12223
rect 21361 12183 21419 12189
rect 21450 12180 21456 12232
rect 21508 12180 21514 12232
rect 21744 12229 21772 12328
rect 22186 12316 22192 12328
rect 22244 12316 22250 12368
rect 22002 12248 22008 12300
rect 22060 12248 22066 12300
rect 22097 12291 22155 12297
rect 22097 12257 22109 12291
rect 22143 12288 22155 12291
rect 22370 12288 22376 12300
rect 22143 12260 22376 12288
rect 22143 12257 22155 12260
rect 22097 12251 22155 12257
rect 22370 12248 22376 12260
rect 22428 12248 22434 12300
rect 22462 12248 22468 12300
rect 22520 12288 22526 12300
rect 24854 12288 24860 12300
rect 22520 12260 24860 12288
rect 22520 12248 22526 12260
rect 24854 12248 24860 12260
rect 24912 12248 24918 12300
rect 21729 12223 21787 12229
rect 21729 12189 21741 12223
rect 21775 12189 21787 12223
rect 21729 12183 21787 12189
rect 21910 12180 21916 12232
rect 21968 12180 21974 12232
rect 22189 12223 22247 12229
rect 22189 12189 22201 12223
rect 22235 12189 22247 12223
rect 22189 12183 22247 12189
rect 22204 12152 22232 12183
rect 22830 12152 22836 12164
rect 20364 12124 21220 12152
rect 21284 12124 22140 12152
rect 22204 12124 22836 12152
rect 20364 12084 20392 12124
rect 17972 12056 20392 12084
rect 20438 12044 20444 12096
rect 20496 12044 20502 12096
rect 20809 12087 20867 12093
rect 20809 12053 20821 12087
rect 20855 12084 20867 12087
rect 21082 12084 21088 12096
rect 20855 12056 21088 12084
rect 20855 12053 20867 12056
rect 20809 12047 20867 12053
rect 21082 12044 21088 12056
rect 21140 12044 21146 12096
rect 21192 12084 21220 12124
rect 21266 12084 21272 12096
rect 21192 12056 21272 12084
rect 21266 12044 21272 12056
rect 21324 12084 21330 12096
rect 21910 12084 21916 12096
rect 21324 12056 21916 12084
rect 21324 12044 21330 12056
rect 21910 12044 21916 12056
rect 21968 12044 21974 12096
rect 22112 12084 22140 12124
rect 22830 12112 22836 12124
rect 22888 12112 22894 12164
rect 23198 12112 23204 12164
rect 23256 12112 23262 12164
rect 22278 12084 22284 12096
rect 22112 12056 22284 12084
rect 22278 12044 22284 12056
rect 22336 12044 22342 12096
rect 1104 11994 25208 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 25208 11994
rect 1104 11920 25208 11942
rect 1670 11840 1676 11892
rect 1728 11880 1734 11892
rect 2133 11883 2191 11889
rect 2133 11880 2145 11883
rect 1728 11852 2145 11880
rect 1728 11840 1734 11852
rect 2133 11849 2145 11852
rect 2179 11849 2191 11883
rect 2133 11843 2191 11849
rect 6546 11840 6552 11892
rect 6604 11880 6610 11892
rect 6825 11883 6883 11889
rect 6825 11880 6837 11883
rect 6604 11852 6837 11880
rect 6604 11840 6610 11852
rect 6825 11849 6837 11852
rect 6871 11849 6883 11883
rect 6825 11843 6883 11849
rect 8294 11840 8300 11892
rect 8352 11880 8358 11892
rect 9674 11880 9680 11892
rect 8352 11852 9680 11880
rect 8352 11840 8358 11852
rect 9674 11840 9680 11852
rect 9732 11880 9738 11892
rect 10134 11880 10140 11892
rect 9732 11852 10140 11880
rect 9732 11840 9738 11852
rect 1949 11815 2007 11821
rect 1949 11781 1961 11815
rect 1995 11812 2007 11815
rect 2501 11815 2559 11821
rect 2501 11812 2513 11815
rect 1995 11784 2513 11812
rect 1995 11781 2007 11784
rect 1949 11775 2007 11781
rect 2501 11781 2513 11784
rect 2547 11812 2559 11815
rect 2869 11815 2927 11821
rect 2869 11812 2881 11815
rect 2547 11784 2881 11812
rect 2547 11781 2559 11784
rect 2501 11775 2559 11781
rect 2869 11781 2881 11784
rect 2915 11781 2927 11815
rect 2869 11775 2927 11781
rect 5718 11772 5724 11824
rect 5776 11772 5782 11824
rect 6135 11815 6193 11821
rect 6135 11781 6147 11815
rect 6181 11812 6193 11815
rect 6638 11812 6644 11824
rect 6181 11784 6644 11812
rect 6181 11781 6193 11784
rect 6135 11775 6193 11781
rect 6638 11772 6644 11784
rect 6696 11772 6702 11824
rect 9876 11812 9904 11852
rect 10134 11840 10140 11852
rect 10192 11840 10198 11892
rect 11514 11840 11520 11892
rect 11572 11880 11578 11892
rect 11572 11852 11836 11880
rect 11572 11840 11578 11852
rect 11011 11815 11069 11821
rect 9876 11784 9982 11812
rect 11011 11781 11023 11815
rect 11057 11812 11069 11815
rect 11422 11812 11428 11824
rect 11057 11784 11428 11812
rect 11057 11781 11069 11784
rect 11011 11775 11069 11781
rect 11422 11772 11428 11784
rect 11480 11812 11486 11824
rect 11808 11821 11836 11852
rect 12250 11840 12256 11892
rect 12308 11840 12314 11892
rect 18046 11840 18052 11892
rect 18104 11880 18110 11892
rect 18233 11883 18291 11889
rect 18233 11880 18245 11883
rect 18104 11852 18245 11880
rect 18104 11840 18110 11852
rect 18233 11849 18245 11852
rect 18279 11849 18291 11883
rect 18233 11843 18291 11849
rect 18506 11840 18512 11892
rect 18564 11880 18570 11892
rect 18601 11883 18659 11889
rect 18601 11880 18613 11883
rect 18564 11852 18613 11880
rect 18564 11840 18570 11852
rect 18601 11849 18613 11852
rect 18647 11849 18659 11883
rect 18601 11843 18659 11849
rect 18782 11840 18788 11892
rect 18840 11880 18846 11892
rect 18840 11852 19012 11880
rect 18840 11840 18846 11852
rect 11793 11815 11851 11821
rect 11480 11784 11744 11812
rect 11480 11772 11486 11784
rect 1670 11704 1676 11756
rect 1728 11704 1734 11756
rect 1765 11747 1823 11753
rect 1765 11713 1777 11747
rect 1811 11713 1823 11747
rect 1765 11707 1823 11713
rect 2041 11747 2099 11753
rect 2041 11713 2053 11747
rect 2087 11744 2099 11747
rect 2314 11744 2320 11756
rect 2087 11716 2320 11744
rect 2087 11713 2099 11716
rect 2041 11707 2099 11713
rect 1780 11608 1808 11707
rect 2314 11704 2320 11716
rect 2372 11704 2378 11756
rect 2593 11747 2651 11753
rect 2593 11713 2605 11747
rect 2639 11744 2651 11747
rect 3326 11744 3332 11756
rect 2639 11716 3332 11744
rect 2639 11713 2651 11716
rect 2593 11707 2651 11713
rect 3326 11704 3332 11716
rect 3384 11704 3390 11756
rect 4709 11747 4767 11753
rect 4709 11713 4721 11747
rect 4755 11744 4767 11747
rect 4798 11744 4804 11756
rect 4755 11716 4804 11744
rect 4755 11713 4767 11716
rect 4709 11707 4767 11713
rect 4798 11704 4804 11716
rect 4856 11704 4862 11756
rect 6730 11704 6736 11756
rect 6788 11704 6794 11756
rect 8113 11747 8171 11753
rect 8113 11713 8125 11747
rect 8159 11744 8171 11747
rect 8662 11744 8668 11756
rect 8159 11716 8668 11744
rect 8159 11713 8171 11716
rect 8113 11707 8171 11713
rect 8662 11704 8668 11716
rect 8720 11704 8726 11756
rect 9214 11704 9220 11756
rect 9272 11704 9278 11756
rect 11606 11704 11612 11756
rect 11664 11704 11670 11756
rect 11716 11744 11744 11784
rect 11793 11781 11805 11815
rect 11839 11781 11851 11815
rect 11793 11775 11851 11781
rect 11885 11815 11943 11821
rect 11885 11781 11897 11815
rect 11931 11812 11943 11815
rect 12066 11812 12072 11824
rect 11931 11784 12072 11812
rect 11931 11781 11943 11784
rect 11885 11775 11943 11781
rect 12066 11772 12072 11784
rect 12124 11772 12130 11824
rect 12802 11812 12808 11824
rect 12176 11784 12808 11812
rect 12176 11753 12204 11784
rect 12802 11772 12808 11784
rect 12860 11772 12866 11824
rect 17954 11772 17960 11824
rect 18012 11812 18018 11824
rect 18693 11815 18751 11821
rect 18693 11812 18705 11815
rect 18012 11784 18705 11812
rect 18012 11772 18018 11784
rect 11982 11747 12040 11753
rect 11716 11742 11836 11744
rect 11982 11742 11994 11747
rect 11716 11716 11994 11742
rect 11808 11714 11994 11716
rect 11982 11713 11994 11714
rect 12028 11713 12040 11747
rect 11982 11707 12040 11713
rect 12161 11747 12219 11753
rect 12161 11713 12173 11747
rect 12207 11713 12219 11747
rect 12161 11707 12219 11713
rect 3142 11636 3148 11688
rect 3200 11676 3206 11688
rect 3421 11679 3479 11685
rect 3421 11676 3433 11679
rect 3200 11648 3433 11676
rect 3200 11636 3206 11648
rect 3421 11645 3433 11648
rect 3467 11645 3479 11679
rect 3421 11639 3479 11645
rect 4062 11636 4068 11688
rect 4120 11676 4126 11688
rect 4157 11679 4215 11685
rect 4157 11676 4169 11679
rect 4120 11648 4169 11676
rect 4120 11636 4126 11648
rect 4157 11645 4169 11648
rect 4203 11645 4215 11679
rect 4157 11639 4215 11645
rect 4341 11679 4399 11685
rect 4341 11645 4353 11679
rect 4387 11676 4399 11679
rect 4614 11676 4620 11688
rect 4387 11648 4620 11676
rect 4387 11645 4399 11648
rect 4341 11639 4399 11645
rect 4614 11636 4620 11648
rect 4672 11636 4678 11688
rect 6914 11636 6920 11688
rect 6972 11636 6978 11688
rect 7834 11636 7840 11688
rect 7892 11676 7898 11688
rect 8205 11679 8263 11685
rect 8205 11676 8217 11679
rect 7892 11648 8217 11676
rect 7892 11636 7898 11648
rect 8205 11645 8217 11648
rect 8251 11645 8263 11679
rect 8205 11639 8263 11645
rect 8297 11679 8355 11685
rect 8297 11645 8309 11679
rect 8343 11645 8355 11679
rect 8297 11639 8355 11645
rect 9585 11679 9643 11685
rect 9585 11645 9597 11679
rect 9631 11676 9643 11679
rect 9766 11676 9772 11688
rect 9631 11648 9772 11676
rect 9631 11645 9643 11648
rect 9585 11639 9643 11645
rect 3605 11611 3663 11617
rect 3605 11608 3617 11611
rect 1780 11580 3617 11608
rect 3605 11577 3617 11580
rect 3651 11577 3663 11611
rect 8312 11608 8340 11639
rect 9766 11636 9772 11648
rect 9824 11636 9830 11688
rect 11793 11679 11851 11685
rect 11793 11645 11805 11679
rect 11839 11676 11851 11679
rect 12176 11676 12204 11707
rect 12342 11704 12348 11756
rect 12400 11704 12406 11756
rect 12621 11747 12679 11753
rect 12621 11713 12633 11747
rect 12667 11744 12679 11747
rect 12667 11716 13124 11744
rect 12667 11713 12679 11716
rect 12621 11707 12679 11713
rect 11839 11648 12204 11676
rect 11839 11645 11851 11648
rect 11793 11639 11851 11645
rect 12710 11636 12716 11688
rect 12768 11636 12774 11688
rect 13096 11676 13124 11716
rect 13170 11704 13176 11756
rect 13228 11704 13234 11756
rect 13354 11704 13360 11756
rect 13412 11704 13418 11756
rect 13906 11704 13912 11756
rect 13964 11704 13970 11756
rect 18138 11704 18144 11756
rect 18196 11704 18202 11756
rect 18432 11753 18460 11784
rect 18693 11781 18705 11784
rect 18739 11781 18751 11815
rect 18893 11815 18951 11821
rect 18893 11812 18905 11815
rect 18693 11775 18751 11781
rect 18800 11784 18905 11812
rect 18417 11747 18475 11753
rect 18417 11713 18429 11747
rect 18463 11713 18475 11747
rect 18417 11707 18475 11713
rect 13265 11679 13323 11685
rect 13265 11676 13277 11679
rect 13096 11648 13277 11676
rect 13265 11645 13277 11648
rect 13311 11676 13323 11679
rect 13725 11679 13783 11685
rect 13725 11676 13737 11679
rect 13311 11648 13737 11676
rect 13311 11645 13323 11648
rect 13265 11639 13323 11645
rect 13725 11645 13737 11648
rect 13771 11645 13783 11679
rect 18156 11676 18184 11704
rect 18800 11676 18828 11784
rect 18893 11781 18905 11784
rect 18939 11781 18951 11815
rect 18893 11775 18951 11781
rect 18156 11648 18828 11676
rect 18984 11676 19012 11852
rect 19058 11840 19064 11892
rect 19116 11840 19122 11892
rect 19521 11883 19579 11889
rect 19521 11849 19533 11883
rect 19567 11880 19579 11883
rect 19886 11880 19892 11892
rect 19567 11852 19892 11880
rect 19567 11849 19579 11852
rect 19521 11843 19579 11849
rect 19886 11840 19892 11852
rect 19944 11840 19950 11892
rect 20990 11880 20996 11892
rect 20088 11852 20996 11880
rect 19076 11744 19104 11840
rect 19337 11747 19395 11753
rect 19337 11744 19349 11747
rect 19076 11716 19349 11744
rect 19337 11713 19349 11716
rect 19383 11713 19395 11747
rect 19337 11707 19395 11713
rect 19978 11704 19984 11756
rect 20036 11704 20042 11756
rect 20088 11753 20116 11852
rect 20990 11840 20996 11852
rect 21048 11840 21054 11892
rect 22373 11883 22431 11889
rect 22373 11849 22385 11883
rect 22419 11880 22431 11883
rect 24578 11880 24584 11892
rect 22419 11852 24584 11880
rect 22419 11849 22431 11852
rect 22373 11843 22431 11849
rect 24578 11840 24584 11852
rect 24636 11840 24642 11892
rect 20073 11747 20131 11753
rect 20073 11713 20085 11747
rect 20119 11713 20131 11747
rect 20073 11707 20131 11713
rect 20254 11704 20260 11756
rect 20312 11704 20318 11756
rect 20349 11747 20407 11753
rect 20349 11713 20361 11747
rect 20395 11713 20407 11747
rect 20349 11707 20407 11713
rect 19153 11679 19211 11685
rect 19153 11676 19165 11679
rect 18984 11648 19165 11676
rect 13725 11639 13783 11645
rect 19153 11645 19165 11648
rect 19199 11676 19211 11679
rect 19610 11676 19616 11688
rect 19199 11648 19616 11676
rect 19199 11645 19211 11648
rect 19153 11639 19211 11645
rect 19610 11636 19616 11648
rect 19668 11636 19674 11688
rect 20162 11636 20168 11688
rect 20220 11676 20226 11688
rect 20364 11676 20392 11707
rect 21910 11704 21916 11756
rect 21968 11704 21974 11756
rect 22005 11747 22063 11753
rect 22005 11713 22017 11747
rect 22051 11713 22063 11747
rect 22005 11707 22063 11713
rect 20220 11648 20392 11676
rect 20220 11636 20226 11648
rect 21358 11636 21364 11688
rect 21416 11676 21422 11688
rect 22020 11676 22048 11707
rect 22186 11704 22192 11756
rect 22244 11704 22250 11756
rect 22370 11676 22376 11688
rect 21416 11648 22376 11676
rect 21416 11636 21422 11648
rect 22370 11636 22376 11648
rect 22428 11676 22434 11688
rect 23106 11676 23112 11688
rect 22428 11648 23112 11676
rect 22428 11636 22434 11648
rect 23106 11636 23112 11648
rect 23164 11636 23170 11688
rect 3605 11571 3663 11577
rect 6288 11580 8340 11608
rect 842 11500 848 11552
rect 900 11540 906 11552
rect 1489 11543 1547 11549
rect 1489 11540 1501 11543
rect 900 11512 1501 11540
rect 900 11500 906 11512
rect 1489 11509 1501 11512
rect 1535 11509 1547 11543
rect 1489 11503 1547 11509
rect 1578 11500 1584 11552
rect 1636 11540 1642 11552
rect 1765 11543 1823 11549
rect 1765 11540 1777 11543
rect 1636 11512 1777 11540
rect 1636 11500 1642 11512
rect 1765 11509 1777 11512
rect 1811 11509 1823 11543
rect 1765 11503 1823 11509
rect 4706 11500 4712 11552
rect 4764 11540 4770 11552
rect 6288 11540 6316 11580
rect 4764 11512 6316 11540
rect 4764 11500 4770 11512
rect 6362 11500 6368 11552
rect 6420 11500 6426 11552
rect 7282 11500 7288 11552
rect 7340 11540 7346 11552
rect 7745 11543 7803 11549
rect 7745 11540 7757 11543
rect 7340 11512 7757 11540
rect 7340 11500 7346 11512
rect 7745 11509 7757 11512
rect 7791 11509 7803 11543
rect 8312 11540 8340 11580
rect 12989 11611 13047 11617
rect 12989 11577 13001 11611
rect 13035 11608 13047 11611
rect 13446 11608 13452 11620
rect 13035 11580 13452 11608
rect 13035 11577 13047 11580
rect 12989 11571 13047 11577
rect 13446 11568 13452 11580
rect 13504 11568 13510 11620
rect 21818 11568 21824 11620
rect 21876 11608 21882 11620
rect 22462 11608 22468 11620
rect 21876 11580 22468 11608
rect 21876 11568 21882 11580
rect 22462 11568 22468 11580
rect 22520 11568 22526 11620
rect 9858 11540 9864 11552
rect 8312 11512 9864 11540
rect 7745 11503 7803 11509
rect 9858 11500 9864 11512
rect 9916 11540 9922 11552
rect 10318 11540 10324 11552
rect 9916 11512 10324 11540
rect 9916 11500 9922 11512
rect 10318 11500 10324 11512
rect 10376 11500 10382 11552
rect 14093 11543 14151 11549
rect 14093 11509 14105 11543
rect 14139 11540 14151 11543
rect 17954 11540 17960 11552
rect 14139 11512 17960 11540
rect 14139 11509 14151 11512
rect 14093 11503 14151 11509
rect 17954 11500 17960 11512
rect 18012 11500 18018 11552
rect 18046 11500 18052 11552
rect 18104 11540 18110 11552
rect 18877 11543 18935 11549
rect 18877 11540 18889 11543
rect 18104 11512 18889 11540
rect 18104 11500 18110 11512
rect 18877 11509 18889 11512
rect 18923 11509 18935 11543
rect 18877 11503 18935 11509
rect 20533 11543 20591 11549
rect 20533 11509 20545 11543
rect 20579 11540 20591 11543
rect 21358 11540 21364 11552
rect 20579 11512 21364 11540
rect 20579 11509 20591 11512
rect 20533 11503 20591 11509
rect 21358 11500 21364 11512
rect 21416 11500 21422 11552
rect 1104 11450 25208 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 25208 11450
rect 1104 11376 25208 11398
rect 1670 11336 1676 11348
rect 1412 11308 1676 11336
rect 1412 11141 1440 11308
rect 1670 11296 1676 11308
rect 1728 11336 1734 11348
rect 3418 11336 3424 11348
rect 1728 11308 3424 11336
rect 1728 11296 1734 11308
rect 3418 11296 3424 11308
rect 3476 11336 3482 11348
rect 4249 11339 4307 11345
rect 4249 11336 4261 11339
rect 3476 11308 4261 11336
rect 3476 11296 3482 11308
rect 4249 11305 4261 11308
rect 4295 11305 4307 11339
rect 4249 11299 4307 11305
rect 6730 11296 6736 11348
rect 6788 11345 6794 11348
rect 6788 11339 6837 11345
rect 6788 11305 6791 11339
rect 6825 11336 6837 11339
rect 8478 11336 8484 11348
rect 6825 11308 8484 11336
rect 6825 11305 6837 11308
rect 6788 11299 6837 11305
rect 6788 11296 6794 11299
rect 8478 11296 8484 11308
rect 8536 11296 8542 11348
rect 8662 11296 8668 11348
rect 8720 11296 8726 11348
rect 9766 11296 9772 11348
rect 9824 11296 9830 11348
rect 15562 11296 15568 11348
rect 15620 11336 15626 11348
rect 17126 11336 17132 11348
rect 15620 11308 17132 11336
rect 15620 11296 15626 11308
rect 17126 11296 17132 11308
rect 17184 11296 17190 11348
rect 19981 11339 20039 11345
rect 19981 11305 19993 11339
rect 20027 11336 20039 11339
rect 20162 11336 20168 11348
rect 20027 11308 20168 11336
rect 20027 11305 20039 11308
rect 19981 11299 20039 11305
rect 20162 11296 20168 11308
rect 20220 11296 20226 11348
rect 20254 11296 20260 11348
rect 20312 11336 20318 11348
rect 20717 11339 20775 11345
rect 20717 11336 20729 11339
rect 20312 11308 20729 11336
rect 20312 11296 20318 11308
rect 20717 11305 20729 11308
rect 20763 11305 20775 11339
rect 20717 11299 20775 11305
rect 21910 11296 21916 11348
rect 21968 11296 21974 11348
rect 22094 11296 22100 11348
rect 22152 11336 22158 11348
rect 22152 11308 22508 11336
rect 22152 11296 22158 11308
rect 10134 11228 10140 11280
rect 10192 11268 10198 11280
rect 10597 11271 10655 11277
rect 10597 11268 10609 11271
rect 10192 11240 10609 11268
rect 10192 11228 10198 11240
rect 10597 11237 10609 11240
rect 10643 11237 10655 11271
rect 10597 11231 10655 11237
rect 11606 11228 11612 11280
rect 11664 11268 11670 11280
rect 12713 11271 12771 11277
rect 12713 11268 12725 11271
rect 11664 11240 12725 11268
rect 11664 11228 11670 11240
rect 12713 11237 12725 11240
rect 12759 11268 12771 11271
rect 12759 11240 13676 11268
rect 12759 11237 12771 11240
rect 12713 11231 12771 11237
rect 1673 11203 1731 11209
rect 1673 11169 1685 11203
rect 1719 11200 1731 11203
rect 1719 11172 4108 11200
rect 1719 11169 1731 11172
rect 1673 11163 1731 11169
rect 1397 11135 1455 11141
rect 1397 11101 1409 11135
rect 1443 11101 1455 11135
rect 1397 11095 1455 11101
rect 1578 11092 1584 11144
rect 1636 11092 1642 11144
rect 3234 11132 3240 11144
rect 3082 11104 3240 11132
rect 3234 11092 3240 11104
rect 3292 11092 3298 11144
rect 4080 11141 4108 11172
rect 4614 11160 4620 11212
rect 4672 11160 4678 11212
rect 5353 11203 5411 11209
rect 5353 11169 5365 11203
rect 5399 11200 5411 11203
rect 6362 11200 6368 11212
rect 5399 11172 6368 11200
rect 5399 11169 5411 11172
rect 5353 11163 5411 11169
rect 6362 11160 6368 11172
rect 6420 11160 6426 11212
rect 6822 11160 6828 11212
rect 6880 11200 6886 11212
rect 6917 11203 6975 11209
rect 6917 11200 6929 11203
rect 6880 11172 6929 11200
rect 6880 11160 6886 11172
rect 6917 11169 6929 11172
rect 6963 11169 6975 11203
rect 6917 11163 6975 11169
rect 7282 11160 7288 11212
rect 7340 11160 7346 11212
rect 7392 11172 8432 11200
rect 4065 11135 4123 11141
rect 4065 11101 4077 11135
rect 4111 11132 4123 11135
rect 4154 11132 4160 11144
rect 4111 11104 4160 11132
rect 4111 11101 4123 11104
rect 4065 11095 4123 11101
rect 4154 11092 4160 11104
rect 4212 11132 4218 11144
rect 4632 11132 4660 11160
rect 4985 11135 5043 11141
rect 4985 11132 4997 11135
rect 4212 11104 4997 11132
rect 4212 11092 4218 11104
rect 4985 11101 4997 11104
rect 5031 11101 5043 11135
rect 4985 11095 5043 11101
rect 6270 11092 6276 11144
rect 6328 11132 6334 11144
rect 7392 11132 7420 11172
rect 6328 11104 7420 11132
rect 6328 11092 6334 11104
rect 8300 11076 8352 11082
rect 1489 11067 1547 11073
rect 1489 11033 1501 11067
rect 1535 11064 1547 11067
rect 1949 11067 2007 11073
rect 1949 11064 1961 11067
rect 1535 11036 1961 11064
rect 1535 11033 1547 11036
rect 1489 11027 1547 11033
rect 1949 11033 1961 11036
rect 1995 11033 2007 11067
rect 1949 11027 2007 11033
rect 4433 11067 4491 11073
rect 4433 11033 4445 11067
rect 4479 11064 4491 11067
rect 4522 11064 4528 11076
rect 4479 11036 4528 11064
rect 4479 11033 4491 11036
rect 4433 11027 4491 11033
rect 4522 11024 4528 11036
rect 4580 11024 4586 11076
rect 4617 11067 4675 11073
rect 4617 11033 4629 11067
rect 4663 11033 4675 11067
rect 4617 11027 4675 11033
rect 3234 10956 3240 11008
rect 3292 10996 3298 11008
rect 3421 10999 3479 11005
rect 3421 10996 3433 10999
rect 3292 10968 3433 10996
rect 3292 10956 3298 10968
rect 3421 10965 3433 10968
rect 3467 10996 3479 10999
rect 4062 10996 4068 11008
rect 3467 10968 4068 10996
rect 3467 10965 3479 10968
rect 3421 10959 3479 10965
rect 4062 10956 4068 10968
rect 4120 10956 4126 11008
rect 4246 10956 4252 11008
rect 4304 10996 4310 11008
rect 4632 10996 4660 11027
rect 5718 11024 5724 11076
rect 5776 11024 5782 11076
rect 8404 11064 8432 11172
rect 10318 11160 10324 11212
rect 10376 11160 10382 11212
rect 12066 11160 12072 11212
rect 12124 11200 12130 11212
rect 12124 11172 13584 11200
rect 12124 11160 12130 11172
rect 13004 11141 13032 11172
rect 10137 11135 10195 11141
rect 10137 11101 10149 11135
rect 10183 11132 10195 11135
rect 12989 11135 13047 11141
rect 10183 11104 11468 11132
rect 10183 11101 10195 11104
rect 10137 11095 10195 11101
rect 11440 11076 11468 11104
rect 12989 11101 13001 11135
rect 13035 11101 13047 11135
rect 12989 11095 13047 11101
rect 13265 11135 13323 11141
rect 13265 11101 13277 11135
rect 13311 11132 13323 11135
rect 13354 11132 13360 11144
rect 13311 11104 13360 11132
rect 13311 11101 13323 11104
rect 13265 11095 13323 11101
rect 13354 11092 13360 11104
rect 13412 11092 13418 11144
rect 13556 11141 13584 11172
rect 13648 11144 13676 11240
rect 20346 11228 20352 11280
rect 20404 11268 20410 11280
rect 20809 11271 20867 11277
rect 20809 11268 20821 11271
rect 20404 11240 20821 11268
rect 20404 11228 20410 11240
rect 20809 11237 20821 11240
rect 20855 11237 20867 11271
rect 20809 11231 20867 11237
rect 21821 11271 21879 11277
rect 21821 11237 21833 11271
rect 21867 11268 21879 11271
rect 22186 11268 22192 11280
rect 21867 11240 22192 11268
rect 21867 11237 21879 11240
rect 21821 11231 21879 11237
rect 22186 11228 22192 11240
rect 22244 11228 22250 11280
rect 14826 11160 14832 11212
rect 14884 11200 14890 11212
rect 15197 11203 15255 11209
rect 15197 11200 15209 11203
rect 14884 11172 15209 11200
rect 14884 11160 14890 11172
rect 15197 11169 15209 11172
rect 15243 11200 15255 11203
rect 15930 11200 15936 11212
rect 15243 11172 15936 11200
rect 15243 11169 15255 11172
rect 15197 11163 15255 11169
rect 15930 11160 15936 11172
rect 15988 11200 15994 11212
rect 16574 11200 16580 11212
rect 15988 11172 16580 11200
rect 15988 11160 15994 11172
rect 16574 11160 16580 11172
rect 16632 11200 16638 11212
rect 17129 11203 17187 11209
rect 17129 11200 17141 11203
rect 16632 11172 17141 11200
rect 16632 11160 16638 11172
rect 17129 11169 17141 11172
rect 17175 11169 17187 11203
rect 17129 11163 17187 11169
rect 20070 11160 20076 11212
rect 20128 11200 20134 11212
rect 20625 11208 20683 11209
rect 20456 11203 20683 11208
rect 20456 11200 20637 11203
rect 20128 11180 20637 11200
rect 20128 11172 20484 11180
rect 20128 11160 20134 11172
rect 13541 11135 13599 11141
rect 13541 11101 13553 11135
rect 13587 11101 13599 11135
rect 13541 11095 13599 11101
rect 13630 11092 13636 11144
rect 13688 11092 13694 11144
rect 13814 11092 13820 11144
rect 13872 11132 13878 11144
rect 13909 11135 13967 11141
rect 13909 11132 13921 11135
rect 13872 11104 13921 11132
rect 13872 11092 13878 11104
rect 13909 11101 13921 11104
rect 13955 11101 13967 11135
rect 13909 11095 13967 11101
rect 15562 11092 15568 11144
rect 15620 11092 15626 11144
rect 19886 11092 19892 11144
rect 19944 11132 19950 11144
rect 20165 11135 20223 11141
rect 20165 11132 20177 11135
rect 19944 11104 20177 11132
rect 19944 11092 19950 11104
rect 20165 11101 20177 11104
rect 20211 11101 20223 11135
rect 20165 11095 20223 11101
rect 20254 11092 20260 11144
rect 20312 11092 20318 11144
rect 20364 11141 20392 11172
rect 20625 11169 20637 11180
rect 20671 11169 20683 11203
rect 20625 11163 20683 11169
rect 21358 11160 21364 11212
rect 21416 11160 21422 11212
rect 21637 11203 21695 11209
rect 21637 11169 21649 11203
rect 21683 11200 21695 11203
rect 22278 11200 22284 11212
rect 21683 11172 22284 11200
rect 21683 11169 21695 11172
rect 21637 11163 21695 11169
rect 22278 11160 22284 11172
rect 22336 11160 22342 11212
rect 20349 11135 20407 11141
rect 20349 11101 20361 11135
rect 20395 11101 20407 11135
rect 20349 11095 20407 11101
rect 20438 11092 20444 11144
rect 20496 11092 20502 11144
rect 20898 11092 20904 11144
rect 20956 11092 20962 11144
rect 21453 11135 21511 11141
rect 21453 11101 21465 11135
rect 21499 11101 21511 11135
rect 21453 11095 21511 11101
rect 10229 11067 10287 11073
rect 10229 11064 10241 11067
rect 8404 11036 10241 11064
rect 10229 11033 10241 11036
rect 10275 11064 10287 11067
rect 10318 11064 10324 11076
rect 10275 11036 10324 11064
rect 10275 11033 10287 11036
rect 10229 11027 10287 11033
rect 10318 11024 10324 11036
rect 10376 11024 10382 11076
rect 10686 11024 10692 11076
rect 10744 11064 10750 11076
rect 10781 11067 10839 11073
rect 10781 11064 10793 11067
rect 10744 11036 10793 11064
rect 10744 11024 10750 11036
rect 10781 11033 10793 11036
rect 10827 11033 10839 11067
rect 10781 11027 10839 11033
rect 11422 11024 11428 11076
rect 11480 11064 11486 11076
rect 13081 11067 13139 11073
rect 13081 11064 13093 11067
rect 11480 11036 13093 11064
rect 11480 11024 11486 11036
rect 13081 11033 13093 11036
rect 13127 11064 13139 11067
rect 13725 11067 13783 11073
rect 13725 11064 13737 11067
rect 13127 11036 13737 11064
rect 13127 11033 13139 11036
rect 13081 11027 13139 11033
rect 13725 11033 13737 11036
rect 13771 11033 13783 11067
rect 13725 11027 13783 11033
rect 16390 11024 16396 11076
rect 16448 11024 16454 11076
rect 16991 11067 17049 11073
rect 16991 11033 17003 11067
rect 17037 11064 17049 11067
rect 17218 11064 17224 11076
rect 17037 11036 17224 11064
rect 17037 11033 17049 11036
rect 16991 11027 17049 11033
rect 17218 11024 17224 11036
rect 17276 11064 17282 11076
rect 17586 11064 17592 11076
rect 17276 11036 17592 11064
rect 17276 11024 17282 11036
rect 17586 11024 17592 11036
rect 17644 11024 17650 11076
rect 18874 11024 18880 11076
rect 18932 11064 18938 11076
rect 21468 11064 21496 11095
rect 21542 11092 21548 11144
rect 21600 11092 21606 11144
rect 22094 11092 22100 11144
rect 22152 11092 22158 11144
rect 22189 11135 22247 11141
rect 22189 11101 22201 11135
rect 22235 11101 22247 11135
rect 22189 11095 22247 11101
rect 22204 11064 22232 11095
rect 22370 11092 22376 11144
rect 22428 11092 22434 11144
rect 22480 11141 22508 11308
rect 22465 11135 22523 11141
rect 22465 11101 22477 11135
rect 22511 11101 22523 11135
rect 22465 11095 22523 11101
rect 22554 11064 22560 11076
rect 18932 11036 20484 11064
rect 21468 11036 22140 11064
rect 22204 11036 22560 11064
rect 18932 11024 18938 11036
rect 8300 11018 8352 11024
rect 20456 11008 20484 11036
rect 4304 10968 4660 10996
rect 4304 10956 4310 10968
rect 10870 10956 10876 11008
rect 10928 10996 10934 11008
rect 12894 10996 12900 11008
rect 10928 10968 12900 10996
rect 10928 10956 10934 10968
rect 12894 10956 12900 10968
rect 12952 10956 12958 11008
rect 13262 10956 13268 11008
rect 13320 10996 13326 11008
rect 13357 10999 13415 11005
rect 13357 10996 13369 10999
rect 13320 10968 13369 10996
rect 13320 10956 13326 10968
rect 13357 10965 13369 10968
rect 13403 10965 13415 10999
rect 13357 10959 13415 10965
rect 13906 10956 13912 11008
rect 13964 10996 13970 11008
rect 19334 10996 19340 11008
rect 13964 10968 19340 10996
rect 13964 10956 13970 10968
rect 19334 10956 19340 10968
rect 19392 10956 19398 11008
rect 20438 10956 20444 11008
rect 20496 10956 20502 11008
rect 22112 10996 22140 11036
rect 22554 11024 22560 11036
rect 22612 11024 22618 11076
rect 23014 11064 23020 11076
rect 22664 11036 23020 11064
rect 22664 10996 22692 11036
rect 23014 11024 23020 11036
rect 23072 11024 23078 11076
rect 22112 10968 22692 10996
rect 1104 10906 25208 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 25208 10906
rect 1104 10832 25208 10854
rect 8938 10792 8944 10804
rect 5460 10764 8944 10792
rect 5460 10733 5488 10764
rect 8938 10752 8944 10764
rect 8996 10752 9002 10804
rect 9030 10752 9036 10804
rect 9088 10792 9094 10804
rect 9171 10795 9229 10801
rect 9171 10792 9183 10795
rect 9088 10764 9183 10792
rect 9088 10752 9094 10764
rect 9171 10761 9183 10764
rect 9217 10792 9229 10795
rect 10870 10792 10876 10804
rect 9217 10764 10876 10792
rect 9217 10761 9229 10764
rect 9171 10755 9229 10761
rect 10870 10752 10876 10764
rect 10928 10752 10934 10804
rect 12894 10752 12900 10804
rect 12952 10792 12958 10804
rect 13814 10792 13820 10804
rect 12952 10764 13820 10792
rect 12952 10752 12958 10764
rect 13814 10752 13820 10764
rect 13872 10792 13878 10804
rect 14277 10795 14335 10801
rect 14277 10792 14289 10795
rect 13872 10764 14289 10792
rect 13872 10752 13878 10764
rect 14277 10761 14289 10764
rect 14323 10761 14335 10795
rect 14277 10755 14335 10761
rect 17126 10752 17132 10804
rect 17184 10752 17190 10804
rect 17586 10752 17592 10804
rect 17644 10752 17650 10804
rect 19886 10752 19892 10804
rect 19944 10792 19950 10804
rect 20898 10792 20904 10804
rect 19944 10764 20904 10792
rect 19944 10752 19950 10764
rect 20898 10752 20904 10764
rect 20956 10752 20962 10804
rect 21542 10752 21548 10804
rect 21600 10752 21606 10804
rect 22281 10795 22339 10801
rect 22281 10761 22293 10795
rect 22327 10792 22339 10795
rect 22370 10792 22376 10804
rect 22327 10764 22376 10792
rect 22327 10761 22339 10764
rect 22281 10755 22339 10761
rect 22370 10752 22376 10764
rect 22428 10752 22434 10804
rect 5445 10727 5503 10733
rect 5445 10693 5457 10727
rect 5491 10693 5503 10727
rect 5445 10687 5503 10693
rect 8294 10684 8300 10736
rect 8352 10684 8358 10736
rect 13633 10727 13691 10733
rect 13633 10724 13645 10727
rect 13280 10696 13645 10724
rect 13280 10668 13308 10696
rect 13633 10693 13645 10696
rect 13679 10724 13691 10727
rect 14185 10727 14243 10733
rect 14185 10724 14197 10727
rect 13679 10696 14197 10724
rect 13679 10693 13691 10696
rect 13633 10687 13691 10693
rect 14185 10693 14197 10696
rect 14231 10693 14243 10727
rect 21818 10724 21824 10736
rect 14185 10687 14243 10693
rect 21100 10696 21824 10724
rect 2774 10616 2780 10668
rect 2832 10616 2838 10668
rect 3053 10659 3111 10665
rect 3053 10625 3065 10659
rect 3099 10656 3111 10659
rect 3142 10656 3148 10668
rect 3099 10628 3148 10656
rect 3099 10625 3111 10628
rect 3053 10619 3111 10625
rect 3142 10616 3148 10628
rect 3200 10616 3206 10668
rect 6914 10616 6920 10668
rect 6972 10656 6978 10668
rect 7377 10659 7435 10665
rect 7377 10656 7389 10659
rect 6972 10628 7389 10656
rect 6972 10616 6978 10628
rect 7377 10625 7389 10628
rect 7423 10625 7435 10659
rect 13262 10656 13268 10668
rect 13223 10628 13268 10656
rect 7377 10619 7435 10625
rect 13262 10616 13268 10628
rect 13320 10616 13326 10668
rect 13354 10616 13360 10668
rect 13412 10616 13418 10668
rect 13446 10616 13452 10668
rect 13504 10616 13510 10668
rect 13722 10616 13728 10668
rect 13780 10616 13786 10668
rect 13814 10616 13820 10668
rect 13872 10616 13878 10668
rect 14093 10659 14151 10665
rect 14093 10625 14105 10659
rect 14139 10625 14151 10659
rect 14093 10619 14151 10625
rect 2961 10591 3019 10597
rect 2961 10557 2973 10591
rect 3007 10588 3019 10591
rect 3418 10588 3424 10600
rect 3007 10560 3424 10588
rect 3007 10557 3019 10560
rect 2961 10551 3019 10557
rect 3418 10548 3424 10560
rect 3476 10548 3482 10600
rect 3970 10548 3976 10600
rect 4028 10588 4034 10600
rect 4246 10588 4252 10600
rect 4028 10560 4252 10588
rect 4028 10548 4034 10560
rect 4246 10548 4252 10560
rect 4304 10548 4310 10600
rect 7742 10548 7748 10600
rect 7800 10548 7806 10600
rect 13464 10588 13492 10616
rect 14108 10588 14136 10619
rect 15930 10616 15936 10668
rect 15988 10616 15994 10668
rect 16758 10616 16764 10668
rect 16816 10656 16822 10668
rect 21100 10665 21128 10696
rect 21818 10684 21824 10696
rect 21876 10684 21882 10736
rect 17497 10659 17555 10665
rect 17497 10656 17509 10659
rect 16816 10628 17509 10656
rect 16816 10616 16822 10628
rect 17497 10625 17509 10628
rect 17543 10625 17555 10659
rect 17497 10619 17555 10625
rect 21085 10659 21143 10665
rect 21085 10625 21097 10659
rect 21131 10625 21143 10659
rect 21085 10619 21143 10625
rect 21266 10616 21272 10668
rect 21324 10616 21330 10668
rect 22462 10616 22468 10668
rect 22520 10616 22526 10668
rect 22649 10659 22707 10665
rect 22649 10625 22661 10659
rect 22695 10656 22707 10659
rect 23382 10656 23388 10668
rect 22695 10628 23388 10656
rect 22695 10625 22707 10628
rect 22649 10619 22707 10625
rect 23382 10616 23388 10628
rect 23440 10616 23446 10668
rect 13464 10560 14136 10588
rect 14461 10591 14519 10597
rect 14461 10557 14473 10591
rect 14507 10557 14519 10591
rect 14461 10551 14519 10557
rect 3510 10480 3516 10532
rect 3568 10520 3574 10532
rect 3568 10492 5396 10520
rect 3568 10480 3574 10492
rect 5368 10464 5396 10492
rect 12406 10492 13676 10520
rect 3053 10455 3111 10461
rect 3053 10421 3065 10455
rect 3099 10452 3111 10455
rect 3142 10452 3148 10464
rect 3099 10424 3148 10452
rect 3099 10421 3111 10424
rect 3053 10415 3111 10421
rect 3142 10412 3148 10424
rect 3200 10412 3206 10464
rect 3237 10455 3295 10461
rect 3237 10421 3249 10455
rect 3283 10452 3295 10455
rect 3326 10452 3332 10464
rect 3283 10424 3332 10452
rect 3283 10421 3295 10424
rect 3237 10415 3295 10421
rect 3326 10412 3332 10424
rect 3384 10412 3390 10464
rect 4154 10412 4160 10464
rect 4212 10452 4218 10464
rect 4614 10452 4620 10464
rect 4212 10424 4620 10452
rect 4212 10412 4218 10424
rect 4614 10412 4620 10424
rect 4672 10412 4678 10464
rect 5350 10412 5356 10464
rect 5408 10452 5414 10464
rect 12406 10452 12434 10492
rect 5408 10424 12434 10452
rect 13173 10455 13231 10461
rect 5408 10412 5414 10424
rect 13173 10421 13185 10455
rect 13219 10452 13231 10455
rect 13538 10452 13544 10464
rect 13219 10424 13544 10452
rect 13219 10421 13231 10424
rect 13173 10415 13231 10421
rect 13538 10412 13544 10424
rect 13596 10412 13602 10464
rect 13648 10452 13676 10492
rect 13722 10480 13728 10532
rect 13780 10520 13786 10532
rect 14476 10520 14504 10551
rect 17310 10548 17316 10600
rect 17368 10588 17374 10600
rect 17681 10591 17739 10597
rect 17681 10588 17693 10591
rect 17368 10560 17693 10588
rect 17368 10548 17374 10560
rect 17681 10557 17693 10560
rect 17727 10557 17739 10591
rect 17681 10551 17739 10557
rect 21542 10548 21548 10600
rect 21600 10548 21606 10600
rect 13780 10492 14504 10520
rect 13780 10480 13786 10492
rect 13906 10452 13912 10464
rect 13648 10424 13912 10452
rect 13906 10412 13912 10424
rect 13964 10412 13970 10464
rect 13998 10412 14004 10464
rect 14056 10412 14062 10464
rect 14366 10412 14372 10464
rect 14424 10452 14430 10464
rect 15194 10452 15200 10464
rect 14424 10424 15200 10452
rect 14424 10412 14430 10424
rect 15194 10412 15200 10424
rect 15252 10412 15258 10464
rect 21174 10412 21180 10464
rect 21232 10452 21238 10464
rect 21361 10455 21419 10461
rect 21361 10452 21373 10455
rect 21232 10424 21373 10452
rect 21232 10412 21238 10424
rect 21361 10421 21373 10424
rect 21407 10421 21419 10455
rect 21361 10415 21419 10421
rect 1104 10362 25208 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 25208 10362
rect 1104 10288 25208 10310
rect 3418 10208 3424 10260
rect 3476 10248 3482 10260
rect 4522 10248 4528 10260
rect 3476 10220 4528 10248
rect 3476 10208 3482 10220
rect 4522 10208 4528 10220
rect 4580 10248 4586 10260
rect 5258 10248 5264 10260
rect 4580 10220 5264 10248
rect 4580 10208 4586 10220
rect 5258 10208 5264 10220
rect 5316 10208 5322 10260
rect 17678 10208 17684 10260
rect 17736 10248 17742 10260
rect 17911 10251 17969 10257
rect 17911 10248 17923 10251
rect 17736 10220 17923 10248
rect 17736 10208 17742 10220
rect 17911 10217 17923 10220
rect 17957 10217 17969 10251
rect 17911 10211 17969 10217
rect 19886 10208 19892 10260
rect 19944 10208 19950 10260
rect 21729 10251 21787 10257
rect 21729 10217 21741 10251
rect 21775 10248 21787 10251
rect 21818 10248 21824 10260
rect 21775 10220 21824 10248
rect 21775 10217 21787 10220
rect 21729 10211 21787 10217
rect 21818 10208 21824 10220
rect 21876 10208 21882 10260
rect 2958 10140 2964 10192
rect 3016 10180 3022 10192
rect 3145 10183 3203 10189
rect 3145 10180 3157 10183
rect 3016 10152 3157 10180
rect 3016 10140 3022 10152
rect 3145 10149 3157 10152
rect 3191 10149 3203 10183
rect 3145 10143 3203 10149
rect 3237 10183 3295 10189
rect 3237 10149 3249 10183
rect 3283 10180 3295 10183
rect 3510 10180 3516 10192
rect 3283 10152 3516 10180
rect 3283 10149 3295 10152
rect 3237 10143 3295 10149
rect 3510 10140 3516 10152
rect 3568 10140 3574 10192
rect 3970 10140 3976 10192
rect 4028 10140 4034 10192
rect 4798 10180 4804 10192
rect 4080 10152 4804 10180
rect 1762 10072 1768 10124
rect 1820 10112 1826 10124
rect 2409 10115 2467 10121
rect 2409 10112 2421 10115
rect 1820 10084 2421 10112
rect 1820 10072 1826 10084
rect 2409 10081 2421 10084
rect 2455 10081 2467 10115
rect 4080 10112 4108 10152
rect 2409 10075 2467 10081
rect 3160 10084 4108 10112
rect 3160 10056 3188 10084
rect 4338 10072 4344 10124
rect 4396 10072 4402 10124
rect 2317 10047 2375 10053
rect 2317 10013 2329 10047
rect 2363 10013 2375 10047
rect 2317 10007 2375 10013
rect 2332 9976 2360 10007
rect 2866 10004 2872 10056
rect 2924 10044 2930 10056
rect 3053 10047 3111 10053
rect 3053 10044 3065 10047
rect 2924 10016 3065 10044
rect 2924 10004 2930 10016
rect 3053 10013 3065 10016
rect 3099 10013 3111 10047
rect 3053 10007 3111 10013
rect 3142 10004 3148 10056
rect 3200 10004 3206 10056
rect 3326 10004 3332 10056
rect 3384 10004 3390 10056
rect 4154 10004 4160 10056
rect 4212 10004 4218 10056
rect 4540 10054 4568 10152
rect 4798 10140 4804 10152
rect 4856 10140 4862 10192
rect 6086 10140 6092 10192
rect 6144 10180 6150 10192
rect 13909 10183 13967 10189
rect 6144 10152 12434 10180
rect 6144 10140 6150 10152
rect 6914 10072 6920 10124
rect 6972 10112 6978 10124
rect 7009 10115 7067 10121
rect 7009 10112 7021 10115
rect 6972 10084 7021 10112
rect 6972 10072 6978 10084
rect 7009 10081 7021 10084
rect 7055 10081 7067 10115
rect 7009 10075 7067 10081
rect 9306 10072 9312 10124
rect 9364 10112 9370 10124
rect 10045 10115 10103 10121
rect 10045 10112 10057 10115
rect 9364 10084 10057 10112
rect 9364 10072 9370 10084
rect 10045 10081 10057 10084
rect 10091 10081 10103 10115
rect 10045 10075 10103 10081
rect 10137 10115 10195 10121
rect 10137 10081 10149 10115
rect 10183 10081 10195 10115
rect 10137 10075 10195 10081
rect 4598 10057 4656 10063
rect 4598 10054 4610 10057
rect 4540 10026 4610 10054
rect 4598 10023 4610 10026
rect 4644 10023 4656 10057
rect 4598 10017 4656 10023
rect 4715 10047 4773 10053
rect 4715 10013 4727 10047
rect 4761 10013 4773 10047
rect 4715 10007 4773 10013
rect 4893 10047 4951 10053
rect 4893 10013 4905 10047
rect 4939 10044 4951 10047
rect 5442 10044 5448 10056
rect 4939 10016 5448 10044
rect 4939 10013 4951 10016
rect 4893 10007 4951 10013
rect 4724 9976 4752 10007
rect 5442 10004 5448 10016
rect 5500 10004 5506 10056
rect 6273 10047 6331 10053
rect 6273 10013 6285 10047
rect 6319 10044 6331 10047
rect 6546 10044 6552 10056
rect 6319 10016 6552 10044
rect 6319 10013 6331 10016
rect 6273 10007 6331 10013
rect 6546 10004 6552 10016
rect 6604 10004 6610 10056
rect 8757 10047 8815 10053
rect 8757 10013 8769 10047
rect 8803 10044 8815 10047
rect 8938 10044 8944 10056
rect 8803 10016 8944 10044
rect 8803 10013 8815 10016
rect 8757 10007 8815 10013
rect 8938 10004 8944 10016
rect 8996 10004 9002 10056
rect 9674 10004 9680 10056
rect 9732 10044 9738 10056
rect 10152 10044 10180 10075
rect 10502 10072 10508 10124
rect 10560 10112 10566 10124
rect 10873 10115 10931 10121
rect 10873 10112 10885 10115
rect 10560 10084 10885 10112
rect 10560 10072 10566 10084
rect 10873 10081 10885 10084
rect 10919 10081 10931 10115
rect 10873 10075 10931 10081
rect 10965 10115 11023 10121
rect 10965 10081 10977 10115
rect 11011 10081 11023 10115
rect 10965 10075 11023 10081
rect 10778 10044 10784 10056
rect 9732 10016 10784 10044
rect 9732 10004 9738 10016
rect 10778 10004 10784 10016
rect 10836 10044 10842 10056
rect 10980 10044 11008 10075
rect 10836 10016 11008 10044
rect 12406 10044 12434 10152
rect 13909 10149 13921 10183
rect 13955 10180 13967 10183
rect 16022 10180 16028 10192
rect 13955 10152 16028 10180
rect 13955 10149 13967 10152
rect 13909 10143 13967 10149
rect 16022 10140 16028 10152
rect 16080 10140 16086 10192
rect 19518 10180 19524 10192
rect 19260 10152 19524 10180
rect 13446 10072 13452 10124
rect 13504 10072 13510 10124
rect 13998 10072 14004 10124
rect 14056 10112 14062 10124
rect 14056 10084 14504 10112
rect 14056 10072 14062 10084
rect 13081 10047 13139 10053
rect 13081 10044 13093 10047
rect 12406 10016 13093 10044
rect 10836 10004 10842 10016
rect 13081 10013 13093 10016
rect 13127 10013 13139 10047
rect 13081 10007 13139 10013
rect 13265 10047 13323 10053
rect 13265 10013 13277 10047
rect 13311 10044 13323 10047
rect 13354 10044 13360 10056
rect 13311 10016 13360 10044
rect 13311 10013 13323 10016
rect 13265 10007 13323 10013
rect 2332 9948 3280 9976
rect 3252 9920 3280 9948
rect 4172 9948 4752 9976
rect 6457 9979 6515 9985
rect 4172 9920 4200 9948
rect 6457 9945 6469 9979
rect 6503 9976 6515 9979
rect 6638 9976 6644 9988
rect 6503 9948 6644 9976
rect 6503 9945 6515 9948
rect 6457 9939 6515 9945
rect 6638 9936 6644 9948
rect 6696 9936 6702 9988
rect 2130 9868 2136 9920
rect 2188 9868 2194 9920
rect 2777 9911 2835 9917
rect 2777 9877 2789 9911
rect 2823 9908 2835 9911
rect 2869 9911 2927 9917
rect 2869 9908 2881 9911
rect 2823 9880 2881 9908
rect 2823 9877 2835 9880
rect 2777 9871 2835 9877
rect 2869 9877 2881 9880
rect 2915 9877 2927 9911
rect 2869 9871 2927 9877
rect 3234 9868 3240 9920
rect 3292 9868 3298 9920
rect 4154 9868 4160 9920
rect 4212 9868 4218 9920
rect 4341 9911 4399 9917
rect 4341 9877 4353 9911
rect 4387 9908 4399 9911
rect 4706 9908 4712 9920
rect 4387 9880 4712 9908
rect 4387 9877 4399 9880
rect 4341 9871 4399 9877
rect 4706 9868 4712 9880
rect 4764 9868 4770 9920
rect 4801 9911 4859 9917
rect 4801 9877 4813 9911
rect 4847 9908 4859 9911
rect 4890 9908 4896 9920
rect 4847 9880 4896 9908
rect 4847 9877 4859 9880
rect 4801 9871 4859 9877
rect 4890 9868 4896 9880
rect 4948 9908 4954 9920
rect 7006 9908 7012 9920
rect 4948 9880 7012 9908
rect 4948 9868 4954 9880
rect 7006 9868 7012 9880
rect 7064 9868 7070 9920
rect 9306 9868 9312 9920
rect 9364 9908 9370 9920
rect 9585 9911 9643 9917
rect 9585 9908 9597 9911
rect 9364 9880 9597 9908
rect 9364 9868 9370 9880
rect 9585 9877 9597 9880
rect 9631 9877 9643 9911
rect 9585 9871 9643 9877
rect 9953 9911 10011 9917
rect 9953 9877 9965 9911
rect 9999 9908 10011 9911
rect 10134 9908 10140 9920
rect 9999 9880 10140 9908
rect 9999 9877 10011 9880
rect 9953 9871 10011 9877
rect 10134 9868 10140 9880
rect 10192 9868 10198 9920
rect 10410 9868 10416 9920
rect 10468 9868 10474 9920
rect 10781 9911 10839 9917
rect 10781 9877 10793 9911
rect 10827 9908 10839 9911
rect 11882 9908 11888 9920
rect 10827 9880 11888 9908
rect 10827 9877 10839 9880
rect 10781 9871 10839 9877
rect 11882 9868 11888 9880
rect 11940 9868 11946 9920
rect 13096 9908 13124 10007
rect 13354 10004 13360 10016
rect 13412 10004 13418 10056
rect 13538 10004 13544 10056
rect 13596 10004 13602 10056
rect 13906 10004 13912 10056
rect 13964 10044 13970 10056
rect 14093 10047 14151 10053
rect 14093 10044 14105 10047
rect 13964 10016 14105 10044
rect 13964 10004 13970 10016
rect 14093 10013 14105 10016
rect 14139 10013 14151 10047
rect 14093 10007 14151 10013
rect 14182 10004 14188 10056
rect 14240 10044 14246 10056
rect 14277 10047 14335 10053
rect 14277 10044 14289 10047
rect 14240 10016 14289 10044
rect 14240 10004 14246 10016
rect 14277 10013 14289 10016
rect 14323 10013 14335 10047
rect 14277 10007 14335 10013
rect 14366 10004 14372 10056
rect 14424 10004 14430 10056
rect 14476 10053 14504 10084
rect 15930 10072 15936 10124
rect 15988 10112 15994 10124
rect 16117 10115 16175 10121
rect 16117 10112 16129 10115
rect 15988 10084 16129 10112
rect 15988 10072 15994 10084
rect 16117 10081 16129 10084
rect 16163 10112 16175 10115
rect 16666 10112 16672 10124
rect 16163 10084 16672 10112
rect 16163 10081 16175 10084
rect 16117 10075 16175 10081
rect 16666 10072 16672 10084
rect 16724 10072 16730 10124
rect 17954 10072 17960 10124
rect 18012 10112 18018 10124
rect 18509 10115 18567 10121
rect 18509 10112 18521 10115
rect 18012 10084 18521 10112
rect 18012 10072 18018 10084
rect 18509 10081 18521 10084
rect 18555 10081 18567 10115
rect 18509 10075 18567 10081
rect 18598 10072 18604 10124
rect 18656 10072 18662 10124
rect 14461 10047 14519 10053
rect 14461 10013 14473 10047
rect 14507 10013 14519 10047
rect 14461 10007 14519 10013
rect 14737 10047 14795 10053
rect 14737 10013 14749 10047
rect 14783 10044 14795 10047
rect 15105 10047 15163 10053
rect 15105 10044 15117 10047
rect 14783 10016 15117 10044
rect 14783 10013 14795 10016
rect 14737 10007 14795 10013
rect 15105 10013 15117 10016
rect 15151 10013 15163 10047
rect 15105 10007 15163 10013
rect 15746 10004 15752 10056
rect 15804 10004 15810 10056
rect 16485 10047 16543 10053
rect 16485 10013 16497 10047
rect 16531 10044 16543 10047
rect 16574 10044 16580 10056
rect 16531 10016 16580 10044
rect 16531 10013 16543 10016
rect 16485 10007 16543 10013
rect 16574 10004 16580 10016
rect 16632 10004 16638 10056
rect 19260 10053 19288 10152
rect 19518 10140 19524 10152
rect 19576 10140 19582 10192
rect 20346 10140 20352 10192
rect 20404 10140 20410 10192
rect 22094 10140 22100 10192
rect 22152 10180 22158 10192
rect 22281 10183 22339 10189
rect 22281 10180 22293 10183
rect 22152 10152 22293 10180
rect 22152 10140 22158 10152
rect 22281 10149 22293 10152
rect 22327 10149 22339 10183
rect 22281 10143 22339 10149
rect 19337 10115 19395 10121
rect 19337 10081 19349 10115
rect 19383 10112 19395 10115
rect 20254 10112 20260 10124
rect 19383 10084 20260 10112
rect 19383 10081 19395 10084
rect 19337 10075 19395 10081
rect 20254 10072 20260 10084
rect 20312 10112 20318 10124
rect 20312 10084 20392 10112
rect 20312 10072 20318 10084
rect 19245 10047 19303 10053
rect 19245 10013 19257 10047
rect 19291 10013 19303 10047
rect 19245 10007 19303 10013
rect 19429 10047 19487 10053
rect 19429 10013 19441 10047
rect 19475 10013 19487 10047
rect 19429 10007 19487 10013
rect 13173 9979 13231 9985
rect 13173 9945 13185 9979
rect 13219 9976 13231 9979
rect 14200 9976 14228 10004
rect 14599 9979 14657 9985
rect 14599 9976 14611 9979
rect 13219 9948 14228 9976
rect 14292 9948 14611 9976
rect 13219 9945 13231 9948
rect 13173 9939 13231 9945
rect 14292 9908 14320 9948
rect 14599 9945 14611 9948
rect 14645 9976 14657 9979
rect 15838 9976 15844 9988
rect 14645 9948 15844 9976
rect 14645 9945 14657 9948
rect 14599 9939 14657 9945
rect 15838 9936 15844 9948
rect 15896 9936 15902 9988
rect 18417 9979 18475 9985
rect 17526 9948 18368 9976
rect 13096 9880 14320 9908
rect 15286 9868 15292 9920
rect 15344 9908 15350 9920
rect 16390 9908 16396 9920
rect 15344 9880 16396 9908
rect 15344 9868 15350 9880
rect 16390 9868 16396 9880
rect 16448 9908 16454 9920
rect 17604 9908 17632 9948
rect 16448 9880 17632 9908
rect 16448 9868 16454 9880
rect 17954 9868 17960 9920
rect 18012 9908 18018 9920
rect 18049 9911 18107 9917
rect 18049 9908 18061 9911
rect 18012 9880 18061 9908
rect 18012 9868 18018 9880
rect 18049 9877 18061 9880
rect 18095 9877 18107 9911
rect 18340 9908 18368 9948
rect 18417 9945 18429 9979
rect 18463 9976 18475 9979
rect 19444 9976 19472 10007
rect 19518 10004 19524 10056
rect 19576 10004 19582 10056
rect 19705 10047 19763 10053
rect 19705 10013 19717 10047
rect 19751 10013 19763 10047
rect 19705 10007 19763 10013
rect 19720 9976 19748 10007
rect 20070 10004 20076 10056
rect 20128 10004 20134 10056
rect 20364 10053 20392 10084
rect 20714 10072 20720 10124
rect 20772 10112 20778 10124
rect 22557 10115 22615 10121
rect 22557 10112 22569 10115
rect 20772 10084 22569 10112
rect 20772 10072 20778 10084
rect 22557 10081 22569 10084
rect 22603 10081 22615 10115
rect 22557 10075 22615 10081
rect 20349 10047 20407 10053
rect 20349 10013 20361 10047
rect 20395 10013 20407 10047
rect 20349 10007 20407 10013
rect 20438 10004 20444 10056
rect 20496 10004 20502 10056
rect 22646 10004 22652 10056
rect 22704 10004 22710 10056
rect 19794 9976 19800 9988
rect 18463 9948 19800 9976
rect 18463 9945 18475 9948
rect 18417 9939 18475 9945
rect 19794 9936 19800 9948
rect 19852 9936 19858 9988
rect 18782 9908 18788 9920
rect 18340 9880 18788 9908
rect 18049 9871 18107 9877
rect 18782 9868 18788 9880
rect 18840 9868 18846 9920
rect 20162 9868 20168 9920
rect 20220 9868 20226 9920
rect 1104 9818 25208 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 25208 9818
rect 1104 9744 25208 9766
rect 4338 9664 4344 9716
rect 4396 9704 4402 9716
rect 4433 9707 4491 9713
rect 4433 9704 4445 9707
rect 4396 9676 4445 9704
rect 4396 9664 4402 9676
rect 4433 9673 4445 9676
rect 4479 9673 4491 9707
rect 4433 9667 4491 9673
rect 4890 9664 4896 9716
rect 4948 9704 4954 9716
rect 5350 9704 5356 9716
rect 4948 9676 5356 9704
rect 4948 9664 4954 9676
rect 5350 9664 5356 9676
rect 5408 9664 5414 9716
rect 6546 9664 6552 9716
rect 6604 9664 6610 9716
rect 8389 9707 8447 9713
rect 8389 9673 8401 9707
rect 8435 9704 8447 9707
rect 9030 9704 9036 9716
rect 8435 9676 9036 9704
rect 8435 9673 8447 9676
rect 8389 9667 8447 9673
rect 9030 9664 9036 9676
rect 9088 9664 9094 9716
rect 10778 9664 10784 9716
rect 10836 9704 10842 9716
rect 10836 9676 11008 9704
rect 10836 9664 10842 9676
rect 2774 9596 2780 9648
rect 2832 9636 2838 9648
rect 2869 9639 2927 9645
rect 2869 9636 2881 9639
rect 2832 9608 2881 9636
rect 2832 9596 2838 9608
rect 2869 9605 2881 9608
rect 2915 9636 2927 9639
rect 3605 9639 3663 9645
rect 3605 9636 3617 9639
rect 2915 9608 3617 9636
rect 2915 9605 2927 9608
rect 2869 9599 2927 9605
rect 3605 9605 3617 9608
rect 3651 9605 3663 9639
rect 4356 9636 4384 9664
rect 4617 9639 4675 9645
rect 4617 9636 4629 9639
rect 3605 9599 3663 9605
rect 3804 9608 4384 9636
rect 4540 9608 4629 9636
rect 3326 9528 3332 9580
rect 3384 9528 3390 9580
rect 3804 9577 3832 9608
rect 3789 9571 3847 9577
rect 3789 9537 3801 9571
rect 3835 9537 3847 9571
rect 3789 9531 3847 9537
rect 4065 9571 4123 9577
rect 4065 9537 4077 9571
rect 4111 9568 4123 9571
rect 4154 9568 4160 9580
rect 4111 9540 4160 9568
rect 4111 9537 4123 9540
rect 4065 9531 4123 9537
rect 4154 9528 4160 9540
rect 4212 9528 4218 9580
rect 4540 9577 4568 9608
rect 4617 9605 4629 9608
rect 4663 9636 4675 9639
rect 5534 9636 5540 9648
rect 4663 9608 5540 9636
rect 4663 9605 4675 9608
rect 4617 9599 4675 9605
rect 5534 9596 5540 9608
rect 5592 9596 5598 9648
rect 6454 9596 6460 9648
rect 6512 9596 6518 9648
rect 6564 9636 6592 9664
rect 6564 9608 6684 9636
rect 4249 9571 4307 9577
rect 4249 9537 4261 9571
rect 4295 9537 4307 9571
rect 4249 9531 4307 9537
rect 4341 9571 4399 9577
rect 4341 9537 4353 9571
rect 4387 9537 4399 9571
rect 4341 9531 4399 9537
rect 4525 9571 4583 9577
rect 4525 9537 4537 9571
rect 4571 9537 4583 9571
rect 4525 9531 4583 9537
rect 3237 9503 3295 9509
rect 3237 9469 3249 9503
rect 3283 9500 3295 9503
rect 3970 9500 3976 9512
rect 3283 9472 3976 9500
rect 3283 9469 3295 9472
rect 3237 9463 3295 9469
rect 3970 9460 3976 9472
rect 4028 9460 4034 9512
rect 4264 9432 4292 9531
rect 4356 9500 4384 9531
rect 4798 9528 4804 9580
rect 4856 9568 4862 9580
rect 4893 9571 4951 9577
rect 4893 9568 4905 9571
rect 4856 9540 4905 9568
rect 4856 9528 4862 9540
rect 4893 9537 4905 9540
rect 4939 9537 4951 9571
rect 4893 9531 4951 9537
rect 5166 9528 5172 9580
rect 5224 9528 5230 9580
rect 5258 9528 5264 9580
rect 5316 9568 5322 9580
rect 5353 9571 5411 9577
rect 5353 9568 5365 9571
rect 5316 9540 5365 9568
rect 5316 9528 5322 9540
rect 5353 9537 5365 9540
rect 5399 9537 5411 9571
rect 5353 9531 5411 9537
rect 5905 9571 5963 9577
rect 5905 9537 5917 9571
rect 5951 9568 5963 9571
rect 6362 9568 6368 9580
rect 5951 9540 6368 9568
rect 5951 9537 5963 9540
rect 5905 9531 5963 9537
rect 6362 9528 6368 9540
rect 6420 9528 6426 9580
rect 6472 9568 6500 9596
rect 6549 9571 6607 9577
rect 6549 9568 6561 9571
rect 6472 9540 6561 9568
rect 6549 9537 6561 9540
rect 6595 9537 6607 9571
rect 6656 9568 6684 9608
rect 6914 9596 6920 9648
rect 6972 9636 6978 9648
rect 8018 9636 8024 9648
rect 6972 9608 8024 9636
rect 6972 9596 6978 9608
rect 8018 9596 8024 9608
rect 8076 9636 8082 9648
rect 8076 9608 9536 9636
rect 8076 9596 8082 9608
rect 9508 9577 9536 9608
rect 10226 9596 10232 9648
rect 10284 9596 10290 9648
rect 10980 9636 11008 9676
rect 14182 9664 14188 9716
rect 14240 9704 14246 9716
rect 15657 9707 15715 9713
rect 14240 9676 15056 9704
rect 14240 9664 14246 9676
rect 10980 9608 11836 9636
rect 7009 9571 7067 9577
rect 7009 9568 7021 9571
rect 6656 9540 7021 9568
rect 6549 9531 6607 9537
rect 7009 9537 7021 9540
rect 7055 9537 7067 9571
rect 7009 9531 7067 9537
rect 7193 9571 7251 9577
rect 7193 9537 7205 9571
rect 7239 9537 7251 9571
rect 9493 9571 9551 9577
rect 7193 9531 7251 9537
rect 7300 9540 8616 9568
rect 4709 9503 4767 9509
rect 4709 9500 4721 9503
rect 4356 9472 4721 9500
rect 4709 9469 4721 9472
rect 4755 9500 4767 9503
rect 5184 9500 5212 9528
rect 4755 9472 5028 9500
rect 5184 9472 6224 9500
rect 4755 9469 4767 9472
rect 4709 9463 4767 9469
rect 4798 9432 4804 9444
rect 4264 9404 4804 9432
rect 4798 9392 4804 9404
rect 4856 9392 4862 9444
rect 5000 9432 5028 9472
rect 5442 9432 5448 9444
rect 5000 9404 5448 9432
rect 5442 9392 5448 9404
rect 5500 9392 5506 9444
rect 6196 9432 6224 9472
rect 6270 9460 6276 9512
rect 6328 9500 6334 9512
rect 6457 9503 6515 9509
rect 6457 9500 6469 9503
rect 6328 9472 6469 9500
rect 6328 9460 6334 9472
rect 6457 9469 6469 9472
rect 6503 9469 6515 9503
rect 6457 9463 6515 9469
rect 6638 9460 6644 9512
rect 6696 9500 6702 9512
rect 7208 9500 7236 9531
rect 6696 9472 7236 9500
rect 6696 9460 6702 9472
rect 7300 9432 7328 9540
rect 7377 9503 7435 9509
rect 7377 9469 7389 9503
rect 7423 9500 7435 9503
rect 7423 9472 8432 9500
rect 7423 9469 7435 9472
rect 7377 9463 7435 9469
rect 6196 9404 7328 9432
rect 7742 9392 7748 9444
rect 7800 9432 7806 9444
rect 8021 9435 8079 9441
rect 8021 9432 8033 9435
rect 7800 9404 8033 9432
rect 7800 9392 7806 9404
rect 8021 9401 8033 9404
rect 8067 9401 8079 9435
rect 8021 9395 8079 9401
rect 3234 9324 3240 9376
rect 3292 9324 3298 9376
rect 3326 9324 3332 9376
rect 3384 9364 3390 9376
rect 3513 9367 3571 9373
rect 3513 9364 3525 9367
rect 3384 9336 3525 9364
rect 3384 9324 3390 9336
rect 3513 9333 3525 9336
rect 3559 9333 3571 9367
rect 3513 9327 3571 9333
rect 4522 9324 4528 9376
rect 4580 9364 4586 9376
rect 4617 9367 4675 9373
rect 4617 9364 4629 9367
rect 4580 9336 4629 9364
rect 4580 9324 4586 9336
rect 4617 9333 4629 9336
rect 4663 9333 4675 9367
rect 4617 9327 4675 9333
rect 5077 9367 5135 9373
rect 5077 9333 5089 9367
rect 5123 9364 5135 9367
rect 5902 9364 5908 9376
rect 5123 9336 5908 9364
rect 5123 9333 5135 9336
rect 5077 9327 5135 9333
rect 5902 9324 5908 9336
rect 5960 9324 5966 9376
rect 6825 9367 6883 9373
rect 6825 9333 6837 9367
rect 6871 9364 6883 9367
rect 7926 9364 7932 9376
rect 6871 9336 7932 9364
rect 6871 9333 6883 9336
rect 6825 9327 6883 9333
rect 7926 9324 7932 9336
rect 7984 9324 7990 9376
rect 8404 9364 8432 9472
rect 8478 9460 8484 9512
rect 8536 9460 8542 9512
rect 8588 9509 8616 9540
rect 9493 9537 9505 9571
rect 9539 9537 9551 9571
rect 9493 9531 9551 9537
rect 11287 9571 11345 9577
rect 11287 9537 11299 9571
rect 11333 9568 11345 9571
rect 11333 9540 11744 9568
rect 11333 9537 11345 9540
rect 11287 9531 11345 9537
rect 8573 9503 8631 9509
rect 8573 9469 8585 9503
rect 8619 9469 8631 9503
rect 8573 9463 8631 9469
rect 9861 9503 9919 9509
rect 9861 9469 9873 9503
rect 9907 9500 9919 9503
rect 9907 9472 11560 9500
rect 9907 9469 9919 9472
rect 9861 9463 9919 9469
rect 11532 9441 11560 9472
rect 11517 9435 11575 9441
rect 11164 9404 11468 9432
rect 11164 9364 11192 9404
rect 8404 9336 11192 9364
rect 11440 9364 11468 9404
rect 11517 9401 11529 9435
rect 11563 9401 11575 9435
rect 11716 9432 11744 9540
rect 11808 9500 11836 9608
rect 11974 9596 11980 9648
rect 12032 9596 12038 9648
rect 13630 9636 13636 9648
rect 12406 9608 13636 9636
rect 11885 9571 11943 9577
rect 11885 9537 11897 9571
rect 11931 9568 11943 9571
rect 12158 9568 12164 9580
rect 11931 9540 12164 9568
rect 11931 9537 11943 9540
rect 11885 9531 11943 9537
rect 12158 9528 12164 9540
rect 12216 9528 12222 9580
rect 12069 9503 12127 9509
rect 12069 9500 12081 9503
rect 11808 9472 12081 9500
rect 12069 9469 12081 9472
rect 12115 9469 12127 9503
rect 12069 9463 12127 9469
rect 12158 9432 12164 9444
rect 11716 9404 12164 9432
rect 11517 9395 11575 9401
rect 12158 9392 12164 9404
rect 12216 9392 12222 9444
rect 12406 9364 12434 9608
rect 13630 9596 13636 9608
rect 13688 9596 13694 9648
rect 15028 9636 15056 9676
rect 15657 9673 15669 9707
rect 15703 9673 15715 9707
rect 15657 9667 15715 9673
rect 15672 9636 15700 9667
rect 16574 9664 16580 9716
rect 16632 9704 16638 9716
rect 16669 9707 16727 9713
rect 16669 9704 16681 9707
rect 16632 9676 16681 9704
rect 16632 9664 16638 9676
rect 16669 9673 16681 9676
rect 16715 9673 16727 9707
rect 16669 9667 16727 9673
rect 17129 9707 17187 9713
rect 17129 9673 17141 9707
rect 17175 9704 17187 9707
rect 17586 9704 17592 9716
rect 17175 9676 17592 9704
rect 17175 9673 17187 9676
rect 17129 9667 17187 9673
rect 17586 9664 17592 9676
rect 17644 9664 17650 9716
rect 19705 9707 19763 9713
rect 19705 9673 19717 9707
rect 19751 9704 19763 9707
rect 20162 9704 20168 9716
rect 19751 9676 20168 9704
rect 19751 9673 19763 9676
rect 19705 9667 19763 9673
rect 20162 9664 20168 9676
rect 20220 9664 20226 9716
rect 21266 9704 21272 9716
rect 20548 9676 21272 9704
rect 13541 9571 13599 9577
rect 13541 9537 13553 9571
rect 13587 9568 13599 9571
rect 14936 9568 14964 9622
rect 15028 9608 15700 9636
rect 16960 9608 17632 9636
rect 15102 9568 15108 9580
rect 13587 9540 14044 9568
rect 14936 9540 15108 9568
rect 13587 9537 13599 9540
rect 13541 9531 13599 9537
rect 13906 9460 13912 9512
rect 13964 9460 13970 9512
rect 14016 9500 14044 9540
rect 15102 9528 15108 9540
rect 15160 9528 15166 9580
rect 15194 9528 15200 9580
rect 15252 9568 15258 9580
rect 15598 9571 15656 9577
rect 15598 9568 15610 9571
rect 15252 9540 15610 9568
rect 15252 9528 15258 9540
rect 15598 9537 15610 9540
rect 15644 9537 15656 9571
rect 16960 9568 16988 9608
rect 15598 9531 15656 9537
rect 16040 9540 16988 9568
rect 17037 9571 17095 9577
rect 14274 9500 14280 9512
rect 14016 9472 14280 9500
rect 14274 9460 14280 9472
rect 14332 9460 14338 9512
rect 15335 9503 15393 9509
rect 15335 9469 15347 9503
rect 15381 9500 15393 9503
rect 15746 9500 15752 9512
rect 15381 9472 15752 9500
rect 15381 9469 15393 9472
rect 15335 9463 15393 9469
rect 15746 9460 15752 9472
rect 15804 9500 15810 9512
rect 16040 9500 16068 9540
rect 17037 9537 17049 9571
rect 17083 9537 17095 9571
rect 17037 9531 17095 9537
rect 15804 9472 16068 9500
rect 15804 9460 15810 9472
rect 16114 9460 16120 9512
rect 16172 9460 16178 9512
rect 17052 9432 17080 9531
rect 17494 9528 17500 9580
rect 17552 9528 17558 9580
rect 17604 9568 17632 9608
rect 18782 9596 18788 9648
rect 18840 9596 18846 9648
rect 19291 9639 19349 9645
rect 19291 9605 19303 9639
rect 19337 9636 19349 9639
rect 19981 9639 20039 9645
rect 19337 9608 19840 9636
rect 19337 9605 19349 9608
rect 19291 9599 19349 9605
rect 19812 9580 19840 9608
rect 19981 9605 19993 9639
rect 20027 9636 20039 9639
rect 20548 9636 20576 9676
rect 21266 9664 21272 9676
rect 21324 9664 21330 9716
rect 20027 9608 20576 9636
rect 20027 9605 20039 9608
rect 19981 9599 20039 9605
rect 17604 9540 18000 9568
rect 17218 9460 17224 9512
rect 17276 9460 17282 9512
rect 17865 9503 17923 9509
rect 17865 9500 17877 9503
rect 17512 9472 17877 9500
rect 14660 9404 17080 9432
rect 11440 9336 12434 9364
rect 12894 9324 12900 9376
rect 12952 9364 12958 9376
rect 14660 9364 14688 9404
rect 12952 9336 14688 9364
rect 12952 9324 12958 9336
rect 15470 9324 15476 9376
rect 15528 9324 15534 9376
rect 15930 9324 15936 9376
rect 15988 9364 15994 9376
rect 16025 9367 16083 9373
rect 16025 9364 16037 9367
rect 15988 9336 16037 9364
rect 15988 9324 15994 9336
rect 16025 9333 16037 9336
rect 16071 9333 16083 9367
rect 17512 9364 17540 9472
rect 17865 9469 17877 9472
rect 17911 9469 17923 9503
rect 17972 9500 18000 9540
rect 19518 9528 19524 9580
rect 19576 9568 19582 9580
rect 19613 9571 19671 9577
rect 19613 9568 19625 9571
rect 19576 9540 19625 9568
rect 19576 9528 19582 9540
rect 19613 9537 19625 9540
rect 19659 9537 19671 9571
rect 19613 9531 19671 9537
rect 19794 9528 19800 9580
rect 19852 9528 19858 9580
rect 19886 9528 19892 9580
rect 19944 9528 19950 9580
rect 20070 9528 20076 9580
rect 20128 9528 20134 9580
rect 20254 9528 20260 9580
rect 20312 9568 20318 9580
rect 20349 9571 20407 9577
rect 20349 9568 20361 9571
rect 20312 9540 20361 9568
rect 20312 9528 20318 9540
rect 20349 9537 20361 9540
rect 20395 9537 20407 9571
rect 20548 9568 20576 9608
rect 20625 9639 20683 9645
rect 20625 9605 20637 9639
rect 20671 9636 20683 9639
rect 20671 9608 20944 9636
rect 20671 9605 20683 9608
rect 20625 9599 20683 9605
rect 20916 9577 20944 9608
rect 20717 9571 20775 9577
rect 20717 9568 20729 9571
rect 20548 9540 20729 9568
rect 20349 9531 20407 9537
rect 20717 9537 20729 9540
rect 20763 9537 20775 9571
rect 20717 9531 20775 9537
rect 20901 9571 20959 9577
rect 20901 9537 20913 9571
rect 20947 9537 20959 9571
rect 20901 9531 20959 9537
rect 20088 9500 20116 9528
rect 17972 9472 20116 9500
rect 17865 9463 17923 9469
rect 20622 9460 20628 9512
rect 20680 9460 20686 9512
rect 20916 9500 20944 9531
rect 21174 9528 21180 9580
rect 21232 9528 21238 9580
rect 21284 9568 21312 9664
rect 21361 9639 21419 9645
rect 21361 9605 21373 9639
rect 21407 9636 21419 9639
rect 22646 9636 22652 9648
rect 21407 9608 22652 9636
rect 21407 9605 21419 9608
rect 21361 9599 21419 9605
rect 22646 9596 22652 9608
rect 22704 9596 22710 9648
rect 21821 9571 21879 9577
rect 21284 9540 21680 9568
rect 21542 9500 21548 9512
rect 20916 9472 21548 9500
rect 21542 9460 21548 9472
rect 21600 9460 21606 9512
rect 21652 9500 21680 9540
rect 21821 9537 21833 9571
rect 21867 9568 21879 9571
rect 21867 9540 22048 9568
rect 21867 9537 21879 9540
rect 21821 9531 21879 9537
rect 21913 9503 21971 9509
rect 21913 9500 21925 9503
rect 21652 9472 21925 9500
rect 21913 9469 21925 9472
rect 21959 9469 21971 9503
rect 21913 9463 21971 9469
rect 20346 9392 20352 9444
rect 20404 9432 20410 9444
rect 20441 9435 20499 9441
rect 20441 9432 20453 9435
rect 20404 9404 20453 9432
rect 20404 9392 20410 9404
rect 20441 9401 20453 9404
rect 20487 9432 20499 9435
rect 20990 9432 20996 9444
rect 20487 9404 20996 9432
rect 20487 9401 20499 9404
rect 20441 9395 20499 9401
rect 20990 9392 20996 9404
rect 21048 9392 21054 9444
rect 21174 9392 21180 9444
rect 21232 9432 21238 9444
rect 22020 9432 22048 9540
rect 21232 9404 22048 9432
rect 22189 9435 22247 9441
rect 21232 9392 21238 9404
rect 22189 9401 22201 9435
rect 22235 9432 22247 9435
rect 22278 9432 22284 9444
rect 22235 9404 22284 9432
rect 22235 9401 22247 9404
rect 22189 9395 22247 9401
rect 22278 9392 22284 9404
rect 22336 9392 22342 9444
rect 17862 9364 17868 9376
rect 17512 9336 17868 9364
rect 16025 9327 16083 9333
rect 17862 9324 17868 9336
rect 17920 9324 17926 9376
rect 18046 9324 18052 9376
rect 18104 9364 18110 9376
rect 19886 9364 19892 9376
rect 18104 9336 19892 9364
rect 18104 9324 18110 9336
rect 19886 9324 19892 9336
rect 19944 9324 19950 9376
rect 21542 9324 21548 9376
rect 21600 9364 21606 9376
rect 21821 9367 21879 9373
rect 21821 9364 21833 9367
rect 21600 9336 21833 9364
rect 21600 9324 21606 9336
rect 21821 9333 21833 9336
rect 21867 9333 21879 9367
rect 21821 9327 21879 9333
rect 1104 9274 25208 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 25208 9274
rect 1104 9200 25208 9222
rect 4430 9120 4436 9172
rect 4488 9160 4494 9172
rect 4798 9160 4804 9172
rect 4488 9132 4804 9160
rect 4488 9120 4494 9132
rect 4798 9120 4804 9132
rect 4856 9120 4862 9172
rect 6086 9120 6092 9172
rect 6144 9120 6150 9172
rect 6270 9120 6276 9172
rect 6328 9120 6334 9172
rect 10226 9120 10232 9172
rect 10284 9160 10290 9172
rect 10962 9160 10968 9172
rect 10284 9132 10968 9160
rect 10284 9120 10290 9132
rect 10962 9120 10968 9132
rect 11020 9120 11026 9172
rect 11882 9120 11888 9172
rect 11940 9160 11946 9172
rect 12023 9163 12081 9169
rect 12023 9160 12035 9163
rect 11940 9132 12035 9160
rect 11940 9120 11946 9132
rect 12023 9129 12035 9132
rect 12069 9160 12081 9163
rect 12342 9160 12348 9172
rect 12069 9132 12348 9160
rect 12069 9129 12081 9132
rect 12023 9123 12081 9129
rect 12342 9120 12348 9132
rect 12400 9120 12406 9172
rect 13630 9120 13636 9172
rect 13688 9160 13694 9172
rect 15378 9160 15384 9172
rect 13688 9132 15384 9160
rect 13688 9120 13694 9132
rect 15378 9120 15384 9132
rect 15436 9160 15442 9172
rect 15930 9160 15936 9172
rect 15436 9132 15936 9160
rect 15436 9120 15442 9132
rect 15930 9120 15936 9132
rect 15988 9120 15994 9172
rect 16114 9120 16120 9172
rect 16172 9160 16178 9172
rect 16807 9163 16865 9169
rect 16807 9160 16819 9163
rect 16172 9132 16819 9160
rect 16172 9120 16178 9132
rect 16807 9129 16819 9132
rect 16853 9160 16865 9163
rect 16853 9132 19380 9160
rect 16853 9129 16865 9132
rect 16807 9123 16865 9129
rect 4985 9095 5043 9101
rect 3436 9064 4936 9092
rect 3050 8984 3056 9036
rect 3108 9024 3114 9036
rect 3108 8996 3372 9024
rect 3108 8984 3114 8996
rect 2774 8916 2780 8968
rect 2832 8956 2838 8968
rect 3344 8965 3372 8996
rect 3436 8965 3464 9064
rect 3513 9027 3571 9033
rect 3513 8993 3525 9027
rect 3559 9024 3571 9027
rect 3789 9027 3847 9033
rect 3789 9024 3801 9027
rect 3559 8996 3801 9024
rect 3559 8993 3571 8996
rect 3513 8987 3571 8993
rect 3789 8993 3801 8996
rect 3835 9024 3847 9027
rect 4062 9024 4068 9036
rect 3835 8996 4068 9024
rect 3835 8993 3847 8996
rect 3789 8987 3847 8993
rect 4062 8984 4068 8996
rect 4120 8984 4126 9036
rect 4338 8984 4344 9036
rect 4396 9024 4402 9036
rect 4617 9027 4675 9033
rect 4617 9024 4629 9027
rect 4396 8996 4629 9024
rect 4396 8984 4402 8996
rect 4617 8993 4629 8996
rect 4663 9024 4675 9027
rect 4798 9024 4804 9036
rect 4663 8996 4804 9024
rect 4663 8993 4675 8996
rect 4617 8987 4675 8993
rect 4798 8984 4804 8996
rect 4856 8984 4862 9036
rect 2869 8959 2927 8965
rect 2869 8956 2881 8959
rect 2832 8928 2881 8956
rect 2832 8916 2838 8928
rect 2869 8925 2881 8928
rect 2915 8925 2927 8959
rect 2869 8919 2927 8925
rect 3145 8959 3203 8965
rect 3145 8925 3157 8959
rect 3191 8925 3203 8959
rect 3145 8919 3203 8925
rect 3329 8959 3387 8965
rect 3329 8925 3341 8959
rect 3375 8925 3387 8959
rect 3329 8919 3387 8925
rect 3421 8959 3479 8965
rect 3421 8925 3433 8959
rect 3467 8925 3479 8959
rect 3421 8919 3479 8925
rect 2498 8780 2504 8832
rect 2556 8820 2562 8832
rect 2685 8823 2743 8829
rect 2685 8820 2697 8823
rect 2556 8792 2697 8820
rect 2556 8780 2562 8792
rect 2685 8789 2697 8792
rect 2731 8789 2743 8823
rect 3160 8820 3188 8919
rect 3436 8888 3464 8919
rect 3602 8916 3608 8968
rect 3660 8916 3666 8968
rect 4157 8959 4215 8965
rect 4157 8925 4169 8959
rect 4203 8956 4215 8959
rect 4706 8956 4712 8968
rect 4203 8928 4712 8956
rect 4203 8925 4215 8928
rect 4157 8919 4215 8925
rect 4706 8916 4712 8928
rect 4764 8916 4770 8968
rect 4908 8965 4936 9064
rect 4985 9061 4997 9095
rect 5031 9092 5043 9095
rect 5534 9092 5540 9104
rect 5031 9064 5540 9092
rect 5031 9061 5043 9064
rect 4985 9055 5043 9061
rect 5534 9052 5540 9064
rect 5592 9092 5598 9104
rect 6638 9092 6644 9104
rect 5592 9064 6644 9092
rect 5592 9052 5598 9064
rect 6638 9052 6644 9064
rect 6696 9052 6702 9104
rect 9582 9092 9588 9104
rect 9416 9064 9588 9092
rect 5626 9024 5632 9036
rect 5092 8996 5632 9024
rect 5092 8965 5120 8996
rect 5626 8984 5632 8996
rect 5684 8984 5690 9036
rect 5718 8984 5724 9036
rect 5776 9024 5782 9036
rect 6549 9027 6607 9033
rect 6549 9024 6561 9027
rect 5776 8996 6561 9024
rect 5776 8984 5782 8996
rect 6549 8993 6561 8996
rect 6595 8993 6607 9027
rect 6549 8987 6607 8993
rect 8018 8984 8024 9036
rect 8076 9024 8082 9036
rect 9416 9033 9444 9064
rect 9582 9052 9588 9064
rect 9640 9052 9646 9104
rect 12805 9095 12863 9101
rect 12805 9061 12817 9095
rect 12851 9061 12863 9095
rect 12805 9055 12863 9061
rect 8297 9027 8355 9033
rect 8297 9024 8309 9027
rect 8076 8996 8309 9024
rect 8076 8984 8082 8996
rect 8297 8993 8309 8996
rect 8343 8993 8355 9027
rect 8297 8987 8355 8993
rect 9401 9027 9459 9033
rect 9401 8993 9413 9027
rect 9447 8993 9459 9027
rect 9401 8987 9459 8993
rect 9493 9027 9551 9033
rect 9493 8993 9505 9027
rect 9539 9024 9551 9027
rect 9674 9024 9680 9036
rect 9539 8996 9680 9024
rect 9539 8993 9551 8996
rect 9493 8987 9551 8993
rect 4893 8959 4951 8965
rect 4893 8925 4905 8959
rect 4939 8925 4951 8959
rect 4893 8919 4951 8925
rect 5077 8959 5135 8965
rect 5077 8925 5089 8959
rect 5123 8925 5135 8959
rect 5077 8919 5135 8925
rect 5169 8959 5227 8965
rect 5169 8925 5181 8959
rect 5215 8956 5227 8959
rect 5258 8956 5264 8968
rect 5215 8928 5264 8956
rect 5215 8925 5227 8928
rect 5169 8919 5227 8925
rect 5258 8916 5264 8928
rect 5316 8916 5322 8968
rect 5350 8916 5356 8968
rect 5408 8916 5414 8968
rect 5445 8959 5503 8965
rect 5445 8925 5457 8959
rect 5491 8925 5503 8959
rect 5445 8919 5503 8925
rect 3510 8888 3516 8900
rect 3436 8860 3516 8888
rect 3510 8848 3516 8860
rect 3568 8848 3574 8900
rect 3988 8860 4200 8888
rect 3418 8820 3424 8832
rect 3160 8792 3424 8820
rect 2685 8783 2743 8789
rect 3418 8780 3424 8792
rect 3476 8780 3482 8832
rect 3786 8780 3792 8832
rect 3844 8780 3850 8832
rect 3988 8829 4016 8860
rect 3973 8823 4031 8829
rect 3973 8789 3985 8823
rect 4019 8789 4031 8823
rect 3973 8783 4031 8789
rect 4062 8780 4068 8832
rect 4120 8780 4126 8832
rect 4172 8820 4200 8860
rect 4246 8848 4252 8900
rect 4304 8848 4310 8900
rect 4430 8848 4436 8900
rect 4488 8848 4494 8900
rect 4798 8848 4804 8900
rect 4856 8888 4862 8900
rect 5460 8888 5488 8919
rect 5534 8916 5540 8968
rect 5592 8916 5598 8968
rect 8312 8956 8340 8987
rect 9674 8984 9680 8996
rect 9732 8984 9738 9036
rect 10410 8984 10416 9036
rect 10468 9024 10474 9036
rect 10597 9027 10655 9033
rect 10597 9024 10609 9027
rect 10468 8996 10609 9024
rect 10468 8984 10474 8996
rect 10597 8993 10609 8996
rect 10643 8993 10655 9027
rect 10597 8987 10655 8993
rect 10778 8984 10784 9036
rect 10836 9024 10842 9036
rect 11790 9024 11796 9036
rect 10836 8996 11796 9024
rect 10836 8984 10842 8996
rect 11790 8984 11796 8996
rect 11848 9024 11854 9036
rect 12820 9024 12848 9055
rect 11848 8996 12664 9024
rect 12820 8996 13492 9024
rect 11848 8984 11854 8996
rect 10229 8959 10287 8965
rect 10229 8956 10241 8959
rect 8312 8928 10241 8956
rect 10229 8925 10241 8928
rect 10275 8925 10287 8959
rect 10229 8919 10287 8925
rect 12158 8916 12164 8968
rect 12216 8956 12222 8968
rect 12253 8959 12311 8965
rect 12253 8956 12265 8959
rect 12216 8928 12265 8956
rect 12216 8916 12222 8928
rect 12253 8925 12265 8928
rect 12299 8925 12311 8959
rect 12253 8919 12311 8925
rect 12342 8916 12348 8968
rect 12400 8956 12406 8968
rect 12526 8956 12532 8968
rect 12400 8928 12532 8956
rect 12400 8916 12406 8928
rect 12526 8916 12532 8928
rect 12584 8916 12590 8968
rect 12636 8965 12664 8996
rect 13464 8965 13492 8996
rect 14274 8984 14280 9036
rect 14332 9024 14338 9036
rect 15013 9027 15071 9033
rect 15013 9024 15025 9027
rect 14332 8996 15025 9024
rect 14332 8984 14338 8996
rect 15013 8993 15025 8996
rect 15059 9024 15071 9027
rect 17494 9024 17500 9036
rect 15059 8996 16712 9024
rect 15059 8993 15071 8996
rect 15013 8987 15071 8993
rect 16684 8968 16712 8996
rect 16960 8996 17500 9024
rect 12621 8959 12679 8965
rect 12621 8925 12633 8959
rect 12667 8956 12679 8959
rect 13173 8959 13231 8965
rect 13173 8956 13185 8959
rect 12667 8928 13185 8956
rect 12667 8925 12679 8928
rect 12621 8919 12679 8925
rect 13173 8925 13185 8928
rect 13219 8925 13231 8959
rect 13173 8919 13231 8925
rect 13265 8959 13323 8965
rect 13265 8925 13277 8959
rect 13311 8925 13323 8959
rect 13265 8919 13323 8925
rect 13449 8959 13507 8965
rect 13449 8925 13461 8959
rect 13495 8925 13507 8959
rect 13449 8919 13507 8925
rect 15381 8959 15439 8965
rect 15381 8925 15393 8959
rect 15427 8956 15439 8959
rect 15470 8956 15476 8968
rect 15427 8928 15476 8956
rect 15427 8925 15439 8928
rect 15381 8919 15439 8925
rect 4856 8860 5488 8888
rect 4856 8848 4862 8860
rect 5902 8848 5908 8900
rect 5960 8888 5966 8900
rect 6730 8888 6736 8900
rect 5960 8860 6736 8888
rect 5960 8848 5966 8860
rect 6730 8848 6736 8860
rect 6788 8848 6794 8900
rect 7282 8848 7288 8900
rect 7340 8848 7346 8900
rect 7926 8848 7932 8900
rect 7984 8888 7990 8900
rect 8021 8891 8079 8897
rect 8021 8888 8033 8891
rect 7984 8860 8033 8888
rect 7984 8848 7990 8860
rect 8021 8857 8033 8860
rect 8067 8857 8079 8891
rect 8021 8851 8079 8857
rect 8846 8848 8852 8900
rect 8904 8888 8910 8900
rect 8904 8860 9352 8888
rect 8904 8848 8910 8860
rect 4816 8820 4844 8848
rect 4172 8792 4844 8820
rect 5813 8823 5871 8829
rect 5813 8789 5825 8823
rect 5859 8820 5871 8823
rect 6105 8823 6163 8829
rect 6105 8820 6117 8823
rect 5859 8792 6117 8820
rect 5859 8789 5871 8792
rect 5813 8783 5871 8789
rect 6105 8789 6117 8792
rect 6151 8789 6163 8823
rect 6105 8783 6163 8789
rect 7374 8780 7380 8832
rect 7432 8820 7438 8832
rect 9324 8829 9352 8860
rect 10962 8848 10968 8900
rect 11020 8848 11026 8900
rect 12437 8891 12495 8897
rect 12437 8857 12449 8891
rect 12483 8857 12495 8891
rect 12437 8851 12495 8857
rect 8941 8823 8999 8829
rect 8941 8820 8953 8823
rect 7432 8792 8953 8820
rect 7432 8780 7438 8792
rect 8941 8789 8953 8792
rect 8987 8789 8999 8823
rect 8941 8783 8999 8789
rect 9309 8823 9367 8829
rect 9309 8789 9321 8823
rect 9355 8820 9367 8823
rect 11882 8820 11888 8832
rect 9355 8792 11888 8820
rect 9355 8789 9367 8792
rect 9309 8783 9367 8789
rect 11882 8780 11888 8792
rect 11940 8820 11946 8832
rect 12452 8820 12480 8851
rect 12894 8848 12900 8900
rect 12952 8848 12958 8900
rect 13081 8891 13139 8897
rect 13081 8857 13093 8891
rect 13127 8857 13139 8891
rect 13280 8888 13308 8919
rect 15470 8916 15476 8928
rect 15528 8916 15534 8968
rect 16666 8916 16672 8968
rect 16724 8956 16730 8968
rect 16960 8965 16988 8996
rect 17494 8984 17500 8996
rect 17552 8984 17558 9036
rect 19352 9033 19380 9132
rect 20622 9120 20628 9172
rect 20680 9160 20686 9172
rect 20717 9163 20775 9169
rect 20717 9160 20729 9163
rect 20680 9132 20729 9160
rect 20680 9120 20686 9132
rect 20717 9129 20729 9132
rect 20763 9129 20775 9163
rect 20717 9123 20775 9129
rect 19797 9095 19855 9101
rect 19797 9061 19809 9095
rect 19843 9092 19855 9095
rect 19843 9064 20668 9092
rect 19843 9061 19855 9064
rect 19797 9055 19855 9061
rect 20640 9036 20668 9064
rect 19337 9027 19395 9033
rect 19337 8993 19349 9027
rect 19383 8993 19395 9027
rect 19337 8987 19395 8993
rect 19886 8984 19892 9036
rect 19944 8984 19950 9036
rect 20622 8984 20628 9036
rect 20680 8984 20686 9036
rect 20732 9024 20760 9123
rect 21361 9095 21419 9101
rect 21361 9061 21373 9095
rect 21407 9092 21419 9095
rect 22462 9092 22468 9104
rect 21407 9064 22468 9092
rect 21407 9061 21419 9064
rect 21361 9055 21419 9061
rect 22462 9052 22468 9064
rect 22520 9052 22526 9104
rect 21085 9027 21143 9033
rect 20732 8996 20944 9024
rect 16945 8959 17003 8965
rect 16945 8956 16957 8959
rect 16724 8928 16957 8956
rect 16724 8916 16730 8928
rect 16945 8925 16957 8928
rect 16991 8925 17003 8959
rect 16945 8919 17003 8925
rect 17034 8916 17040 8968
rect 17092 8956 17098 8968
rect 17313 8959 17371 8965
rect 17313 8956 17325 8959
rect 17092 8928 17325 8956
rect 17092 8916 17098 8928
rect 17313 8925 17325 8928
rect 17359 8925 17371 8959
rect 18782 8956 18788 8968
rect 17313 8919 17371 8925
rect 18340 8928 18788 8956
rect 13081 8851 13139 8857
rect 13188 8860 13308 8888
rect 13096 8820 13124 8851
rect 13188 8832 13216 8860
rect 16390 8848 16396 8900
rect 16448 8848 16454 8900
rect 18340 8874 18368 8928
rect 18782 8916 18788 8928
rect 18840 8916 18846 8968
rect 19058 8916 19064 8968
rect 19116 8956 19122 8968
rect 19429 8959 19487 8965
rect 19429 8956 19441 8959
rect 19116 8928 19441 8956
rect 19116 8916 19122 8928
rect 19429 8925 19441 8928
rect 19475 8925 19487 8959
rect 19429 8919 19487 8925
rect 20070 8916 20076 8968
rect 20128 8916 20134 8968
rect 20533 8959 20591 8965
rect 20533 8925 20545 8959
rect 20579 8956 20591 8959
rect 20714 8956 20720 8968
rect 20579 8928 20720 8956
rect 20579 8925 20591 8928
rect 20533 8919 20591 8925
rect 20714 8916 20720 8928
rect 20772 8916 20778 8968
rect 20349 8891 20407 8897
rect 20349 8888 20361 8891
rect 19260 8860 20361 8888
rect 11940 8792 13124 8820
rect 11940 8780 11946 8792
rect 13170 8780 13176 8832
rect 13228 8780 13234 8832
rect 13633 8823 13691 8829
rect 13633 8789 13645 8823
rect 13679 8820 13691 8823
rect 16758 8820 16764 8832
rect 13679 8792 16764 8820
rect 13679 8789 13691 8792
rect 13633 8783 13691 8789
rect 16758 8780 16764 8792
rect 16816 8780 16822 8832
rect 17402 8780 17408 8832
rect 17460 8820 17466 8832
rect 18739 8823 18797 8829
rect 18739 8820 18751 8823
rect 17460 8792 18751 8820
rect 17460 8780 17466 8792
rect 18739 8789 18751 8792
rect 18785 8820 18797 8823
rect 19260 8820 19288 8860
rect 20349 8857 20361 8860
rect 20395 8888 20407 8891
rect 20438 8888 20444 8900
rect 20395 8860 20444 8888
rect 20395 8857 20407 8860
rect 20349 8851 20407 8857
rect 20438 8848 20444 8860
rect 20496 8848 20502 8900
rect 20916 8888 20944 8996
rect 21085 8993 21097 9027
rect 21131 9024 21143 9027
rect 21821 9027 21879 9033
rect 21821 9024 21833 9027
rect 21131 8996 21833 9024
rect 21131 8993 21143 8996
rect 21085 8987 21143 8993
rect 21821 8993 21833 8996
rect 21867 8993 21879 9027
rect 21821 8987 21879 8993
rect 20990 8916 20996 8968
rect 21048 8916 21054 8968
rect 21450 8916 21456 8968
rect 21508 8916 21514 8968
rect 21546 8959 21604 8965
rect 21546 8925 21558 8959
rect 21592 8925 21604 8959
rect 21546 8919 21604 8925
rect 21560 8888 21588 8919
rect 20916 8860 21588 8888
rect 18785 8792 19288 8820
rect 20257 8823 20315 8829
rect 18785 8789 18797 8792
rect 18739 8783 18797 8789
rect 20257 8789 20269 8823
rect 20303 8820 20315 8823
rect 21174 8820 21180 8832
rect 20303 8792 21180 8820
rect 20303 8789 20315 8792
rect 20257 8783 20315 8789
rect 21174 8780 21180 8792
rect 21232 8780 21238 8832
rect 1104 8730 25208 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 25208 8730
rect 1104 8656 25208 8678
rect 3234 8576 3240 8628
rect 3292 8616 3298 8628
rect 3421 8619 3479 8625
rect 3421 8616 3433 8619
rect 3292 8588 3433 8616
rect 3292 8576 3298 8588
rect 3421 8585 3433 8588
rect 3467 8585 3479 8619
rect 4062 8616 4068 8628
rect 3421 8579 3479 8585
rect 3528 8588 4068 8616
rect 2958 8548 2964 8560
rect 2792 8520 2964 8548
rect 2498 8440 2504 8492
rect 2556 8440 2562 8492
rect 2792 8489 2820 8520
rect 2958 8508 2964 8520
rect 3016 8548 3022 8560
rect 3528 8548 3556 8588
rect 4062 8576 4068 8588
rect 4120 8576 4126 8628
rect 4154 8576 4160 8628
rect 4212 8616 4218 8628
rect 4433 8619 4491 8625
rect 4212 8588 4384 8616
rect 4212 8576 4218 8588
rect 3016 8520 3556 8548
rect 3881 8551 3939 8557
rect 3016 8508 3022 8520
rect 3881 8517 3893 8551
rect 3927 8548 3939 8551
rect 4356 8548 4384 8588
rect 4433 8585 4445 8619
rect 4479 8616 4491 8619
rect 4798 8616 4804 8628
rect 4479 8588 4804 8616
rect 4479 8585 4491 8588
rect 4433 8579 4491 8585
rect 4798 8576 4804 8588
rect 4856 8576 4862 8628
rect 5258 8576 5264 8628
rect 5316 8576 5322 8628
rect 8018 8576 8024 8628
rect 8076 8616 8082 8628
rect 12713 8619 12771 8625
rect 8076 8588 8984 8616
rect 8076 8576 8082 8588
rect 3927 8520 4200 8548
rect 4356 8520 7144 8548
rect 3927 8517 3939 8520
rect 3881 8511 3939 8517
rect 4172 8492 4200 8520
rect 2777 8483 2835 8489
rect 2777 8449 2789 8483
rect 2823 8449 2835 8483
rect 2777 8443 2835 8449
rect 2866 8440 2872 8492
rect 2924 8440 2930 8492
rect 3050 8440 3056 8492
rect 3108 8440 3114 8492
rect 3142 8440 3148 8492
rect 3200 8440 3206 8492
rect 3234 8440 3240 8492
rect 3292 8440 3298 8492
rect 3697 8483 3755 8489
rect 3697 8449 3709 8483
rect 3743 8449 3755 8483
rect 3697 8443 3755 8449
rect 3793 8483 3851 8489
rect 3793 8449 3805 8483
rect 3839 8480 3851 8483
rect 3970 8480 3976 8492
rect 3839 8452 3976 8480
rect 3839 8449 3851 8452
rect 3793 8443 3851 8449
rect 3712 8412 3740 8443
rect 3970 8440 3976 8452
rect 4028 8440 4034 8492
rect 4065 8483 4123 8489
rect 4065 8449 4077 8483
rect 4111 8449 4123 8483
rect 4065 8443 4123 8449
rect 4080 8412 4108 8443
rect 4154 8440 4160 8492
rect 4212 8440 4218 8492
rect 4338 8440 4344 8492
rect 4396 8440 4402 8492
rect 4798 8480 4804 8492
rect 4448 8452 4804 8480
rect 4448 8412 4476 8452
rect 4798 8440 4804 8452
rect 4856 8440 4862 8492
rect 5166 8440 5172 8492
rect 5224 8440 5230 8492
rect 5258 8440 5264 8492
rect 5316 8480 5322 8492
rect 5353 8483 5411 8489
rect 5353 8480 5365 8483
rect 5316 8452 5365 8480
rect 5316 8440 5322 8452
rect 5353 8449 5365 8452
rect 5399 8480 5411 8483
rect 5534 8480 5540 8492
rect 5399 8452 5540 8480
rect 5399 8449 5411 8452
rect 5353 8443 5411 8449
rect 5534 8440 5540 8452
rect 5592 8440 5598 8492
rect 5629 8483 5687 8489
rect 5629 8449 5641 8483
rect 5675 8480 5687 8483
rect 5718 8480 5724 8492
rect 5675 8452 5724 8480
rect 5675 8449 5687 8452
rect 5629 8443 5687 8449
rect 5718 8440 5724 8452
rect 5776 8440 5782 8492
rect 6914 8440 6920 8492
rect 6972 8480 6978 8492
rect 7009 8483 7067 8489
rect 7009 8480 7021 8483
rect 6972 8452 7021 8480
rect 6972 8440 6978 8452
rect 7009 8449 7021 8452
rect 7055 8449 7067 8483
rect 7116 8480 7144 8520
rect 8202 8508 8208 8560
rect 8260 8508 8266 8560
rect 8846 8508 8852 8560
rect 8904 8508 8910 8560
rect 7282 8480 7288 8492
rect 7116 8452 7288 8480
rect 7009 8443 7067 8449
rect 7282 8440 7288 8452
rect 7340 8440 7346 8492
rect 7374 8440 7380 8492
rect 7432 8440 7438 8492
rect 2700 8384 2820 8412
rect 3712 8384 4016 8412
rect 4080 8384 4476 8412
rect 2222 8304 2228 8356
rect 2280 8304 2286 8356
rect 2593 8279 2651 8285
rect 2593 8245 2605 8279
rect 2639 8276 2651 8279
rect 2700 8276 2728 8384
rect 2792 8344 2820 8384
rect 3234 8344 3240 8356
rect 2792 8316 3240 8344
rect 3234 8304 3240 8316
rect 3292 8344 3298 8356
rect 3513 8347 3571 8353
rect 3513 8344 3525 8347
rect 3292 8316 3525 8344
rect 3292 8304 3298 8316
rect 3513 8313 3525 8316
rect 3559 8313 3571 8347
rect 3513 8307 3571 8313
rect 3988 8288 4016 8384
rect 4706 8372 4712 8424
rect 4764 8372 4770 8424
rect 8220 8412 8248 8508
rect 8956 8489 8984 8588
rect 12713 8585 12725 8619
rect 12759 8616 12771 8619
rect 12894 8616 12900 8628
rect 12759 8588 12900 8616
rect 12759 8585 12771 8588
rect 12713 8579 12771 8585
rect 12894 8576 12900 8588
rect 12952 8576 12958 8628
rect 17034 8576 17040 8628
rect 17092 8576 17098 8628
rect 17402 8576 17408 8628
rect 17460 8576 17466 8628
rect 20254 8576 20260 8628
rect 20312 8616 20318 8628
rect 21450 8616 21456 8628
rect 20312 8588 21456 8616
rect 20312 8576 20318 8588
rect 21450 8576 21456 8588
rect 21508 8576 21514 8628
rect 8941 8483 8999 8489
rect 8941 8449 8953 8483
rect 8987 8449 8999 8483
rect 8941 8443 8999 8449
rect 9306 8440 9312 8492
rect 9364 8440 9370 8492
rect 10060 8412 10088 8534
rect 16022 8508 16028 8560
rect 16080 8548 16086 8560
rect 17497 8551 17555 8557
rect 17497 8548 17509 8551
rect 16080 8520 17509 8548
rect 16080 8508 16086 8520
rect 17497 8517 17509 8520
rect 17543 8517 17555 8551
rect 17497 8511 17555 8517
rect 10134 8440 10140 8492
rect 10192 8480 10198 8492
rect 10778 8480 10784 8492
rect 10192 8452 10784 8480
rect 10192 8440 10198 8452
rect 10778 8440 10784 8452
rect 10836 8440 10842 8492
rect 12526 8440 12532 8492
rect 12584 8480 12590 8492
rect 12802 8480 12808 8492
rect 12584 8452 12808 8480
rect 12584 8440 12590 8452
rect 12802 8440 12808 8452
rect 12860 8440 12866 8492
rect 13354 8440 13360 8492
rect 13412 8480 13418 8492
rect 13449 8483 13507 8489
rect 13449 8480 13461 8483
rect 13412 8452 13461 8480
rect 13412 8440 13418 8452
rect 13449 8449 13461 8452
rect 13495 8480 13507 8483
rect 17218 8480 17224 8492
rect 13495 8452 17224 8480
rect 13495 8449 13507 8452
rect 13449 8443 13507 8449
rect 17218 8440 17224 8452
rect 17276 8440 17282 8492
rect 20438 8440 20444 8492
rect 20496 8440 20502 8492
rect 20625 8483 20683 8489
rect 20625 8449 20637 8483
rect 20671 8480 20683 8483
rect 20714 8480 20720 8492
rect 20671 8452 20720 8480
rect 20671 8449 20683 8452
rect 20625 8443 20683 8449
rect 20714 8440 20720 8452
rect 20772 8440 20778 8492
rect 10226 8412 10232 8424
rect 8220 8384 10232 8412
rect 10226 8372 10232 8384
rect 10284 8372 10290 8424
rect 12158 8372 12164 8424
rect 12216 8412 12222 8424
rect 12345 8415 12403 8421
rect 12345 8412 12357 8415
rect 12216 8384 12357 8412
rect 12216 8372 12222 8384
rect 12345 8381 12357 8384
rect 12391 8381 12403 8415
rect 12345 8375 12403 8381
rect 15930 8372 15936 8424
rect 15988 8412 15994 8424
rect 17589 8415 17647 8421
rect 17589 8412 17601 8415
rect 15988 8384 17601 8412
rect 15988 8372 15994 8384
rect 17589 8381 17601 8384
rect 17635 8412 17647 8415
rect 18598 8412 18604 8424
rect 17635 8384 18604 8412
rect 17635 8381 17647 8384
rect 17589 8375 17647 8381
rect 18598 8372 18604 8384
rect 18656 8372 18662 8424
rect 4890 8344 4896 8356
rect 4816 8316 4896 8344
rect 2639 8248 2728 8276
rect 2639 8245 2651 8248
rect 2593 8239 2651 8245
rect 3970 8236 3976 8288
rect 4028 8276 4034 8288
rect 4816 8285 4844 8316
rect 4890 8304 4896 8316
rect 4948 8344 4954 8356
rect 6362 8344 6368 8356
rect 4948 8316 6368 8344
rect 4948 8304 4954 8316
rect 6362 8304 6368 8316
rect 6420 8304 6426 8356
rect 4249 8279 4307 8285
rect 4249 8276 4261 8279
rect 4028 8248 4261 8276
rect 4028 8236 4034 8248
rect 4249 8245 4261 8248
rect 4295 8245 4307 8279
rect 4249 8239 4307 8245
rect 4801 8279 4859 8285
rect 4801 8245 4813 8279
rect 4847 8245 4859 8279
rect 4801 8239 4859 8245
rect 5166 8236 5172 8288
rect 5224 8276 5230 8288
rect 5626 8276 5632 8288
rect 5224 8248 5632 8276
rect 5224 8236 5230 8248
rect 5626 8236 5632 8248
rect 5684 8276 5690 8288
rect 5721 8279 5779 8285
rect 5721 8276 5733 8279
rect 5684 8248 5733 8276
rect 5684 8236 5690 8248
rect 5721 8245 5733 8248
rect 5767 8276 5779 8279
rect 7190 8276 7196 8288
rect 5767 8248 7196 8276
rect 5767 8245 5779 8248
rect 5721 8239 5779 8245
rect 7190 8236 7196 8248
rect 7248 8236 7254 8288
rect 12986 8236 12992 8288
rect 13044 8276 13050 8288
rect 13630 8276 13636 8288
rect 13044 8248 13636 8276
rect 13044 8236 13050 8248
rect 13630 8236 13636 8248
rect 13688 8236 13694 8288
rect 1104 8186 25208 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 25208 8186
rect 1104 8112 25208 8134
rect 2685 8075 2743 8081
rect 2685 8041 2697 8075
rect 2731 8041 2743 8075
rect 2685 8035 2743 8041
rect 2869 8075 2927 8081
rect 2869 8041 2881 8075
rect 2915 8072 2927 8075
rect 3050 8072 3056 8084
rect 2915 8044 3056 8072
rect 2915 8041 2927 8044
rect 2869 8035 2927 8041
rect 2700 7936 2728 8035
rect 3050 8032 3056 8044
rect 3108 8032 3114 8084
rect 3326 8032 3332 8084
rect 3384 8032 3390 8084
rect 3602 8032 3608 8084
rect 3660 8032 3666 8084
rect 12250 8032 12256 8084
rect 12308 8072 12314 8084
rect 12345 8075 12403 8081
rect 12345 8072 12357 8075
rect 12308 8044 12357 8072
rect 12308 8032 12314 8044
rect 12345 8041 12357 8044
rect 12391 8041 12403 8075
rect 12345 8035 12403 8041
rect 16071 8075 16129 8081
rect 16071 8041 16083 8075
rect 16117 8072 16129 8075
rect 16574 8072 16580 8084
rect 16117 8044 16580 8072
rect 16117 8041 16129 8044
rect 16071 8035 16129 8041
rect 16574 8032 16580 8044
rect 16632 8072 16638 8084
rect 17770 8072 17776 8084
rect 16632 8044 17776 8072
rect 16632 8032 16638 8044
rect 17770 8032 17776 8044
rect 17828 8032 17834 8084
rect 2958 7964 2964 8016
rect 3016 7964 3022 8016
rect 5258 8004 5264 8016
rect 3160 7976 5264 8004
rect 3160 7948 3188 7976
rect 5258 7964 5264 7976
rect 5316 7964 5322 8016
rect 6362 7964 6368 8016
rect 6420 8004 6426 8016
rect 6457 8007 6515 8013
rect 6457 8004 6469 8007
rect 6420 7976 6469 8004
rect 6420 7964 6426 7976
rect 6457 7973 6469 7976
rect 6503 8004 6515 8007
rect 6914 8004 6920 8016
rect 6503 7976 6920 8004
rect 6503 7973 6515 7976
rect 6457 7967 6515 7973
rect 6914 7964 6920 7976
rect 6972 7964 6978 8016
rect 12713 8007 12771 8013
rect 12713 7973 12725 8007
rect 12759 8004 12771 8007
rect 12759 7976 13216 8004
rect 12759 7973 12771 7976
rect 12713 7967 12771 7973
rect 3142 7936 3148 7948
rect 2700 7908 3148 7936
rect 3142 7896 3148 7908
rect 3200 7896 3206 7948
rect 3234 7896 3240 7948
rect 3292 7896 3298 7948
rect 3694 7896 3700 7948
rect 3752 7936 3758 7948
rect 4890 7936 4896 7948
rect 3752 7908 4108 7936
rect 3752 7896 3758 7908
rect 3329 7871 3387 7877
rect 3329 7837 3341 7871
rect 3375 7837 3387 7871
rect 3329 7831 3387 7837
rect 2501 7803 2559 7809
rect 2501 7769 2513 7803
rect 2547 7800 2559 7803
rect 3344 7800 3372 7831
rect 3418 7828 3424 7880
rect 3476 7828 3482 7880
rect 3605 7871 3663 7877
rect 3605 7837 3617 7871
rect 3651 7868 3663 7871
rect 3651 7840 3924 7868
rect 3651 7837 3663 7840
rect 3605 7831 3663 7837
rect 3896 7812 3924 7840
rect 3970 7828 3976 7880
rect 4028 7828 4034 7880
rect 4080 7877 4108 7908
rect 4172 7908 4896 7936
rect 4065 7871 4123 7877
rect 4065 7837 4077 7871
rect 4111 7837 4123 7871
rect 4065 7831 4123 7837
rect 3789 7803 3847 7809
rect 3789 7800 3801 7803
rect 2547 7772 3280 7800
rect 3344 7772 3801 7800
rect 2547 7769 2559 7772
rect 2501 7763 2559 7769
rect 2711 7735 2769 7741
rect 2711 7701 2723 7735
rect 2757 7732 2769 7735
rect 2866 7732 2872 7744
rect 2757 7704 2872 7732
rect 2757 7701 2769 7704
rect 2711 7695 2769 7701
rect 2866 7692 2872 7704
rect 2924 7692 2930 7744
rect 3252 7732 3280 7772
rect 3789 7769 3801 7772
rect 3835 7769 3847 7803
rect 3789 7763 3847 7769
rect 3878 7760 3884 7812
rect 3936 7800 3942 7812
rect 4172 7800 4200 7908
rect 4890 7896 4896 7908
rect 4948 7896 4954 7948
rect 5718 7896 5724 7948
rect 5776 7936 5782 7948
rect 5997 7939 6055 7945
rect 5997 7936 6009 7939
rect 5776 7908 6009 7936
rect 5776 7896 5782 7908
rect 5997 7905 6009 7908
rect 6043 7905 6055 7939
rect 7469 7939 7527 7945
rect 7469 7936 7481 7939
rect 5997 7899 6055 7905
rect 6656 7908 7481 7936
rect 4249 7871 4307 7877
rect 4249 7837 4261 7871
rect 4295 7837 4307 7871
rect 4249 7831 4307 7837
rect 3936 7772 4200 7800
rect 4264 7800 4292 7831
rect 4338 7828 4344 7880
rect 4396 7828 4402 7880
rect 5442 7828 5448 7880
rect 5500 7828 5506 7880
rect 6012 7868 6040 7899
rect 6656 7877 6684 7908
rect 7469 7905 7481 7908
rect 7515 7905 7527 7939
rect 7469 7899 7527 7905
rect 12986 7896 12992 7948
rect 13044 7896 13050 7948
rect 13188 7945 13216 7976
rect 13814 7964 13820 8016
rect 13872 7964 13878 8016
rect 13173 7939 13231 7945
rect 13173 7905 13185 7939
rect 13219 7936 13231 7939
rect 13219 7908 13676 7936
rect 13219 7905 13231 7908
rect 13173 7899 13231 7905
rect 6365 7871 6423 7877
rect 6365 7868 6377 7871
rect 6012 7840 6377 7868
rect 6365 7837 6377 7840
rect 6411 7837 6423 7871
rect 6365 7831 6423 7837
rect 6549 7871 6607 7877
rect 6549 7837 6561 7871
rect 6595 7837 6607 7871
rect 6549 7831 6607 7837
rect 6641 7871 6699 7877
rect 6641 7837 6653 7871
rect 6687 7837 6699 7871
rect 6641 7831 6699 7837
rect 4706 7800 4712 7812
rect 4264 7772 4712 7800
rect 3936 7760 3942 7772
rect 4706 7760 4712 7772
rect 4764 7760 4770 7812
rect 5460 7800 5488 7828
rect 6564 7800 6592 7831
rect 6730 7828 6736 7880
rect 6788 7868 6794 7880
rect 6825 7871 6883 7877
rect 6825 7868 6837 7871
rect 6788 7840 6837 7868
rect 6788 7828 6794 7840
rect 6825 7837 6837 7840
rect 6871 7837 6883 7871
rect 6825 7831 6883 7837
rect 6914 7828 6920 7880
rect 6972 7828 6978 7880
rect 7101 7871 7159 7877
rect 7101 7837 7113 7871
rect 7147 7868 7159 7871
rect 7190 7868 7196 7880
rect 7147 7840 7196 7868
rect 7147 7837 7159 7840
rect 7101 7831 7159 7837
rect 7190 7828 7196 7840
rect 7248 7828 7254 7880
rect 7282 7828 7288 7880
rect 7340 7868 7346 7880
rect 7561 7871 7619 7877
rect 7561 7868 7573 7871
rect 7340 7840 7573 7868
rect 7340 7828 7346 7840
rect 7561 7837 7573 7840
rect 7607 7868 7619 7871
rect 9674 7868 9680 7880
rect 7607 7840 9680 7868
rect 7607 7837 7619 7840
rect 7561 7831 7619 7837
rect 9674 7828 9680 7840
rect 9732 7828 9738 7880
rect 12342 7828 12348 7880
rect 12400 7828 12406 7880
rect 12434 7828 12440 7880
rect 12492 7828 12498 7880
rect 13081 7871 13139 7877
rect 13081 7837 13093 7871
rect 13127 7837 13139 7871
rect 13081 7831 13139 7837
rect 5184 7772 6592 7800
rect 13096 7800 13124 7831
rect 13262 7828 13268 7880
rect 13320 7868 13326 7880
rect 13648 7877 13676 7908
rect 14274 7896 14280 7948
rect 14332 7896 14338 7948
rect 13541 7871 13599 7877
rect 13541 7868 13553 7871
rect 13320 7840 13553 7868
rect 13320 7828 13326 7840
rect 13541 7837 13553 7840
rect 13587 7837 13599 7871
rect 13541 7831 13599 7837
rect 13633 7871 13691 7877
rect 13633 7837 13645 7871
rect 13679 7837 13691 7871
rect 13633 7831 13691 7837
rect 14642 7828 14648 7880
rect 14700 7828 14706 7880
rect 18506 7828 18512 7880
rect 18564 7828 18570 7880
rect 13170 7800 13176 7812
rect 13096 7772 13176 7800
rect 3896 7732 3924 7760
rect 3252 7704 3924 7732
rect 4246 7692 4252 7744
rect 4304 7732 4310 7744
rect 5184 7732 5212 7772
rect 13170 7760 13176 7772
rect 13228 7800 13234 7812
rect 13817 7803 13875 7809
rect 13817 7800 13829 7803
rect 13228 7772 13829 7800
rect 13228 7760 13234 7772
rect 13817 7769 13829 7772
rect 13863 7769 13875 7803
rect 16390 7800 16396 7812
rect 15686 7772 16396 7800
rect 13817 7763 13875 7769
rect 16390 7760 16396 7772
rect 16448 7760 16454 7812
rect 4304 7704 5212 7732
rect 4304 7692 4310 7704
rect 5442 7692 5448 7744
rect 5500 7692 5506 7744
rect 5902 7692 5908 7744
rect 5960 7732 5966 7744
rect 6181 7735 6239 7741
rect 6181 7732 6193 7735
rect 5960 7704 6193 7732
rect 5960 7692 5966 7704
rect 6181 7701 6193 7704
rect 6227 7701 6239 7735
rect 6181 7695 6239 7701
rect 6730 7692 6736 7744
rect 6788 7732 6794 7744
rect 7285 7735 7343 7741
rect 7285 7732 7297 7735
rect 6788 7704 7297 7732
rect 6788 7692 6794 7704
rect 7285 7701 7297 7704
rect 7331 7701 7343 7735
rect 7285 7695 7343 7701
rect 7374 7692 7380 7744
rect 7432 7732 7438 7744
rect 13354 7732 13360 7744
rect 7432 7704 13360 7732
rect 7432 7692 7438 7704
rect 13354 7692 13360 7704
rect 13412 7692 13418 7744
rect 13446 7692 13452 7744
rect 13504 7692 13510 7744
rect 18782 7692 18788 7744
rect 18840 7692 18846 7744
rect 1104 7642 25208 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 25208 7642
rect 1104 7568 25208 7590
rect 2866 7488 2872 7540
rect 2924 7528 2930 7540
rect 4062 7528 4068 7540
rect 2924 7500 4068 7528
rect 2924 7488 2930 7500
rect 4062 7488 4068 7500
rect 4120 7488 4126 7540
rect 4154 7488 4160 7540
rect 4212 7528 4218 7540
rect 4338 7528 4344 7540
rect 4212 7500 4344 7528
rect 4212 7488 4218 7500
rect 4338 7488 4344 7500
rect 4396 7488 4402 7540
rect 4893 7531 4951 7537
rect 4893 7497 4905 7531
rect 4939 7528 4951 7531
rect 5258 7528 5264 7540
rect 4939 7500 5264 7528
rect 4939 7497 4951 7500
rect 4893 7491 4951 7497
rect 5258 7488 5264 7500
rect 5316 7488 5322 7540
rect 5350 7488 5356 7540
rect 5408 7488 5414 7540
rect 6917 7531 6975 7537
rect 6917 7497 6929 7531
rect 6963 7528 6975 7531
rect 7374 7528 7380 7540
rect 6963 7500 7380 7528
rect 6963 7497 6975 7500
rect 6917 7491 6975 7497
rect 7374 7488 7380 7500
rect 7432 7488 7438 7540
rect 9033 7531 9091 7537
rect 9033 7497 9045 7531
rect 9079 7528 9091 7531
rect 9398 7528 9404 7540
rect 9079 7500 9404 7528
rect 9079 7497 9091 7500
rect 9033 7491 9091 7497
rect 9398 7488 9404 7500
rect 9456 7488 9462 7540
rect 10229 7531 10287 7537
rect 10229 7497 10241 7531
rect 10275 7528 10287 7531
rect 10318 7528 10324 7540
rect 10275 7500 10324 7528
rect 10275 7497 10287 7500
rect 10229 7491 10287 7497
rect 10318 7488 10324 7500
rect 10376 7488 10382 7540
rect 11977 7531 12035 7537
rect 11977 7497 11989 7531
rect 12023 7528 12035 7531
rect 13262 7528 13268 7540
rect 12023 7500 13268 7528
rect 12023 7497 12035 7500
rect 11977 7491 12035 7497
rect 13262 7488 13268 7500
rect 13320 7488 13326 7540
rect 14277 7531 14335 7537
rect 14277 7497 14289 7531
rect 14323 7528 14335 7531
rect 14642 7528 14648 7540
rect 14323 7500 14648 7528
rect 14323 7497 14335 7500
rect 14277 7491 14335 7497
rect 14642 7488 14648 7500
rect 14700 7488 14706 7540
rect 19610 7528 19616 7540
rect 17972 7500 19616 7528
rect 3602 7420 3608 7472
rect 3660 7460 3666 7472
rect 5077 7463 5135 7469
rect 5077 7460 5089 7463
rect 3660 7432 4568 7460
rect 3660 7420 3666 7432
rect 3142 7392 3148 7404
rect 3103 7364 3148 7392
rect 3142 7352 3148 7364
rect 3200 7352 3206 7404
rect 3237 7395 3295 7401
rect 3237 7361 3249 7395
rect 3283 7392 3295 7395
rect 3510 7392 3516 7404
rect 3283 7364 3516 7392
rect 3283 7361 3295 7364
rect 3237 7355 3295 7361
rect 3510 7352 3516 7364
rect 3568 7352 3574 7404
rect 3878 7352 3884 7404
rect 3936 7392 3942 7404
rect 4065 7395 4123 7401
rect 4065 7392 4077 7395
rect 3936 7364 4077 7392
rect 3936 7352 3942 7364
rect 4065 7361 4077 7364
rect 4111 7361 4123 7395
rect 4065 7355 4123 7361
rect 4246 7352 4252 7404
rect 4304 7352 4310 7404
rect 4540 7401 4568 7432
rect 4632 7432 5089 7460
rect 4632 7401 4660 7432
rect 5077 7429 5089 7432
rect 5123 7460 5135 7463
rect 5166 7460 5172 7472
rect 5123 7432 5172 7460
rect 5123 7429 5135 7432
rect 5077 7423 5135 7429
rect 5166 7420 5172 7432
rect 5224 7420 5230 7472
rect 5368 7460 5396 7488
rect 5368 7432 5856 7460
rect 4341 7395 4399 7401
rect 4341 7361 4353 7395
rect 4387 7361 4399 7395
rect 4341 7355 4399 7361
rect 4525 7395 4583 7401
rect 4525 7361 4537 7395
rect 4571 7361 4583 7395
rect 4525 7355 4583 7361
rect 4617 7395 4675 7401
rect 4617 7361 4629 7395
rect 4663 7361 4675 7395
rect 4617 7355 4675 7361
rect 4801 7395 4859 7401
rect 4801 7361 4813 7395
rect 4847 7392 4859 7395
rect 5261 7395 5319 7401
rect 5261 7392 5273 7395
rect 4847 7364 5273 7392
rect 4847 7361 4859 7364
rect 4801 7355 4859 7361
rect 5261 7361 5273 7364
rect 5307 7392 5319 7395
rect 5350 7392 5356 7404
rect 5307 7364 5356 7392
rect 5307 7361 5319 7364
rect 5261 7355 5319 7361
rect 4356 7324 4384 7355
rect 5350 7352 5356 7364
rect 5408 7392 5414 7404
rect 5828 7401 5856 7432
rect 6730 7420 6736 7472
rect 6788 7420 6794 7472
rect 11808 7432 12388 7460
rect 5537 7395 5595 7401
rect 5537 7392 5549 7395
rect 5408 7364 5549 7392
rect 5408 7352 5414 7364
rect 5537 7361 5549 7364
rect 5583 7361 5595 7395
rect 5537 7355 5595 7361
rect 5813 7395 5871 7401
rect 5813 7361 5825 7395
rect 5859 7361 5871 7395
rect 5813 7355 5871 7361
rect 4890 7324 4896 7336
rect 4356 7296 4896 7324
rect 4890 7284 4896 7296
rect 4948 7284 4954 7336
rect 4433 7259 4491 7265
rect 4433 7225 4445 7259
rect 4479 7256 4491 7259
rect 4982 7256 4988 7268
rect 4479 7228 4988 7256
rect 4479 7225 4491 7228
rect 4433 7219 4491 7225
rect 4982 7216 4988 7228
rect 5040 7256 5046 7268
rect 5828 7256 5856 7355
rect 5902 7352 5908 7404
rect 5960 7352 5966 7404
rect 6546 7352 6552 7404
rect 6604 7352 6610 7404
rect 6748 7256 6776 7420
rect 8941 7395 8999 7401
rect 8941 7361 8953 7395
rect 8987 7392 8999 7395
rect 9858 7392 9864 7404
rect 8987 7364 9864 7392
rect 8987 7361 8999 7364
rect 8941 7355 8999 7361
rect 9858 7352 9864 7364
rect 9916 7352 9922 7404
rect 10134 7352 10140 7404
rect 10192 7352 10198 7404
rect 10781 7395 10839 7401
rect 10781 7361 10793 7395
rect 10827 7361 10839 7395
rect 10781 7355 10839 7361
rect 9217 7327 9275 7333
rect 9217 7293 9229 7327
rect 9263 7324 9275 7327
rect 9674 7324 9680 7336
rect 9263 7296 9680 7324
rect 9263 7293 9275 7296
rect 9217 7287 9275 7293
rect 9674 7284 9680 7296
rect 9732 7324 9738 7336
rect 10321 7327 10379 7333
rect 10321 7324 10333 7327
rect 9732 7296 10333 7324
rect 9732 7284 9738 7296
rect 10321 7293 10333 7296
rect 10367 7293 10379 7327
rect 10321 7287 10379 7293
rect 5040 7228 5856 7256
rect 5920 7228 6776 7256
rect 10796 7256 10824 7355
rect 11698 7352 11704 7404
rect 11756 7352 11762 7404
rect 11808 7401 11836 7432
rect 12360 7404 12388 7432
rect 13630 7420 13636 7472
rect 13688 7460 13694 7472
rect 14921 7463 14979 7469
rect 13688 7432 14872 7460
rect 13688 7420 13694 7432
rect 11793 7395 11851 7401
rect 11793 7361 11805 7395
rect 11839 7361 11851 7395
rect 11793 7355 11851 7361
rect 12069 7395 12127 7401
rect 12069 7361 12081 7395
rect 12115 7361 12127 7395
rect 12069 7355 12127 7361
rect 11977 7327 12035 7333
rect 11977 7293 11989 7327
rect 12023 7324 12035 7327
rect 12084 7324 12112 7355
rect 12250 7352 12256 7404
rect 12308 7352 12314 7404
rect 12342 7352 12348 7404
rect 12400 7392 12406 7404
rect 12529 7395 12587 7401
rect 12529 7392 12541 7395
rect 12400 7364 12541 7392
rect 12400 7352 12406 7364
rect 12529 7361 12541 7364
rect 12575 7392 12587 7395
rect 12894 7392 12900 7404
rect 12575 7364 12900 7392
rect 12575 7361 12587 7364
rect 12529 7355 12587 7361
rect 12894 7352 12900 7364
rect 12952 7352 12958 7404
rect 13173 7395 13231 7401
rect 13173 7361 13185 7395
rect 13219 7361 13231 7395
rect 13173 7355 13231 7361
rect 12434 7324 12440 7336
rect 12023 7296 12440 7324
rect 12023 7293 12035 7296
rect 11977 7287 12035 7293
rect 12434 7284 12440 7296
rect 12492 7284 12498 7336
rect 12713 7327 12771 7333
rect 12713 7293 12725 7327
rect 12759 7324 12771 7327
rect 13081 7327 13139 7333
rect 13081 7324 13093 7327
rect 12759 7296 13093 7324
rect 12759 7293 12771 7296
rect 12713 7287 12771 7293
rect 13081 7293 13093 7296
rect 13127 7293 13139 7327
rect 13188 7324 13216 7355
rect 13446 7352 13452 7404
rect 13504 7392 13510 7404
rect 14553 7395 14611 7401
rect 14553 7392 14565 7395
rect 13504 7364 14565 7392
rect 13504 7352 13510 7364
rect 14553 7361 14565 7364
rect 14599 7361 14611 7395
rect 14553 7355 14611 7361
rect 13814 7324 13820 7336
rect 13188 7296 13820 7324
rect 13081 7287 13139 7293
rect 13814 7284 13820 7296
rect 13872 7324 13878 7336
rect 14844 7333 14872 7432
rect 14921 7429 14933 7463
rect 14967 7460 14979 7463
rect 16574 7460 16580 7472
rect 14967 7432 16580 7460
rect 14967 7429 14979 7432
rect 14921 7423 14979 7429
rect 16574 7420 16580 7432
rect 16632 7420 16638 7472
rect 17221 7463 17279 7469
rect 17221 7429 17233 7463
rect 17267 7460 17279 7463
rect 17972 7460 18000 7500
rect 19610 7488 19616 7500
rect 19668 7537 19674 7540
rect 19668 7531 19717 7537
rect 19668 7497 19671 7531
rect 19705 7497 19717 7531
rect 19668 7491 19717 7497
rect 19668 7488 19674 7491
rect 17267 7432 18000 7460
rect 17267 7429 17279 7432
rect 17221 7423 17279 7429
rect 18598 7420 18604 7472
rect 18656 7420 18662 7472
rect 16942 7352 16948 7404
rect 17000 7352 17006 7404
rect 17126 7352 17132 7404
rect 17184 7352 17190 7404
rect 17313 7395 17371 7401
rect 17313 7361 17325 7395
rect 17359 7361 17371 7395
rect 18233 7395 18291 7401
rect 18233 7392 18245 7395
rect 17313 7355 17371 7361
rect 17512 7364 18245 7392
rect 14461 7327 14519 7333
rect 14461 7324 14473 7327
rect 13872 7296 14473 7324
rect 13872 7284 13878 7296
rect 14461 7293 14473 7296
rect 14507 7293 14519 7327
rect 14461 7287 14519 7293
rect 14829 7327 14887 7333
rect 14829 7293 14841 7327
rect 14875 7324 14887 7327
rect 17218 7324 17224 7336
rect 14875 7296 17224 7324
rect 14875 7293 14887 7296
rect 14829 7287 14887 7293
rect 17218 7284 17224 7296
rect 17276 7324 17282 7336
rect 17328 7324 17356 7355
rect 17276 7296 17356 7324
rect 17276 7284 17282 7296
rect 13541 7259 13599 7265
rect 10796 7228 11928 7256
rect 5040 7216 5046 7228
rect 3234 7148 3240 7200
rect 3292 7188 3298 7200
rect 4801 7191 4859 7197
rect 4801 7188 4813 7191
rect 3292 7160 4813 7188
rect 3292 7148 3298 7160
rect 4801 7157 4813 7160
rect 4847 7157 4859 7191
rect 4801 7151 4859 7157
rect 5629 7191 5687 7197
rect 5629 7157 5641 7191
rect 5675 7188 5687 7191
rect 5920 7188 5948 7228
rect 5675 7160 5948 7188
rect 5675 7157 5687 7160
rect 5629 7151 5687 7157
rect 5994 7148 6000 7200
rect 6052 7148 6058 7200
rect 8294 7148 8300 7200
rect 8352 7188 8358 7200
rect 8573 7191 8631 7197
rect 8573 7188 8585 7191
rect 8352 7160 8585 7188
rect 8352 7148 8358 7160
rect 8573 7157 8585 7160
rect 8619 7157 8631 7191
rect 8573 7151 8631 7157
rect 9766 7148 9772 7200
rect 9824 7148 9830 7200
rect 10318 7148 10324 7200
rect 10376 7188 10382 7200
rect 10686 7188 10692 7200
rect 10376 7160 10692 7188
rect 10376 7148 10382 7160
rect 10686 7148 10692 7160
rect 10744 7148 10750 7200
rect 11900 7188 11928 7228
rect 13541 7225 13553 7259
rect 13587 7256 13599 7259
rect 13722 7256 13728 7268
rect 13587 7228 13728 7256
rect 13587 7225 13599 7228
rect 13541 7219 13599 7225
rect 13722 7216 13728 7228
rect 13780 7216 13786 7268
rect 17512 7265 17540 7364
rect 18233 7361 18245 7364
rect 18279 7361 18291 7395
rect 18233 7355 18291 7361
rect 17865 7327 17923 7333
rect 17865 7293 17877 7327
rect 17911 7324 17923 7327
rect 18138 7324 18144 7336
rect 17911 7296 18144 7324
rect 17911 7293 17923 7296
rect 17865 7287 17923 7293
rect 18138 7284 18144 7296
rect 18196 7284 18202 7336
rect 17497 7259 17555 7265
rect 17497 7225 17509 7259
rect 17543 7225 17555 7259
rect 21358 7256 21364 7268
rect 17497 7219 17555 7225
rect 19536 7228 21364 7256
rect 19536 7188 19564 7228
rect 21358 7216 21364 7228
rect 21416 7216 21422 7268
rect 11900 7160 19564 7188
rect 1104 7098 25208 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 25208 7098
rect 1104 7024 25208 7046
rect 3602 6944 3608 6996
rect 3660 6944 3666 6996
rect 4617 6987 4675 6993
rect 4617 6953 4629 6987
rect 4663 6984 4675 6987
rect 4706 6984 4712 6996
rect 4663 6956 4712 6984
rect 4663 6953 4675 6956
rect 4617 6947 4675 6953
rect 3053 6919 3111 6925
rect 3053 6885 3065 6919
rect 3099 6916 3111 6919
rect 3878 6916 3884 6928
rect 3099 6888 3884 6916
rect 3099 6885 3111 6888
rect 3053 6879 3111 6885
rect 3878 6876 3884 6888
rect 3936 6876 3942 6928
rect 2130 6808 2136 6860
rect 2188 6848 2194 6860
rect 2498 6848 2504 6860
rect 2188 6820 2504 6848
rect 2188 6808 2194 6820
rect 2498 6808 2504 6820
rect 2556 6808 2562 6860
rect 2961 6851 3019 6857
rect 2961 6817 2973 6851
rect 3007 6848 3019 6851
rect 4632 6848 4660 6947
rect 4706 6944 4712 6956
rect 4764 6944 4770 6996
rect 4890 6944 4896 6996
rect 4948 6944 4954 6996
rect 5074 6944 5080 6996
rect 5132 6984 5138 6996
rect 5537 6987 5595 6993
rect 5537 6984 5549 6987
rect 5132 6956 5549 6984
rect 5132 6944 5138 6956
rect 5537 6953 5549 6956
rect 5583 6953 5595 6987
rect 9582 6984 9588 6996
rect 5537 6947 5595 6953
rect 8772 6956 9588 6984
rect 8772 6916 8800 6956
rect 9582 6944 9588 6956
rect 9640 6944 9646 6996
rect 10134 6944 10140 6996
rect 10192 6984 10198 6996
rect 11054 6993 11060 6996
rect 11011 6987 11060 6993
rect 11011 6984 11023 6987
rect 10192 6956 11023 6984
rect 10192 6944 10198 6956
rect 11011 6953 11023 6956
rect 11057 6953 11060 6987
rect 11011 6947 11060 6953
rect 11054 6944 11060 6947
rect 11112 6984 11118 6996
rect 11606 6984 11612 6996
rect 11112 6956 11612 6984
rect 11112 6944 11118 6956
rect 11606 6944 11612 6956
rect 11664 6944 11670 6996
rect 11698 6944 11704 6996
rect 11756 6984 11762 6996
rect 12069 6987 12127 6993
rect 12069 6984 12081 6987
rect 11756 6956 12081 6984
rect 11756 6944 11762 6956
rect 12069 6953 12081 6956
rect 12115 6984 12127 6987
rect 12250 6984 12256 6996
rect 12115 6956 12256 6984
rect 12115 6953 12127 6956
rect 12069 6947 12127 6953
rect 12250 6944 12256 6956
rect 12308 6944 12314 6996
rect 12526 6944 12532 6996
rect 12584 6984 12590 6996
rect 12713 6987 12771 6993
rect 12713 6984 12725 6987
rect 12584 6956 12725 6984
rect 12584 6944 12590 6956
rect 12713 6953 12725 6956
rect 12759 6953 12771 6987
rect 12713 6947 12771 6953
rect 16393 6987 16451 6993
rect 16393 6953 16405 6987
rect 16439 6984 16451 6987
rect 16942 6984 16948 6996
rect 16439 6956 16948 6984
rect 16439 6953 16451 6956
rect 16393 6947 16451 6953
rect 16942 6944 16948 6956
rect 17000 6944 17006 6996
rect 18598 6944 18604 6996
rect 18656 6984 18662 6996
rect 19978 6984 19984 6996
rect 18656 6956 19984 6984
rect 18656 6944 18662 6956
rect 19978 6944 19984 6956
rect 20036 6944 20042 6996
rect 20714 6944 20720 6996
rect 20772 6984 20778 6996
rect 21039 6987 21097 6993
rect 21039 6984 21051 6987
rect 20772 6956 21051 6984
rect 20772 6944 20778 6956
rect 21039 6953 21051 6956
rect 21085 6953 21097 6987
rect 21039 6947 21097 6953
rect 12158 6916 12164 6928
rect 8680 6888 8800 6916
rect 11532 6888 12164 6916
rect 3007 6820 3464 6848
rect 3007 6817 3019 6820
rect 2961 6811 3019 6817
rect 2222 6740 2228 6792
rect 2280 6780 2286 6792
rect 3436 6789 3464 6820
rect 4080 6820 4660 6848
rect 4709 6851 4767 6857
rect 2317 6783 2375 6789
rect 2317 6780 2329 6783
rect 2280 6752 2329 6780
rect 2280 6740 2286 6752
rect 2317 6749 2329 6752
rect 2363 6749 2375 6783
rect 2317 6743 2375 6749
rect 3237 6783 3295 6789
rect 3237 6749 3249 6783
rect 3283 6749 3295 6783
rect 3237 6743 3295 6749
rect 3421 6783 3479 6789
rect 3421 6749 3433 6783
rect 3467 6780 3479 6783
rect 3510 6780 3516 6792
rect 3467 6752 3516 6780
rect 3467 6749 3479 6752
rect 3421 6743 3479 6749
rect 2409 6715 2467 6721
rect 2409 6681 2421 6715
rect 2455 6712 2467 6715
rect 3142 6712 3148 6724
rect 2455 6684 3148 6712
rect 2455 6681 2467 6684
rect 2409 6675 2467 6681
rect 3142 6672 3148 6684
rect 3200 6712 3206 6724
rect 3252 6712 3280 6743
rect 3510 6740 3516 6752
rect 3568 6740 3574 6792
rect 4080 6789 4108 6820
rect 4709 6817 4721 6851
rect 4755 6848 4767 6851
rect 4890 6848 4896 6860
rect 4755 6820 4896 6848
rect 4755 6817 4767 6820
rect 4709 6811 4767 6817
rect 4890 6808 4896 6820
rect 4948 6808 4954 6860
rect 5258 6808 5264 6860
rect 5316 6848 5322 6860
rect 5316 6820 5948 6848
rect 5316 6808 5322 6820
rect 3605 6783 3663 6789
rect 3605 6749 3617 6783
rect 3651 6780 3663 6783
rect 4065 6783 4123 6789
rect 3651 6752 4016 6780
rect 3651 6749 3663 6752
rect 3605 6743 3663 6749
rect 3620 6712 3648 6743
rect 3200 6684 3648 6712
rect 3200 6672 3206 6684
rect 1670 6604 1676 6656
rect 1728 6644 1734 6656
rect 1949 6647 2007 6653
rect 1949 6644 1961 6647
rect 1728 6616 1961 6644
rect 1728 6604 1734 6616
rect 1949 6613 1961 6616
rect 1995 6613 2007 6647
rect 1949 6607 2007 6613
rect 3878 6604 3884 6656
rect 3936 6604 3942 6656
rect 3988 6644 4016 6752
rect 4065 6749 4077 6783
rect 4111 6749 4123 6783
rect 4065 6743 4123 6749
rect 4154 6740 4160 6792
rect 4212 6780 4218 6792
rect 4341 6783 4399 6789
rect 4341 6780 4353 6783
rect 4212 6752 4353 6780
rect 4212 6740 4218 6752
rect 4341 6749 4353 6752
rect 4387 6749 4399 6783
rect 4341 6743 4399 6749
rect 4433 6783 4491 6789
rect 4433 6749 4445 6783
rect 4479 6749 4491 6783
rect 4433 6743 4491 6749
rect 4525 6783 4583 6789
rect 4525 6749 4537 6783
rect 4571 6749 4583 6783
rect 4525 6743 4583 6749
rect 5077 6783 5135 6789
rect 5077 6749 5089 6783
rect 5123 6780 5135 6783
rect 5350 6780 5356 6792
rect 5123 6752 5356 6780
rect 5123 6749 5135 6752
rect 5077 6743 5135 6749
rect 4246 6672 4252 6724
rect 4304 6672 4310 6724
rect 4448 6644 4476 6743
rect 3988 6616 4476 6644
rect 4540 6644 4568 6743
rect 5350 6740 5356 6752
rect 5408 6780 5414 6792
rect 5736 6789 5764 6820
rect 5920 6789 5948 6820
rect 7006 6808 7012 6860
rect 7064 6848 7070 6860
rect 7745 6851 7803 6857
rect 7745 6848 7757 6851
rect 7064 6820 7757 6848
rect 7064 6808 7070 6820
rect 7745 6817 7757 6820
rect 7791 6817 7803 6851
rect 7745 6811 7803 6817
rect 8478 6808 8484 6860
rect 8536 6808 8542 6860
rect 8680 6857 8708 6888
rect 8665 6851 8723 6857
rect 8665 6817 8677 6851
rect 8711 6817 8723 6851
rect 8665 6811 8723 6817
rect 9585 6851 9643 6857
rect 9585 6817 9597 6851
rect 9631 6848 9643 6851
rect 9766 6848 9772 6860
rect 9631 6820 9772 6848
rect 9631 6817 9643 6820
rect 9585 6811 9643 6817
rect 9766 6808 9772 6820
rect 9824 6808 9830 6860
rect 5628 6783 5686 6789
rect 5628 6780 5640 6783
rect 5408 6752 5640 6780
rect 5408 6740 5414 6752
rect 5628 6749 5640 6752
rect 5674 6749 5686 6783
rect 5628 6743 5686 6749
rect 5721 6783 5779 6789
rect 5721 6749 5733 6783
rect 5767 6749 5779 6783
rect 5721 6743 5779 6749
rect 5813 6783 5871 6789
rect 5813 6749 5825 6783
rect 5859 6749 5871 6783
rect 5813 6743 5871 6749
rect 5906 6783 5964 6789
rect 5906 6749 5918 6783
rect 5952 6749 5964 6783
rect 5906 6743 5964 6749
rect 7653 6783 7711 6789
rect 7653 6749 7665 6783
rect 7699 6780 7711 6783
rect 7834 6780 7840 6792
rect 7699 6752 7840 6780
rect 7699 6749 7711 6752
rect 7653 6743 7711 6749
rect 5644 6712 5672 6743
rect 5828 6712 5856 6743
rect 7834 6740 7840 6752
rect 7892 6740 7898 6792
rect 8018 6740 8024 6792
rect 8076 6780 8082 6792
rect 9217 6783 9275 6789
rect 9217 6780 9229 6783
rect 8076 6752 9229 6780
rect 8076 6740 8082 6752
rect 9217 6749 9229 6752
rect 9263 6749 9275 6783
rect 9217 6743 9275 6749
rect 6822 6712 6828 6724
rect 5644 6684 6828 6712
rect 6822 6672 6828 6684
rect 6880 6672 6886 6724
rect 10134 6672 10140 6724
rect 10192 6672 10198 6724
rect 11146 6672 11152 6724
rect 11204 6712 11210 6724
rect 11532 6721 11560 6888
rect 12158 6876 12164 6888
rect 12216 6916 12222 6928
rect 12621 6919 12679 6925
rect 12216 6888 12359 6916
rect 12216 6876 12222 6888
rect 11606 6808 11612 6860
rect 11664 6848 11670 6860
rect 12331 6848 12359 6888
rect 12621 6885 12633 6919
rect 12667 6916 12679 6919
rect 12894 6916 12900 6928
rect 12667 6888 12900 6916
rect 12667 6885 12679 6888
rect 12621 6879 12679 6885
rect 12894 6876 12900 6888
rect 12952 6876 12958 6928
rect 16025 6851 16083 6857
rect 11664 6820 12204 6848
rect 12331 6820 12388 6848
rect 11664 6808 11670 6820
rect 12176 6774 12204 6820
rect 12360 6789 12388 6820
rect 16025 6817 16037 6851
rect 16071 6848 16083 6851
rect 17126 6848 17132 6860
rect 16071 6820 17132 6848
rect 16071 6817 16083 6820
rect 16025 6811 16083 6817
rect 17126 6808 17132 6820
rect 17184 6808 17190 6860
rect 18046 6808 18052 6860
rect 18104 6808 18110 6860
rect 18138 6808 18144 6860
rect 18196 6848 18202 6860
rect 19245 6851 19303 6857
rect 19245 6848 19257 6851
rect 18196 6820 19257 6848
rect 18196 6808 18202 6820
rect 19245 6817 19257 6820
rect 19291 6848 19303 6851
rect 20806 6848 20812 6860
rect 19291 6820 20812 6848
rect 19291 6817 19303 6820
rect 19245 6811 19303 6817
rect 20806 6808 20812 6820
rect 20864 6808 20870 6860
rect 12348 6783 12406 6789
rect 12232 6777 12290 6783
rect 12232 6774 12244 6777
rect 12176 6746 12244 6774
rect 12232 6743 12244 6746
rect 12278 6743 12290 6777
rect 12348 6749 12360 6783
rect 12394 6749 12406 6783
rect 12348 6743 12406 6749
rect 12232 6737 12290 6743
rect 12434 6740 12440 6792
rect 12492 6740 12498 6792
rect 12618 6740 12624 6792
rect 12676 6740 12682 6792
rect 12894 6740 12900 6792
rect 12952 6740 12958 6792
rect 12989 6783 13047 6789
rect 12989 6749 13001 6783
rect 13035 6749 13047 6783
rect 16117 6783 16175 6789
rect 16117 6780 16129 6783
rect 12989 6743 13047 6749
rect 15672 6752 16129 6780
rect 11517 6715 11575 6721
rect 11517 6712 11529 6715
rect 11204 6684 11529 6712
rect 11204 6672 11210 6684
rect 11517 6681 11529 6684
rect 11563 6681 11575 6715
rect 11517 6675 11575 6681
rect 11606 6672 11612 6724
rect 11664 6712 11670 6724
rect 11701 6715 11759 6721
rect 11701 6712 11713 6715
rect 11664 6684 11713 6712
rect 11664 6672 11670 6684
rect 11701 6681 11713 6684
rect 11747 6681 11759 6715
rect 11701 6675 11759 6681
rect 11790 6672 11796 6724
rect 11848 6672 11854 6724
rect 11882 6672 11888 6724
rect 11940 6672 11946 6724
rect 12802 6672 12808 6724
rect 12860 6712 12866 6724
rect 13004 6712 13032 6743
rect 15672 6724 15700 6752
rect 16117 6749 16129 6752
rect 16163 6749 16175 6783
rect 16117 6743 16175 6749
rect 17405 6783 17463 6789
rect 17405 6749 17417 6783
rect 17451 6749 17463 6783
rect 17405 6743 17463 6749
rect 12860 6684 13032 6712
rect 12860 6672 12866 6684
rect 15654 6672 15660 6724
rect 15712 6672 15718 6724
rect 15841 6715 15899 6721
rect 15841 6681 15853 6715
rect 15887 6712 15899 6715
rect 16209 6715 16267 6721
rect 16209 6712 16221 6715
rect 15887 6684 16221 6712
rect 15887 6681 15899 6684
rect 15841 6675 15899 6681
rect 16209 6681 16221 6684
rect 16255 6681 16267 6715
rect 16209 6675 16267 6681
rect 16393 6715 16451 6721
rect 16393 6681 16405 6715
rect 16439 6712 16451 6715
rect 16574 6712 16580 6724
rect 16439 6684 16580 6712
rect 16439 6681 16451 6684
rect 16393 6675 16451 6681
rect 6181 6647 6239 6653
rect 6181 6644 6193 6647
rect 4540 6616 6193 6644
rect 6181 6613 6193 6616
rect 6227 6644 6239 6647
rect 6546 6644 6552 6656
rect 6227 6616 6552 6644
rect 6227 6613 6239 6616
rect 6181 6607 6239 6613
rect 6546 6604 6552 6616
rect 6604 6604 6610 6656
rect 7193 6647 7251 6653
rect 7193 6613 7205 6647
rect 7239 6644 7251 6647
rect 7282 6644 7288 6656
rect 7239 6616 7288 6644
rect 7239 6613 7251 6616
rect 7193 6607 7251 6613
rect 7282 6604 7288 6616
rect 7340 6604 7346 6656
rect 7558 6604 7564 6656
rect 7616 6604 7622 6656
rect 8021 6647 8079 6653
rect 8021 6613 8033 6647
rect 8067 6644 8079 6647
rect 8110 6644 8116 6656
rect 8067 6616 8116 6644
rect 8067 6613 8079 6616
rect 8021 6607 8079 6613
rect 8110 6604 8116 6616
rect 8168 6604 8174 6656
rect 8389 6647 8447 6653
rect 8389 6613 8401 6647
rect 8435 6644 8447 6647
rect 9582 6644 9588 6656
rect 8435 6616 9588 6644
rect 8435 6613 8447 6616
rect 8389 6607 8447 6613
rect 9582 6604 9588 6616
rect 9640 6604 9646 6656
rect 11808 6644 11836 6672
rect 12250 6644 12256 6656
rect 11808 6616 12256 6644
rect 12250 6604 12256 6616
rect 12308 6604 12314 6656
rect 13722 6604 13728 6656
rect 13780 6644 13786 6656
rect 15856 6644 15884 6675
rect 16574 6672 16580 6684
rect 16632 6712 16638 6724
rect 17218 6712 17224 6724
rect 16632 6684 17224 6712
rect 16632 6672 16638 6684
rect 17218 6672 17224 6684
rect 17276 6672 17282 6724
rect 17420 6712 17448 6743
rect 19058 6740 19064 6792
rect 19116 6740 19122 6792
rect 19610 6740 19616 6792
rect 19668 6740 19674 6792
rect 18417 6715 18475 6721
rect 18417 6712 18429 6715
rect 17420 6684 18429 6712
rect 18417 6681 18429 6684
rect 18463 6681 18475 6715
rect 18417 6675 18475 6681
rect 19978 6672 19984 6724
rect 20036 6672 20042 6724
rect 13780 6616 15884 6644
rect 13780 6604 13786 6616
rect 17310 6604 17316 6656
rect 17368 6604 17374 6656
rect 17494 6604 17500 6656
rect 17552 6604 17558 6656
rect 1104 6554 25208 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 25208 6554
rect 1104 6480 25208 6502
rect 2498 6400 2504 6452
rect 2556 6440 2562 6452
rect 2556 6412 3096 6440
rect 2556 6400 2562 6412
rect 1670 6332 1676 6384
rect 1728 6332 1734 6384
rect 3068 6372 3096 6412
rect 3142 6400 3148 6452
rect 3200 6400 3206 6452
rect 3605 6443 3663 6449
rect 3605 6409 3617 6443
rect 3651 6440 3663 6443
rect 3786 6440 3792 6452
rect 3651 6412 3792 6440
rect 3651 6409 3663 6412
rect 3605 6403 3663 6409
rect 3786 6400 3792 6412
rect 3844 6400 3850 6452
rect 4246 6400 4252 6452
rect 4304 6440 4310 6452
rect 5442 6440 5448 6452
rect 4304 6412 5448 6440
rect 4304 6400 4310 6412
rect 5442 6400 5448 6412
rect 5500 6400 5506 6452
rect 5994 6400 6000 6452
rect 6052 6440 6058 6452
rect 6733 6443 6791 6449
rect 6733 6440 6745 6443
rect 6052 6412 6745 6440
rect 6052 6400 6058 6412
rect 6733 6409 6745 6412
rect 6779 6409 6791 6443
rect 6733 6403 6791 6409
rect 6822 6400 6828 6452
rect 6880 6400 6886 6452
rect 10134 6400 10140 6452
rect 10192 6440 10198 6452
rect 10505 6443 10563 6449
rect 10505 6440 10517 6443
rect 10192 6412 10517 6440
rect 10192 6400 10198 6412
rect 10505 6409 10517 6412
rect 10551 6409 10563 6443
rect 10505 6403 10563 6409
rect 10870 6400 10876 6452
rect 10928 6440 10934 6452
rect 11790 6440 11796 6452
rect 10928 6412 11796 6440
rect 10928 6400 10934 6412
rect 11790 6400 11796 6412
rect 11848 6400 11854 6452
rect 13173 6443 13231 6449
rect 13173 6409 13185 6443
rect 13219 6409 13231 6443
rect 13173 6403 13231 6409
rect 14369 6443 14427 6449
rect 14369 6409 14381 6443
rect 14415 6440 14427 6443
rect 15654 6440 15660 6452
rect 14415 6412 15660 6440
rect 14415 6409 14427 6412
rect 14369 6403 14427 6409
rect 3068 6344 3924 6372
rect 2806 6276 2912 6304
rect 2884 6248 2912 6276
rect 1394 6196 1400 6248
rect 1452 6196 1458 6248
rect 2866 6196 2872 6248
rect 2924 6196 2930 6248
rect 3602 6196 3608 6248
rect 3660 6236 3666 6248
rect 3896 6245 3924 6344
rect 7745 6307 7803 6313
rect 7745 6273 7757 6307
rect 7791 6304 7803 6307
rect 8018 6304 8024 6316
rect 7791 6276 8024 6304
rect 7791 6273 7803 6276
rect 7745 6267 7803 6273
rect 8018 6264 8024 6276
rect 8076 6264 8082 6316
rect 8110 6264 8116 6316
rect 8168 6264 8174 6316
rect 9030 6264 9036 6316
rect 9088 6304 9094 6316
rect 9140 6304 9168 6358
rect 9582 6332 9588 6384
rect 9640 6372 9646 6384
rect 12529 6375 12587 6381
rect 9640 6344 12359 6372
rect 9640 6332 9646 6344
rect 10134 6304 10140 6316
rect 9088 6276 10140 6304
rect 9088 6264 9094 6276
rect 10134 6264 10140 6276
rect 10192 6264 10198 6316
rect 10318 6264 10324 6316
rect 10376 6304 10382 6316
rect 10413 6307 10471 6313
rect 10413 6304 10425 6307
rect 10376 6276 10425 6304
rect 10376 6264 10382 6276
rect 10413 6273 10425 6276
rect 10459 6273 10471 6307
rect 10413 6267 10471 6273
rect 11517 6307 11575 6313
rect 11517 6273 11529 6307
rect 11563 6273 11575 6307
rect 11517 6267 11575 6273
rect 3697 6239 3755 6245
rect 3697 6236 3709 6239
rect 3660 6208 3709 6236
rect 3660 6196 3666 6208
rect 3697 6205 3709 6208
rect 3743 6205 3755 6239
rect 3697 6199 3755 6205
rect 3881 6239 3939 6245
rect 3881 6205 3893 6239
rect 3927 6236 3939 6239
rect 6454 6236 6460 6248
rect 3927 6208 6460 6236
rect 3927 6205 3939 6208
rect 3881 6199 3939 6205
rect 6454 6196 6460 6208
rect 6512 6236 6518 6248
rect 6917 6239 6975 6245
rect 6917 6236 6929 6239
rect 6512 6208 6929 6236
rect 6512 6196 6518 6208
rect 6917 6205 6929 6208
rect 6963 6205 6975 6239
rect 11532 6236 11560 6267
rect 11698 6264 11704 6316
rect 11756 6264 11762 6316
rect 12331 6310 12359 6344
rect 12529 6341 12541 6375
rect 12575 6372 12587 6375
rect 12802 6372 12808 6384
rect 12575 6344 12808 6372
rect 12575 6341 12587 6344
rect 12529 6335 12587 6341
rect 12802 6332 12808 6344
rect 12860 6332 12866 6384
rect 13005 6375 13063 6381
rect 13005 6372 13017 6375
rect 12912 6344 13017 6372
rect 12428 6313 12486 6319
rect 12428 6310 12440 6313
rect 12331 6282 12440 6310
rect 12428 6279 12440 6282
rect 12474 6279 12486 6313
rect 12428 6273 12486 6279
rect 11882 6236 11888 6248
rect 11532 6208 11888 6236
rect 6917 6199 6975 6205
rect 11882 6196 11888 6208
rect 11940 6196 11946 6248
rect 3234 6060 3240 6112
rect 3292 6060 3298 6112
rect 6365 6103 6423 6109
rect 6365 6069 6377 6103
rect 6411 6100 6423 6103
rect 6546 6100 6552 6112
rect 6411 6072 6552 6100
rect 6411 6069 6423 6072
rect 6365 6063 6423 6069
rect 6546 6060 6552 6072
rect 6604 6060 6610 6112
rect 11609 6103 11667 6109
rect 11609 6069 11621 6103
rect 11655 6100 11667 6103
rect 11698 6100 11704 6112
rect 11655 6072 11704 6100
rect 11655 6069 11667 6072
rect 11609 6063 11667 6069
rect 11698 6060 11704 6072
rect 11756 6060 11762 6112
rect 12452 6100 12480 6273
rect 12710 6264 12716 6316
rect 12768 6304 12774 6316
rect 12912 6304 12940 6344
rect 13005 6341 13017 6344
rect 13051 6341 13063 6375
rect 13188 6372 13216 6403
rect 15654 6400 15660 6412
rect 15712 6400 15718 6452
rect 16482 6400 16488 6452
rect 16540 6400 16546 6452
rect 17494 6440 17500 6452
rect 16592 6412 17500 6440
rect 14185 6375 14243 6381
rect 14185 6372 14197 6375
rect 13188 6344 14197 6372
rect 13005 6335 13063 6341
rect 14185 6341 14197 6344
rect 14231 6341 14243 6375
rect 14185 6335 14243 6341
rect 14734 6332 14740 6384
rect 14792 6372 14798 6384
rect 15013 6375 15071 6381
rect 15013 6372 15025 6375
rect 14792 6344 15025 6372
rect 14792 6332 14798 6344
rect 15013 6341 15025 6344
rect 15059 6341 15071 6375
rect 16347 6375 16405 6381
rect 16347 6372 16359 6375
rect 15013 6335 15071 6341
rect 15764 6344 16359 6372
rect 12768 6276 12940 6304
rect 13449 6307 13507 6313
rect 12768 6264 12774 6276
rect 13449 6273 13461 6307
rect 13495 6273 13507 6307
rect 13449 6267 13507 6273
rect 13464 6236 13492 6267
rect 13630 6264 13636 6316
rect 13688 6264 13694 6316
rect 13722 6264 13728 6316
rect 13780 6264 13786 6316
rect 14001 6307 14059 6313
rect 14001 6273 14013 6307
rect 14047 6273 14059 6307
rect 14001 6267 14059 6273
rect 14016 6236 14044 6267
rect 14550 6264 14556 6316
rect 14608 6304 14614 6316
rect 14829 6307 14887 6313
rect 14829 6304 14841 6307
rect 14608 6276 14841 6304
rect 14608 6264 14614 6276
rect 14829 6273 14841 6276
rect 14875 6273 14887 6307
rect 14829 6267 14887 6273
rect 12728 6208 14044 6236
rect 14844 6236 14872 6267
rect 14918 6264 14924 6316
rect 14976 6264 14982 6316
rect 15197 6307 15255 6313
rect 15197 6273 15209 6307
rect 15243 6304 15255 6307
rect 15565 6307 15623 6313
rect 15565 6304 15577 6307
rect 15243 6276 15577 6304
rect 15243 6273 15255 6276
rect 15197 6267 15255 6273
rect 15565 6273 15577 6276
rect 15611 6304 15623 6307
rect 15654 6304 15660 6316
rect 15611 6276 15660 6304
rect 15611 6273 15623 6276
rect 15565 6267 15623 6273
rect 15654 6264 15660 6276
rect 15712 6264 15718 6316
rect 15764 6313 15792 6344
rect 16347 6341 16359 6344
rect 16393 6372 16405 6375
rect 16500 6372 16528 6400
rect 16393 6344 16528 6372
rect 16393 6341 16405 6344
rect 16347 6335 16405 6341
rect 15749 6307 15807 6313
rect 15749 6273 15761 6307
rect 15795 6273 15807 6307
rect 15749 6267 15807 6273
rect 16025 6307 16083 6313
rect 16025 6273 16037 6307
rect 16071 6273 16083 6307
rect 16025 6267 16083 6273
rect 15470 6236 15476 6248
rect 14844 6208 15476 6236
rect 12728 6177 12756 6208
rect 15470 6196 15476 6208
rect 15528 6196 15534 6248
rect 16040 6236 16068 6267
rect 16114 6264 16120 6316
rect 16172 6264 16178 6316
rect 16206 6264 16212 6316
rect 16264 6264 16270 6316
rect 16485 6307 16543 6313
rect 16485 6273 16497 6307
rect 16531 6304 16543 6307
rect 16592 6304 16620 6412
rect 17494 6400 17500 6412
rect 17552 6400 17558 6452
rect 19610 6400 19616 6452
rect 19668 6440 19674 6452
rect 20533 6443 20591 6449
rect 20533 6440 20545 6443
rect 19668 6412 20545 6440
rect 19668 6400 19674 6412
rect 20533 6409 20545 6412
rect 20579 6409 20591 6443
rect 20533 6403 20591 6409
rect 20714 6400 20720 6452
rect 20772 6440 20778 6452
rect 20993 6443 21051 6449
rect 20993 6440 21005 6443
rect 20772 6412 21005 6440
rect 20772 6400 20778 6412
rect 20993 6409 21005 6412
rect 21039 6409 21051 6443
rect 20993 6403 21051 6409
rect 21542 6400 21548 6452
rect 21600 6400 21606 6452
rect 18782 6372 18788 6384
rect 18078 6344 18788 6372
rect 18782 6332 18788 6344
rect 18840 6372 18846 6384
rect 18840 6344 19090 6372
rect 18840 6332 18846 6344
rect 16531 6276 16620 6304
rect 16531 6273 16543 6276
rect 16485 6267 16543 6273
rect 16666 6264 16672 6316
rect 16724 6264 16730 6316
rect 20901 6307 20959 6313
rect 20901 6273 20913 6307
rect 20947 6273 20959 6307
rect 20901 6267 20959 6273
rect 16390 6236 16396 6248
rect 15580 6208 16396 6236
rect 12713 6171 12771 6177
rect 12713 6137 12725 6171
rect 12759 6137 12771 6171
rect 12713 6131 12771 6137
rect 14642 6128 14648 6180
rect 14700 6128 14706 6180
rect 15580 6177 15608 6208
rect 16390 6196 16396 6208
rect 16448 6196 16454 6248
rect 17037 6239 17095 6245
rect 17037 6236 17049 6239
rect 16592 6208 17049 6236
rect 15565 6171 15623 6177
rect 15565 6137 15577 6171
rect 15611 6137 15623 6171
rect 15565 6131 15623 6137
rect 15841 6171 15899 6177
rect 15841 6137 15853 6171
rect 15887 6168 15899 6171
rect 16592 6168 16620 6208
rect 17037 6205 17049 6208
rect 17083 6205 17095 6239
rect 17037 6199 17095 6205
rect 17494 6196 17500 6248
rect 17552 6236 17558 6248
rect 20073 6239 20131 6245
rect 20073 6236 20085 6239
rect 17552 6208 20085 6236
rect 17552 6196 17558 6208
rect 20073 6205 20085 6208
rect 20119 6205 20131 6239
rect 20073 6199 20131 6205
rect 20441 6239 20499 6245
rect 20441 6205 20453 6239
rect 20487 6236 20499 6239
rect 20806 6236 20812 6248
rect 20487 6208 20812 6236
rect 20487 6205 20499 6208
rect 20441 6199 20499 6205
rect 20806 6196 20812 6208
rect 20864 6196 20870 6248
rect 15887 6140 16620 6168
rect 15887 6137 15899 6140
rect 15841 6131 15899 6137
rect 18046 6128 18052 6180
rect 18104 6168 18110 6180
rect 18463 6171 18521 6177
rect 18463 6168 18475 6171
rect 18104 6140 18475 6168
rect 18104 6128 18110 6140
rect 18463 6137 18475 6140
rect 18509 6137 18521 6171
rect 18463 6131 18521 6137
rect 18647 6171 18705 6177
rect 18647 6137 18659 6171
rect 18693 6168 18705 6171
rect 18966 6168 18972 6180
rect 18693 6140 18972 6168
rect 18693 6137 18705 6140
rect 18647 6131 18705 6137
rect 18966 6128 18972 6140
rect 19024 6128 19030 6180
rect 12989 6103 13047 6109
rect 12989 6100 13001 6103
rect 12452 6072 13001 6100
rect 12989 6069 13001 6072
rect 13035 6100 13047 6103
rect 13078 6100 13084 6112
rect 13035 6072 13084 6100
rect 13035 6069 13047 6072
rect 12989 6063 13047 6069
rect 13078 6060 13084 6072
rect 13136 6060 13142 6112
rect 13262 6060 13268 6112
rect 13320 6060 13326 6112
rect 18782 6060 18788 6112
rect 18840 6100 18846 6112
rect 20916 6100 20944 6267
rect 21358 6264 21364 6316
rect 21416 6304 21422 6316
rect 24670 6304 24676 6316
rect 21416 6276 24676 6304
rect 21416 6264 21422 6276
rect 24670 6264 24676 6276
rect 24728 6264 24734 6316
rect 21082 6196 21088 6248
rect 21140 6196 21146 6248
rect 18840 6072 20944 6100
rect 18840 6060 18846 6072
rect 1104 6010 25208 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 25208 6010
rect 1104 5936 25208 5958
rect 1752 5899 1810 5905
rect 1752 5865 1764 5899
rect 1798 5896 1810 5899
rect 3234 5896 3240 5908
rect 1798 5868 3240 5896
rect 1798 5865 1810 5868
rect 1752 5859 1810 5865
rect 3234 5856 3240 5868
rect 3292 5856 3298 5908
rect 5077 5899 5135 5905
rect 5077 5865 5089 5899
rect 5123 5896 5135 5899
rect 5350 5896 5356 5908
rect 5123 5868 5356 5896
rect 5123 5865 5135 5868
rect 5077 5859 5135 5865
rect 5350 5856 5356 5868
rect 5408 5856 5414 5908
rect 7558 5856 7564 5908
rect 7616 5896 7622 5908
rect 8665 5899 8723 5905
rect 8665 5896 8677 5899
rect 7616 5868 8677 5896
rect 7616 5856 7622 5868
rect 8665 5865 8677 5868
rect 8711 5865 8723 5899
rect 8665 5859 8723 5865
rect 1394 5720 1400 5772
rect 1452 5760 1458 5772
rect 1489 5763 1547 5769
rect 1489 5760 1501 5763
rect 1452 5732 1501 5760
rect 1452 5720 1458 5732
rect 1489 5729 1501 5732
rect 1535 5760 1547 5763
rect 3694 5760 3700 5772
rect 1535 5732 3700 5760
rect 1535 5729 1547 5732
rect 1489 5723 1547 5729
rect 3694 5720 3700 5732
rect 3752 5760 3758 5772
rect 4614 5760 4620 5772
rect 3752 5732 4620 5760
rect 3752 5720 3758 5732
rect 4614 5720 4620 5732
rect 4672 5720 4678 5772
rect 6546 5720 6552 5772
rect 6604 5720 6610 5772
rect 6825 5763 6883 5769
rect 6825 5729 6837 5763
rect 6871 5760 6883 5763
rect 6917 5763 6975 5769
rect 6917 5760 6929 5763
rect 6871 5732 6929 5760
rect 6871 5729 6883 5732
rect 6825 5723 6883 5729
rect 6917 5729 6929 5732
rect 6963 5760 6975 5763
rect 8018 5760 8024 5772
rect 6963 5732 8024 5760
rect 6963 5729 6975 5732
rect 6917 5723 6975 5729
rect 8018 5720 8024 5732
rect 8076 5720 8082 5772
rect 2866 5652 2872 5704
rect 2924 5652 2930 5704
rect 7282 5652 7288 5704
rect 7340 5652 7346 5704
rect 8680 5692 8708 5859
rect 10410 5856 10416 5908
rect 10468 5896 10474 5908
rect 10870 5896 10876 5908
rect 10468 5868 10876 5896
rect 10468 5856 10474 5868
rect 10870 5856 10876 5868
rect 10928 5856 10934 5908
rect 11330 5896 11336 5908
rect 11164 5868 11336 5896
rect 10502 5788 10508 5840
rect 10560 5828 10566 5840
rect 11054 5828 11060 5840
rect 10560 5800 11060 5828
rect 10560 5788 10566 5800
rect 11054 5788 11060 5800
rect 11112 5788 11118 5840
rect 10229 5763 10287 5769
rect 10229 5729 10241 5763
rect 10275 5760 10287 5763
rect 11164 5760 11192 5868
rect 11330 5856 11336 5868
rect 11388 5856 11394 5908
rect 13265 5899 13323 5905
rect 13265 5865 13277 5899
rect 13311 5896 13323 5899
rect 13630 5896 13636 5908
rect 13311 5868 13636 5896
rect 13311 5865 13323 5868
rect 13265 5859 13323 5865
rect 13630 5856 13636 5868
rect 13688 5856 13694 5908
rect 16206 5856 16212 5908
rect 16264 5896 16270 5908
rect 16301 5899 16359 5905
rect 16301 5896 16313 5899
rect 16264 5868 16313 5896
rect 16264 5856 16270 5868
rect 16301 5865 16313 5868
rect 16347 5865 16359 5899
rect 16301 5859 16359 5865
rect 17129 5899 17187 5905
rect 17129 5865 17141 5899
rect 17175 5896 17187 5899
rect 17494 5896 17500 5908
rect 17175 5868 17500 5896
rect 17175 5865 17187 5868
rect 17129 5859 17187 5865
rect 17494 5856 17500 5868
rect 17552 5856 17558 5908
rect 21082 5896 21088 5908
rect 18616 5868 21088 5896
rect 11882 5788 11888 5840
rect 11940 5828 11946 5840
rect 12253 5831 12311 5837
rect 12253 5828 12265 5831
rect 11940 5800 12265 5828
rect 11940 5788 11946 5800
rect 12253 5797 12265 5800
rect 12299 5797 12311 5831
rect 12253 5791 12311 5797
rect 15470 5788 15476 5840
rect 15528 5828 15534 5840
rect 15528 5800 16206 5828
rect 15528 5788 15534 5800
rect 10275 5732 11192 5760
rect 11793 5763 11851 5769
rect 10275 5729 10287 5732
rect 10229 5723 10287 5729
rect 11793 5729 11805 5763
rect 11839 5760 11851 5763
rect 12161 5763 12219 5769
rect 12161 5760 12173 5763
rect 11839 5732 12173 5760
rect 11839 5729 11851 5732
rect 11793 5723 11851 5729
rect 12161 5729 12173 5732
rect 12207 5729 12219 5763
rect 15657 5763 15715 5769
rect 15657 5760 15669 5763
rect 12161 5723 12219 5729
rect 14844 5732 15669 5760
rect 10597 5695 10655 5701
rect 10597 5692 10609 5695
rect 8680 5664 10609 5692
rect 10597 5661 10609 5664
rect 10643 5661 10655 5695
rect 10597 5655 10655 5661
rect 6086 5584 6092 5636
rect 6144 5624 6150 5636
rect 7006 5624 7012 5636
rect 6144 5596 7012 5624
rect 6144 5584 6150 5596
rect 7006 5584 7012 5596
rect 7064 5584 7070 5636
rect 9030 5624 9036 5636
rect 8326 5596 9036 5624
rect 9030 5584 9036 5596
rect 9088 5584 9094 5636
rect 10410 5584 10416 5636
rect 10468 5584 10474 5636
rect 10502 5584 10508 5636
rect 10560 5584 10566 5636
rect 3237 5559 3295 5565
rect 3237 5525 3249 5559
rect 3283 5556 3295 5559
rect 3602 5556 3608 5568
rect 3283 5528 3608 5556
rect 3283 5525 3295 5528
rect 3237 5519 3295 5525
rect 3602 5516 3608 5528
rect 3660 5516 3666 5568
rect 10612 5556 10640 5655
rect 10870 5652 10876 5704
rect 10928 5652 10934 5704
rect 11146 5692 11152 5704
rect 10980 5664 11152 5692
rect 10781 5627 10839 5633
rect 10781 5593 10793 5627
rect 10827 5624 10839 5627
rect 10980 5624 11008 5664
rect 11146 5652 11152 5664
rect 11204 5652 11210 5704
rect 11241 5695 11299 5701
rect 11241 5661 11253 5695
rect 11287 5661 11299 5695
rect 11241 5655 11299 5661
rect 10827 5596 11008 5624
rect 10827 5593 10839 5596
rect 10781 5587 10839 5593
rect 11054 5584 11060 5636
rect 11112 5584 11118 5636
rect 11256 5568 11284 5655
rect 11698 5652 11704 5704
rect 11756 5652 11762 5704
rect 11992 5664 12434 5692
rect 11330 5584 11336 5636
rect 11388 5624 11394 5636
rect 11992 5624 12020 5664
rect 12406 5624 12434 5664
rect 12802 5652 12808 5704
rect 12860 5692 12866 5704
rect 13265 5695 13323 5701
rect 13265 5692 13277 5695
rect 12860 5664 13277 5692
rect 12860 5652 12866 5664
rect 13265 5661 13277 5664
rect 13311 5661 13323 5695
rect 14550 5692 14556 5704
rect 13265 5655 13323 5661
rect 13648 5664 14556 5692
rect 12621 5627 12679 5633
rect 12621 5624 12633 5627
rect 11388 5596 12020 5624
rect 12084 5596 12296 5624
rect 12406 5596 12633 5624
rect 11388 5584 11394 5596
rect 11238 5556 11244 5568
rect 10612 5528 11244 5556
rect 11238 5516 11244 5528
rect 11296 5516 11302 5568
rect 11425 5559 11483 5565
rect 11425 5525 11437 5559
rect 11471 5556 11483 5559
rect 11882 5556 11888 5568
rect 11471 5528 11888 5556
rect 11471 5525 11483 5528
rect 11425 5519 11483 5525
rect 11882 5516 11888 5528
rect 11940 5516 11946 5568
rect 12084 5565 12112 5596
rect 12069 5559 12127 5565
rect 12069 5525 12081 5559
rect 12115 5525 12127 5559
rect 12268 5556 12296 5596
rect 12621 5593 12633 5596
rect 12667 5593 12679 5627
rect 12621 5587 12679 5593
rect 12989 5627 13047 5633
rect 12989 5593 13001 5627
rect 13035 5593 13047 5627
rect 12989 5587 13047 5593
rect 12710 5556 12716 5568
rect 12268 5528 12716 5556
rect 12069 5519 12127 5525
rect 12710 5516 12716 5528
rect 12768 5556 12774 5568
rect 13004 5556 13032 5587
rect 13078 5584 13084 5636
rect 13136 5624 13142 5636
rect 13173 5627 13231 5633
rect 13173 5624 13185 5627
rect 13136 5596 13185 5624
rect 13136 5584 13142 5596
rect 13173 5593 13185 5596
rect 13219 5624 13231 5627
rect 13648 5624 13676 5664
rect 14550 5652 14556 5664
rect 14608 5652 14614 5704
rect 14734 5652 14740 5704
rect 14792 5652 14798 5704
rect 14844 5633 14872 5732
rect 15657 5729 15669 5732
rect 15703 5760 15715 5763
rect 15703 5732 16068 5760
rect 15703 5729 15715 5732
rect 15657 5723 15715 5729
rect 14918 5652 14924 5704
rect 14976 5652 14982 5704
rect 15289 5695 15347 5701
rect 15289 5661 15301 5695
rect 15335 5661 15347 5695
rect 15289 5655 15347 5661
rect 15749 5695 15807 5701
rect 15749 5661 15761 5695
rect 15795 5661 15807 5695
rect 15749 5655 15807 5661
rect 13219 5596 13676 5624
rect 14829 5627 14887 5633
rect 13219 5593 13231 5596
rect 13173 5587 13231 5593
rect 14829 5593 14841 5627
rect 14875 5593 14887 5627
rect 15304 5624 15332 5655
rect 15562 5624 15568 5636
rect 14829 5587 14887 5593
rect 15120 5596 15568 5624
rect 12768 5528 13032 5556
rect 12768 5516 12774 5528
rect 13630 5516 13636 5568
rect 13688 5556 13694 5568
rect 14642 5556 14648 5568
rect 13688 5528 14648 5556
rect 13688 5516 13694 5528
rect 14642 5516 14648 5528
rect 14700 5556 14706 5568
rect 14844 5556 14872 5587
rect 15120 5565 15148 5596
rect 15562 5584 15568 5596
rect 15620 5624 15626 5636
rect 15764 5624 15792 5655
rect 15930 5652 15936 5704
rect 15988 5652 15994 5704
rect 16040 5701 16068 5732
rect 16178 5701 16206 5800
rect 16390 5788 16396 5840
rect 16448 5828 16454 5840
rect 16448 5800 17172 5828
rect 16448 5788 16454 5800
rect 16666 5720 16672 5772
rect 16724 5720 16730 5772
rect 16025 5695 16083 5701
rect 16025 5661 16037 5695
rect 16071 5661 16083 5695
rect 16025 5655 16083 5661
rect 16163 5695 16221 5701
rect 16163 5661 16175 5695
rect 16209 5661 16221 5695
rect 16163 5655 16221 5661
rect 16574 5652 16580 5704
rect 16632 5652 16638 5704
rect 17144 5701 17172 5800
rect 17218 5788 17224 5840
rect 17276 5828 17282 5840
rect 17276 5800 17540 5828
rect 17276 5788 17282 5800
rect 17310 5720 17316 5772
rect 17368 5760 17374 5772
rect 17368 5732 17448 5760
rect 17368 5720 17374 5732
rect 17420 5701 17448 5732
rect 17512 5701 17540 5800
rect 18509 5763 18567 5769
rect 18509 5729 18521 5763
rect 18555 5760 18567 5763
rect 18616 5760 18644 5868
rect 21082 5856 21088 5868
rect 21140 5856 21146 5908
rect 19061 5831 19119 5837
rect 19061 5797 19073 5831
rect 19107 5797 19119 5831
rect 19061 5791 19119 5797
rect 18555 5732 18644 5760
rect 19076 5760 19104 5791
rect 20717 5763 20775 5769
rect 20717 5760 20729 5763
rect 19076 5732 20729 5760
rect 18555 5729 18567 5732
rect 18509 5723 18567 5729
rect 20717 5729 20729 5732
rect 20763 5729 20775 5763
rect 20717 5723 20775 5729
rect 17129 5695 17187 5701
rect 17129 5661 17141 5695
rect 17175 5661 17187 5695
rect 17129 5655 17187 5661
rect 17405 5695 17463 5701
rect 17405 5661 17417 5695
rect 17451 5661 17463 5695
rect 17512 5695 17591 5701
rect 17512 5664 17545 5695
rect 17405 5655 17463 5661
rect 17533 5661 17545 5664
rect 17579 5692 17591 5695
rect 18524 5692 18552 5723
rect 20806 5720 20812 5772
rect 20864 5760 20870 5772
rect 21085 5763 21143 5769
rect 21085 5760 21097 5763
rect 20864 5732 21097 5760
rect 20864 5720 20870 5732
rect 21085 5729 21097 5732
rect 21131 5760 21143 5763
rect 21818 5760 21824 5772
rect 21131 5732 21824 5760
rect 21131 5729 21143 5732
rect 21085 5723 21143 5729
rect 21818 5720 21824 5732
rect 21876 5720 21882 5772
rect 17579 5664 18552 5692
rect 18601 5695 18659 5701
rect 17579 5661 17591 5664
rect 17533 5655 17591 5661
rect 18601 5661 18613 5695
rect 18647 5692 18659 5695
rect 19291 5695 19349 5701
rect 19291 5692 19303 5695
rect 18647 5664 19303 5692
rect 18647 5661 18659 5664
rect 18601 5655 18659 5661
rect 19291 5661 19303 5664
rect 19337 5692 19349 5695
rect 19518 5692 19524 5704
rect 19337 5664 19524 5692
rect 19337 5661 19349 5664
rect 19291 5655 19349 5661
rect 19518 5652 19524 5664
rect 19576 5652 19582 5704
rect 17313 5627 17371 5633
rect 17313 5624 17325 5627
rect 15620 5596 15792 5624
rect 16316 5596 17325 5624
rect 15620 5584 15626 5596
rect 14700 5528 14872 5556
rect 15105 5559 15163 5565
rect 14700 5516 14706 5528
rect 15105 5525 15117 5559
rect 15151 5525 15163 5559
rect 15105 5519 15163 5525
rect 15286 5516 15292 5568
rect 15344 5556 15350 5568
rect 15381 5559 15439 5565
rect 15381 5556 15393 5559
rect 15344 5528 15393 5556
rect 15344 5516 15350 5528
rect 15381 5525 15393 5528
rect 15427 5525 15439 5559
rect 15381 5519 15439 5525
rect 15470 5516 15476 5568
rect 15528 5516 15534 5568
rect 15657 5559 15715 5565
rect 15657 5525 15669 5559
rect 15703 5556 15715 5559
rect 16114 5556 16120 5568
rect 15703 5528 16120 5556
rect 15703 5525 15715 5528
rect 15657 5519 15715 5525
rect 16114 5516 16120 5528
rect 16172 5556 16178 5568
rect 16316 5556 16344 5596
rect 17313 5593 17325 5596
rect 17359 5593 17371 5627
rect 18782 5624 18788 5636
rect 17313 5587 17371 5593
rect 18524 5596 18788 5624
rect 16172 5528 16344 5556
rect 16945 5559 17003 5565
rect 16172 5516 16178 5528
rect 16945 5525 16957 5559
rect 16991 5556 17003 5559
rect 18524 5556 18552 5596
rect 18782 5584 18788 5596
rect 18840 5584 18846 5636
rect 19978 5584 19984 5636
rect 20036 5584 20042 5636
rect 16991 5528 18552 5556
rect 16991 5525 17003 5528
rect 16945 5519 17003 5525
rect 18690 5516 18696 5568
rect 18748 5516 18754 5568
rect 1104 5466 25208 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 25208 5466
rect 1104 5392 25208 5414
rect 5258 5312 5264 5364
rect 5316 5352 5322 5364
rect 5445 5355 5503 5361
rect 5445 5352 5457 5355
rect 5316 5324 5457 5352
rect 5316 5312 5322 5324
rect 5445 5321 5457 5324
rect 5491 5321 5503 5355
rect 10318 5352 10324 5364
rect 5445 5315 5503 5321
rect 6748 5324 10324 5352
rect 3878 5244 3884 5296
rect 3936 5284 3942 5296
rect 3973 5287 4031 5293
rect 3973 5284 3985 5287
rect 3936 5256 3985 5284
rect 3936 5244 3942 5256
rect 3973 5253 3985 5256
rect 4019 5253 4031 5287
rect 6086 5284 6092 5296
rect 5198 5270 6092 5284
rect 3973 5247 4031 5253
rect 5184 5256 6092 5270
rect 3694 5176 3700 5228
rect 3752 5176 3758 5228
rect 2866 5108 2872 5160
rect 2924 5148 2930 5160
rect 5184 5148 5212 5256
rect 6086 5244 6092 5256
rect 6144 5244 6150 5296
rect 6748 5293 6776 5324
rect 10318 5312 10324 5324
rect 10376 5312 10382 5364
rect 11054 5312 11060 5364
rect 11112 5352 11118 5364
rect 13449 5355 13507 5361
rect 13449 5352 13461 5355
rect 11112 5324 13461 5352
rect 11112 5312 11118 5324
rect 13449 5321 13461 5324
rect 13495 5352 13507 5355
rect 14734 5352 14740 5364
rect 13495 5324 14740 5352
rect 13495 5321 13507 5324
rect 13449 5315 13507 5321
rect 6733 5287 6791 5293
rect 6733 5253 6745 5287
rect 6779 5253 6791 5287
rect 6733 5247 6791 5253
rect 9030 5244 9036 5296
rect 9088 5244 9094 5296
rect 9723 5287 9781 5293
rect 9723 5253 9735 5287
rect 9769 5284 9781 5287
rect 9858 5284 9864 5296
rect 9769 5256 9864 5284
rect 9769 5253 9781 5256
rect 9723 5247 9781 5253
rect 9858 5244 9864 5256
rect 9916 5244 9922 5296
rect 12250 5244 12256 5296
rect 12308 5284 12314 5296
rect 13541 5287 13599 5293
rect 13541 5284 13553 5287
rect 12308 5256 13553 5284
rect 12308 5244 12314 5256
rect 13541 5253 13553 5256
rect 13587 5284 13599 5287
rect 14001 5287 14059 5293
rect 14001 5284 14013 5287
rect 13587 5256 14013 5284
rect 13587 5253 13599 5256
rect 13541 5247 13599 5253
rect 14001 5253 14013 5256
rect 14047 5253 14059 5287
rect 14001 5247 14059 5253
rect 14200 5247 14228 5324
rect 14734 5312 14740 5324
rect 14792 5312 14798 5364
rect 15286 5312 15292 5364
rect 15344 5352 15350 5364
rect 15930 5352 15936 5364
rect 15344 5324 15936 5352
rect 15344 5312 15350 5324
rect 15930 5312 15936 5324
rect 15988 5312 15994 5364
rect 16025 5355 16083 5361
rect 16025 5321 16037 5355
rect 16071 5352 16083 5355
rect 16666 5352 16672 5364
rect 16071 5324 16672 5352
rect 16071 5321 16083 5324
rect 16025 5315 16083 5321
rect 16666 5312 16672 5324
rect 16724 5312 16730 5364
rect 19889 5355 19947 5361
rect 19889 5321 19901 5355
rect 19935 5352 19947 5355
rect 19978 5352 19984 5364
rect 19935 5324 19984 5352
rect 19935 5321 19947 5324
rect 19889 5315 19947 5321
rect 19978 5312 19984 5324
rect 20036 5312 20042 5364
rect 14190 5241 14248 5247
rect 15562 5244 15568 5296
rect 15620 5284 15626 5296
rect 15948 5284 15976 5312
rect 16574 5284 16580 5296
rect 15620 5256 15792 5284
rect 15948 5256 16580 5284
rect 15620 5244 15626 5256
rect 7929 5219 7987 5225
rect 7929 5185 7941 5219
rect 7975 5216 7987 5219
rect 8018 5216 8024 5228
rect 7975 5188 8024 5216
rect 7975 5185 7987 5188
rect 7929 5179 7987 5185
rect 8018 5176 8024 5188
rect 8076 5176 8082 5228
rect 8294 5176 8300 5228
rect 8352 5176 8358 5228
rect 11330 5176 11336 5228
rect 11388 5216 11394 5228
rect 11609 5219 11667 5225
rect 11609 5216 11621 5219
rect 11388 5188 11621 5216
rect 11388 5176 11394 5188
rect 11609 5185 11621 5188
rect 11655 5185 11667 5219
rect 11609 5179 11667 5185
rect 11698 5176 11704 5228
rect 11756 5176 11762 5228
rect 11793 5219 11851 5225
rect 11793 5185 11805 5219
rect 11839 5216 11851 5219
rect 12618 5216 12624 5228
rect 11839 5188 12624 5216
rect 11839 5185 11851 5188
rect 11793 5179 11851 5185
rect 12618 5176 12624 5188
rect 12676 5216 12682 5228
rect 12897 5219 12955 5225
rect 12897 5216 12909 5219
rect 12676 5188 12909 5216
rect 12676 5176 12682 5188
rect 12897 5185 12909 5188
rect 12943 5185 12955 5219
rect 12897 5179 12955 5185
rect 13078 5176 13084 5228
rect 13136 5176 13142 5228
rect 13357 5219 13415 5225
rect 13357 5185 13369 5219
rect 13403 5185 13415 5219
rect 13357 5179 13415 5185
rect 2924 5120 5212 5148
rect 2924 5108 2930 5120
rect 11882 5108 11888 5160
rect 11940 5108 11946 5160
rect 12986 5108 12992 5160
rect 13044 5148 13050 5160
rect 13372 5148 13400 5179
rect 13630 5176 13636 5228
rect 13688 5216 13694 5228
rect 13817 5219 13875 5225
rect 13817 5216 13829 5219
rect 13688 5188 13829 5216
rect 13688 5176 13694 5188
rect 13817 5185 13829 5188
rect 13863 5185 13875 5219
rect 13817 5179 13875 5185
rect 14093 5219 14151 5225
rect 14093 5185 14105 5219
rect 14139 5185 14151 5219
rect 14190 5207 14202 5241
rect 14236 5207 14248 5241
rect 14190 5201 14248 5207
rect 14093 5179 14151 5185
rect 14108 5148 14136 5179
rect 15654 5176 15660 5228
rect 15712 5176 15718 5228
rect 15764 5225 15792 5256
rect 16574 5244 16580 5256
rect 16632 5244 16638 5296
rect 15750 5219 15808 5225
rect 15750 5185 15762 5219
rect 15796 5185 15808 5219
rect 15750 5179 15808 5185
rect 20073 5219 20131 5225
rect 20073 5185 20085 5219
rect 20119 5216 20131 5219
rect 21542 5216 21548 5228
rect 20119 5188 21548 5216
rect 20119 5185 20131 5188
rect 20073 5179 20131 5185
rect 21542 5176 21548 5188
rect 21600 5176 21606 5228
rect 14918 5148 14924 5160
rect 13044 5120 14924 5148
rect 13044 5108 13050 5120
rect 14918 5108 14924 5120
rect 14976 5108 14982 5160
rect 11238 5040 11244 5092
rect 11296 5080 11302 5092
rect 13173 5083 13231 5089
rect 13173 5080 13185 5083
rect 11296 5052 13185 5080
rect 11296 5040 11302 5052
rect 13173 5049 13185 5052
rect 13219 5080 13231 5083
rect 13630 5080 13636 5092
rect 13219 5052 13636 5080
rect 13219 5049 13231 5052
rect 13173 5043 13231 5049
rect 13630 5040 13636 5052
rect 13688 5040 13694 5092
rect 13725 5083 13783 5089
rect 13725 5049 13737 5083
rect 13771 5080 13783 5083
rect 13906 5080 13912 5092
rect 13771 5052 13912 5080
rect 13771 5049 13783 5052
rect 13725 5043 13783 5049
rect 13906 5040 13912 5052
rect 13964 5040 13970 5092
rect 6641 5015 6699 5021
rect 6641 4981 6653 5015
rect 6687 5012 6699 5015
rect 7098 5012 7104 5024
rect 6687 4984 7104 5012
rect 6687 4981 6699 4984
rect 6641 4975 6699 4981
rect 7098 4972 7104 4984
rect 7156 4972 7162 5024
rect 12069 5015 12127 5021
rect 12069 4981 12081 5015
rect 12115 5012 12127 5015
rect 12894 5012 12900 5024
rect 12115 4984 12900 5012
rect 12115 4981 12127 4984
rect 12069 4975 12127 4981
rect 12894 4972 12900 4984
rect 12952 4972 12958 5024
rect 12989 5015 13047 5021
rect 12989 4981 13001 5015
rect 13035 5012 13047 5015
rect 13354 5012 13360 5024
rect 13035 4984 13360 5012
rect 13035 4981 13047 4984
rect 12989 4975 13047 4981
rect 13354 4972 13360 4984
rect 13412 4972 13418 5024
rect 13814 4972 13820 5024
rect 13872 4972 13878 5024
rect 1104 4922 25208 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 25208 4922
rect 1104 4848 25208 4870
rect 12989 4675 13047 4681
rect 12989 4641 13001 4675
rect 13035 4672 13047 4675
rect 13262 4672 13268 4684
rect 13035 4644 13268 4672
rect 13035 4641 13047 4644
rect 12989 4635 13047 4641
rect 13262 4632 13268 4644
rect 13320 4632 13326 4684
rect 12894 4564 12900 4616
rect 12952 4564 12958 4616
rect 13265 4471 13323 4477
rect 13265 4437 13277 4471
rect 13311 4468 13323 4471
rect 15102 4468 15108 4480
rect 13311 4440 15108 4468
rect 13311 4437 13323 4440
rect 13265 4431 13323 4437
rect 15102 4428 15108 4440
rect 15160 4428 15166 4480
rect 1104 4378 25208 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 25208 4378
rect 1104 4304 25208 4326
rect 15286 4224 15292 4276
rect 15344 4224 15350 4276
rect 15102 4156 15108 4208
rect 15160 4196 15166 4208
rect 15381 4199 15439 4205
rect 15381 4196 15393 4199
rect 15160 4168 15393 4196
rect 15160 4156 15166 4168
rect 15381 4165 15393 4168
rect 15427 4165 15439 4199
rect 15381 4159 15439 4165
rect 15488 4168 15700 4196
rect 13354 4088 13360 4140
rect 13412 4088 13418 4140
rect 13541 4131 13599 4137
rect 13541 4097 13553 4131
rect 13587 4128 13599 4131
rect 13722 4128 13728 4140
rect 13587 4100 13728 4128
rect 13587 4097 13599 4100
rect 13541 4091 13599 4097
rect 13722 4088 13728 4100
rect 13780 4088 13786 4140
rect 13817 4131 13875 4137
rect 13817 4097 13829 4131
rect 13863 4128 13875 4131
rect 13906 4128 13912 4140
rect 13863 4100 13912 4128
rect 13863 4097 13875 4100
rect 13817 4091 13875 4097
rect 13906 4088 13912 4100
rect 13964 4088 13970 4140
rect 14093 4131 14151 4137
rect 14093 4097 14105 4131
rect 14139 4097 14151 4131
rect 14093 4091 14151 4097
rect 13372 4060 13400 4088
rect 14108 4060 14136 4091
rect 14918 4088 14924 4140
rect 14976 4128 14982 4140
rect 15488 4128 15516 4168
rect 14976 4100 15516 4128
rect 15565 4131 15623 4137
rect 14976 4088 14982 4100
rect 15565 4097 15577 4131
rect 15611 4097 15623 4131
rect 15565 4091 15623 4097
rect 13372 4032 14136 4060
rect 14182 4020 14188 4072
rect 14240 4020 14246 4072
rect 14829 4063 14887 4069
rect 14829 4029 14841 4063
rect 14875 4029 14887 4063
rect 14829 4023 14887 4029
rect 13541 3995 13599 4001
rect 13541 3961 13553 3995
rect 13587 3992 13599 3995
rect 14844 3992 14872 4023
rect 13587 3964 14872 3992
rect 13587 3961 13599 3964
rect 13541 3955 13599 3961
rect 14369 3927 14427 3933
rect 14369 3893 14381 3927
rect 14415 3924 14427 3927
rect 15194 3924 15200 3936
rect 14415 3896 15200 3924
rect 14415 3893 14427 3896
rect 14369 3887 14427 3893
rect 15194 3884 15200 3896
rect 15252 3924 15258 3936
rect 15580 3924 15608 4091
rect 15672 4060 15700 4168
rect 15749 4131 15807 4137
rect 15749 4097 15761 4131
rect 15795 4128 15807 4131
rect 16025 4131 16083 4137
rect 16025 4128 16037 4131
rect 15795 4100 16037 4128
rect 15795 4097 15807 4100
rect 15749 4091 15807 4097
rect 16025 4097 16037 4100
rect 16071 4097 16083 4131
rect 16025 4091 16083 4097
rect 16209 4131 16267 4137
rect 16209 4097 16221 4131
rect 16255 4128 16267 4131
rect 18690 4128 18696 4140
rect 16255 4100 18696 4128
rect 16255 4097 16267 4100
rect 16209 4091 16267 4097
rect 18690 4088 18696 4100
rect 18748 4088 18754 4140
rect 15841 4063 15899 4069
rect 15841 4060 15853 4063
rect 15672 4032 15853 4060
rect 15841 4029 15853 4032
rect 15887 4029 15899 4063
rect 15841 4023 15899 4029
rect 15252 3896 15608 3924
rect 15252 3884 15258 3896
rect 1104 3834 25208 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 25208 3834
rect 1104 3760 25208 3782
rect 14093 3723 14151 3729
rect 14093 3689 14105 3723
rect 14139 3720 14151 3723
rect 14182 3720 14188 3732
rect 14139 3692 14188 3720
rect 14139 3689 14151 3692
rect 14093 3683 14151 3689
rect 14182 3680 14188 3692
rect 14240 3680 14246 3732
rect 14829 3723 14887 3729
rect 14829 3689 14841 3723
rect 14875 3720 14887 3723
rect 14918 3720 14924 3732
rect 14875 3692 14924 3720
rect 14875 3689 14887 3692
rect 14829 3683 14887 3689
rect 14918 3680 14924 3692
rect 14976 3680 14982 3732
rect 24670 3680 24676 3732
rect 24728 3680 24734 3732
rect 13906 3544 13912 3596
rect 13964 3584 13970 3596
rect 15102 3584 15108 3596
rect 13964 3556 14320 3584
rect 13964 3544 13970 3556
rect 13814 3476 13820 3528
rect 13872 3516 13878 3528
rect 14292 3525 14320 3556
rect 14752 3556 15108 3584
rect 14752 3525 14780 3556
rect 15102 3544 15108 3556
rect 15160 3544 15166 3596
rect 14093 3519 14151 3525
rect 14093 3516 14105 3519
rect 13872 3488 14105 3516
rect 13872 3476 13878 3488
rect 14093 3485 14105 3488
rect 14139 3485 14151 3519
rect 14093 3479 14151 3485
rect 14277 3519 14335 3525
rect 14277 3485 14289 3519
rect 14323 3485 14335 3519
rect 14277 3479 14335 3485
rect 14737 3519 14795 3525
rect 14737 3485 14749 3519
rect 14783 3485 14795 3519
rect 14737 3479 14795 3485
rect 14921 3519 14979 3525
rect 14921 3485 14933 3519
rect 14967 3516 14979 3519
rect 15194 3516 15200 3528
rect 14967 3488 15200 3516
rect 14967 3485 14979 3488
rect 14921 3479 14979 3485
rect 15194 3476 15200 3488
rect 15252 3476 15258 3528
rect 24854 3476 24860 3528
rect 24912 3476 24918 3528
rect 1104 3290 25208 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 25208 3290
rect 1104 3216 25208 3238
rect 1104 2746 25208 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 25208 2746
rect 1104 2672 25208 2694
rect 1104 2202 25208 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 25208 2202
rect 1104 2128 25208 2150
<< via1 >>
rect 4874 26086 4926 26138
rect 4938 26086 4990 26138
rect 5002 26086 5054 26138
rect 5066 26086 5118 26138
rect 5130 26086 5182 26138
rect 9220 25959 9272 25968
rect 9220 25925 9229 25959
rect 9229 25925 9263 25959
rect 9263 25925 9272 25959
rect 9220 25916 9272 25925
rect 9864 25959 9916 25968
rect 9864 25925 9873 25959
rect 9873 25925 9907 25959
rect 9907 25925 9916 25959
rect 9864 25916 9916 25925
rect 10508 25959 10560 25968
rect 10508 25925 10517 25959
rect 10517 25925 10551 25959
rect 10551 25925 10560 25959
rect 10508 25916 10560 25925
rect 12348 25916 12400 25968
rect 13728 25959 13780 25968
rect 13728 25925 13737 25959
rect 13737 25925 13771 25959
rect 13771 25925 13780 25959
rect 13728 25916 13780 25925
rect 14372 25959 14424 25968
rect 14372 25925 14381 25959
rect 14381 25925 14415 25959
rect 14415 25925 14424 25959
rect 14372 25916 14424 25925
rect 15016 25959 15068 25968
rect 15016 25925 15025 25959
rect 15025 25925 15059 25959
rect 15059 25925 15068 25959
rect 15016 25916 15068 25925
rect 17592 25959 17644 25968
rect 17592 25925 17601 25959
rect 17601 25925 17635 25959
rect 17635 25925 17644 25959
rect 17592 25916 17644 25925
rect 18236 25959 18288 25968
rect 18236 25925 18245 25959
rect 18245 25925 18279 25959
rect 18279 25925 18288 25959
rect 18236 25916 18288 25925
rect 4712 25848 4764 25900
rect 10876 25848 10928 25900
rect 11704 25891 11756 25900
rect 11704 25857 11713 25891
rect 11713 25857 11747 25891
rect 11747 25857 11756 25891
rect 11704 25848 11756 25857
rect 12992 25891 13044 25900
rect 12992 25857 13001 25891
rect 13001 25857 13035 25891
rect 13035 25857 13044 25891
rect 12992 25848 13044 25857
rect 15568 25891 15620 25900
rect 15568 25857 15577 25891
rect 15577 25857 15611 25891
rect 15611 25857 15620 25891
rect 15568 25848 15620 25857
rect 16212 25891 16264 25900
rect 16212 25857 16221 25891
rect 16221 25857 16255 25891
rect 16255 25857 16264 25891
rect 16212 25848 16264 25857
rect 4620 25780 4672 25832
rect 10600 25780 10652 25832
rect 17500 25780 17552 25832
rect 12808 25712 12860 25764
rect 13912 25755 13964 25764
rect 13912 25721 13921 25755
rect 13921 25721 13955 25755
rect 13955 25721 13964 25755
rect 13912 25712 13964 25721
rect 14648 25712 14700 25764
rect 17776 25712 17828 25764
rect 18420 25755 18472 25764
rect 18420 25721 18429 25755
rect 18429 25721 18463 25755
rect 18463 25721 18472 25755
rect 18420 25712 18472 25721
rect 2044 25644 2096 25696
rect 4804 25644 4856 25696
rect 9312 25687 9364 25696
rect 9312 25653 9321 25687
rect 9321 25653 9355 25687
rect 9355 25653 9364 25687
rect 9312 25644 9364 25653
rect 10140 25644 10192 25696
rect 11060 25687 11112 25696
rect 11060 25653 11069 25687
rect 11069 25653 11103 25687
rect 11103 25653 11112 25687
rect 11060 25644 11112 25653
rect 11888 25687 11940 25696
rect 11888 25653 11897 25687
rect 11897 25653 11931 25687
rect 11931 25653 11940 25687
rect 11888 25644 11940 25653
rect 13820 25644 13872 25696
rect 16948 25644 17000 25696
rect 17408 25644 17460 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 4620 25440 4672 25492
rect 4712 25483 4764 25492
rect 4712 25449 4721 25483
rect 4721 25449 4755 25483
rect 4755 25449 4764 25483
rect 4712 25440 4764 25449
rect 2044 25347 2096 25356
rect 2044 25313 2053 25347
rect 2053 25313 2087 25347
rect 2087 25313 2096 25347
rect 2044 25304 2096 25313
rect 3700 25304 3752 25356
rect 1400 25236 1452 25288
rect 4160 25236 4212 25288
rect 4712 25279 4764 25288
rect 4712 25245 4721 25279
rect 4721 25245 4755 25279
rect 4755 25245 4764 25279
rect 4712 25236 4764 25245
rect 4804 25279 4856 25288
rect 4804 25245 4813 25279
rect 4813 25245 4847 25279
rect 4847 25245 4856 25279
rect 4804 25236 4856 25245
rect 6000 25279 6052 25288
rect 6000 25245 6009 25279
rect 6009 25245 6043 25279
rect 6043 25245 6052 25279
rect 6000 25236 6052 25245
rect 3056 25168 3108 25220
rect 5356 25168 5408 25220
rect 7380 25168 7432 25220
rect 12072 25304 12124 25356
rect 8484 25236 8536 25288
rect 11060 25279 11112 25288
rect 11060 25245 11069 25279
rect 11069 25245 11103 25279
rect 11103 25245 11112 25279
rect 11060 25236 11112 25245
rect 12992 25279 13044 25288
rect 12992 25245 13001 25279
rect 13001 25245 13035 25279
rect 13035 25245 13044 25279
rect 12992 25236 13044 25245
rect 13360 25347 13412 25356
rect 13360 25313 13369 25347
rect 13369 25313 13403 25347
rect 13403 25313 13412 25347
rect 13360 25304 13412 25313
rect 19524 25304 19576 25356
rect 15292 25236 15344 25288
rect 15476 25236 15528 25288
rect 24860 25279 24912 25288
rect 24860 25245 24869 25279
rect 24869 25245 24903 25279
rect 24903 25245 24912 25279
rect 24860 25236 24912 25245
rect 4804 25100 4856 25152
rect 5264 25100 5316 25152
rect 7564 25100 7616 25152
rect 8392 25100 8444 25152
rect 8576 25100 8628 25152
rect 9220 25211 9272 25220
rect 9220 25177 9229 25211
rect 9229 25177 9263 25211
rect 9263 25177 9272 25211
rect 9220 25168 9272 25177
rect 9956 25168 10008 25220
rect 11336 25168 11388 25220
rect 12716 25211 12768 25220
rect 12716 25177 12725 25211
rect 12725 25177 12759 25211
rect 12759 25177 12768 25211
rect 12716 25168 12768 25177
rect 15844 25211 15896 25220
rect 15844 25177 15853 25211
rect 15853 25177 15887 25211
rect 15887 25177 15896 25211
rect 15844 25168 15896 25177
rect 16856 25168 16908 25220
rect 19432 25168 19484 25220
rect 21088 25168 21140 25220
rect 10508 25100 10560 25152
rect 10968 25143 11020 25152
rect 10968 25109 10977 25143
rect 10977 25109 11011 25143
rect 11011 25109 11020 25143
rect 10968 25100 11020 25109
rect 11244 25143 11296 25152
rect 11244 25109 11253 25143
rect 11253 25109 11287 25143
rect 11287 25109 11296 25143
rect 11244 25100 11296 25109
rect 13544 25100 13596 25152
rect 17592 25100 17644 25152
rect 20996 25143 21048 25152
rect 20996 25109 21005 25143
rect 21005 25109 21039 25143
rect 21039 25109 21048 25143
rect 20996 25100 21048 25109
rect 4874 24998 4926 25050
rect 4938 24998 4990 25050
rect 5002 24998 5054 25050
rect 5066 24998 5118 25050
rect 5130 24998 5182 25050
rect 3056 24896 3108 24948
rect 6000 24896 6052 24948
rect 9220 24896 9272 24948
rect 14740 24896 14792 24948
rect 8760 24828 8812 24880
rect 8484 24803 8536 24812
rect 8484 24769 8493 24803
rect 8493 24769 8527 24803
rect 8527 24769 8536 24803
rect 8484 24760 8536 24769
rect 8668 24760 8720 24812
rect 9220 24803 9272 24812
rect 9220 24769 9229 24803
rect 9229 24769 9263 24803
rect 9263 24769 9272 24803
rect 9220 24760 9272 24769
rect 9404 24803 9456 24812
rect 9404 24769 9413 24803
rect 9413 24769 9447 24803
rect 9447 24769 9456 24803
rect 9404 24760 9456 24769
rect 1400 24692 1452 24744
rect 1768 24735 1820 24744
rect 1768 24701 1777 24735
rect 1777 24701 1811 24735
rect 1811 24701 1820 24735
rect 1768 24692 1820 24701
rect 3884 24735 3936 24744
rect 3884 24701 3893 24735
rect 3893 24701 3927 24735
rect 3927 24701 3936 24735
rect 3884 24692 3936 24701
rect 4528 24692 4580 24744
rect 8208 24735 8260 24744
rect 8208 24701 8217 24735
rect 8217 24701 8251 24735
rect 8251 24701 8260 24735
rect 8208 24692 8260 24701
rect 10784 24760 10836 24812
rect 12532 24760 12584 24812
rect 14464 24760 14516 24812
rect 15844 24896 15896 24948
rect 19892 24896 19944 24948
rect 17592 24828 17644 24880
rect 12716 24735 12768 24744
rect 12716 24701 12725 24735
rect 12725 24701 12759 24735
rect 12759 24701 12768 24735
rect 12716 24692 12768 24701
rect 12992 24692 13044 24744
rect 8760 24624 8812 24676
rect 9956 24624 10008 24676
rect 3332 24599 3384 24608
rect 3332 24565 3341 24599
rect 3341 24565 3375 24599
rect 3375 24565 3384 24599
rect 3332 24556 3384 24565
rect 7196 24556 7248 24608
rect 8392 24556 8444 24608
rect 8484 24556 8536 24608
rect 9036 24556 9088 24608
rect 10232 24556 10284 24608
rect 12900 24599 12952 24608
rect 12900 24565 12909 24599
rect 12909 24565 12943 24599
rect 12943 24565 12952 24599
rect 12900 24556 12952 24565
rect 13360 24735 13412 24744
rect 13360 24701 13369 24735
rect 13369 24701 13403 24735
rect 13403 24701 13412 24735
rect 13360 24692 13412 24701
rect 13728 24692 13780 24744
rect 14924 24735 14976 24744
rect 14924 24701 14933 24735
rect 14933 24701 14967 24735
rect 14967 24701 14976 24735
rect 14924 24692 14976 24701
rect 15476 24624 15528 24676
rect 15016 24599 15068 24608
rect 15016 24565 15025 24599
rect 15025 24565 15059 24599
rect 15059 24565 15068 24599
rect 15016 24556 15068 24565
rect 16028 24803 16080 24812
rect 16028 24769 16037 24803
rect 16037 24769 16071 24803
rect 16071 24769 16080 24803
rect 16028 24760 16080 24769
rect 16120 24735 16172 24744
rect 16120 24701 16129 24735
rect 16129 24701 16163 24735
rect 16163 24701 16172 24735
rect 16120 24692 16172 24701
rect 17132 24803 17184 24812
rect 17132 24769 17141 24803
rect 17141 24769 17175 24803
rect 17175 24769 17184 24803
rect 17132 24760 17184 24769
rect 17224 24803 17276 24812
rect 17224 24769 17233 24803
rect 17233 24769 17267 24803
rect 17267 24769 17276 24803
rect 17224 24760 17276 24769
rect 17868 24828 17920 24880
rect 17316 24692 17368 24744
rect 17132 24624 17184 24676
rect 17776 24803 17828 24812
rect 17776 24769 17785 24803
rect 17785 24769 17819 24803
rect 17819 24769 17828 24803
rect 17776 24760 17828 24769
rect 17500 24735 17552 24744
rect 17500 24701 17509 24735
rect 17509 24701 17543 24735
rect 17543 24701 17552 24735
rect 17500 24692 17552 24701
rect 17684 24692 17736 24744
rect 18144 24760 18196 24812
rect 21088 24828 21140 24880
rect 21548 24828 21600 24880
rect 19432 24760 19484 24812
rect 21364 24760 21416 24812
rect 22376 24760 22428 24812
rect 22652 24803 22704 24812
rect 22652 24769 22661 24803
rect 22661 24769 22695 24803
rect 22695 24769 22704 24803
rect 22652 24760 22704 24769
rect 19340 24692 19392 24744
rect 19524 24735 19576 24744
rect 19524 24701 19533 24735
rect 19533 24701 19567 24735
rect 19567 24701 19576 24735
rect 19524 24692 19576 24701
rect 19800 24735 19852 24744
rect 19800 24701 19809 24735
rect 19809 24701 19843 24735
rect 19843 24701 19852 24735
rect 19800 24692 19852 24701
rect 19432 24556 19484 24608
rect 20812 24624 20864 24676
rect 20536 24556 20588 24608
rect 21180 24556 21232 24608
rect 23020 24556 23072 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 3884 24352 3936 24404
rect 4252 24395 4304 24404
rect 4252 24361 4261 24395
rect 4261 24361 4295 24395
rect 4295 24361 4304 24395
rect 4252 24352 4304 24361
rect 4344 24352 4396 24404
rect 4804 24352 4856 24404
rect 7196 24352 7248 24404
rect 8300 24352 8352 24404
rect 8392 24395 8444 24404
rect 8392 24361 8401 24395
rect 8401 24361 8435 24395
rect 8435 24361 8444 24395
rect 8392 24352 8444 24361
rect 8576 24352 8628 24404
rect 10508 24352 10560 24404
rect 11152 24352 11204 24404
rect 12716 24352 12768 24404
rect 13360 24352 13412 24404
rect 16120 24352 16172 24404
rect 17224 24395 17276 24404
rect 17224 24361 17233 24395
rect 17233 24361 17267 24395
rect 17267 24361 17276 24395
rect 17224 24352 17276 24361
rect 17316 24352 17368 24404
rect 1768 24284 1820 24336
rect 4620 24327 4672 24336
rect 4620 24293 4629 24327
rect 4629 24293 4663 24327
rect 4663 24293 4672 24327
rect 4620 24284 4672 24293
rect 3700 24216 3752 24268
rect 8116 24284 8168 24336
rect 9220 24284 9272 24336
rect 10784 24327 10836 24336
rect 10784 24293 10793 24327
rect 10793 24293 10827 24327
rect 10827 24293 10836 24327
rect 10784 24284 10836 24293
rect 3240 24191 3292 24200
rect 3240 24157 3249 24191
rect 3249 24157 3283 24191
rect 3283 24157 3292 24191
rect 3240 24148 3292 24157
rect 2044 24123 2096 24132
rect 2044 24089 2053 24123
rect 2053 24089 2087 24123
rect 2087 24089 2096 24123
rect 2044 24080 2096 24089
rect 3424 24191 3476 24200
rect 3424 24157 3433 24191
rect 3433 24157 3467 24191
rect 3467 24157 3476 24191
rect 3424 24148 3476 24157
rect 3608 24191 3660 24200
rect 3608 24157 3617 24191
rect 3617 24157 3651 24191
rect 3651 24157 3660 24191
rect 3608 24148 3660 24157
rect 3884 24191 3936 24200
rect 3884 24157 3893 24191
rect 3893 24157 3927 24191
rect 3927 24157 3936 24191
rect 3884 24148 3936 24157
rect 4160 24148 4212 24200
rect 2780 24055 2832 24064
rect 2780 24021 2789 24055
rect 2789 24021 2823 24055
rect 2823 24021 2832 24055
rect 2780 24012 2832 24021
rect 2872 24055 2924 24064
rect 2872 24021 2881 24055
rect 2881 24021 2915 24055
rect 2915 24021 2924 24055
rect 2872 24012 2924 24021
rect 3608 24012 3660 24064
rect 4068 24012 4120 24064
rect 4804 24191 4856 24200
rect 4804 24157 4813 24191
rect 4813 24157 4847 24191
rect 4847 24157 4856 24191
rect 4804 24148 4856 24157
rect 5264 24148 5316 24200
rect 6184 24080 6236 24132
rect 4528 24055 4580 24064
rect 4528 24021 4537 24055
rect 4537 24021 4571 24055
rect 4571 24021 4580 24055
rect 4528 24012 4580 24021
rect 4712 24012 4764 24064
rect 5264 24012 5316 24064
rect 6920 24012 6972 24064
rect 7472 24080 7524 24132
rect 7564 24123 7616 24132
rect 7564 24089 7573 24123
rect 7573 24089 7607 24123
rect 7607 24089 7616 24123
rect 7564 24080 7616 24089
rect 7380 24055 7432 24064
rect 7380 24021 7407 24055
rect 7407 24021 7432 24055
rect 7380 24012 7432 24021
rect 8208 24216 8260 24268
rect 8668 24216 8720 24268
rect 17040 24284 17092 24336
rect 18880 24395 18932 24404
rect 18880 24361 18889 24395
rect 18889 24361 18923 24395
rect 18923 24361 18932 24395
rect 18880 24352 18932 24361
rect 7840 24191 7892 24200
rect 7840 24157 7849 24191
rect 7849 24157 7883 24191
rect 7883 24157 7892 24191
rect 7840 24148 7892 24157
rect 8392 24148 8444 24200
rect 10416 24191 10468 24200
rect 10416 24157 10425 24191
rect 10425 24157 10459 24191
rect 10459 24157 10468 24191
rect 10416 24148 10468 24157
rect 10508 24191 10560 24200
rect 10508 24157 10517 24191
rect 10517 24157 10551 24191
rect 10551 24157 10560 24191
rect 10508 24148 10560 24157
rect 10784 24148 10836 24200
rect 11152 24191 11204 24200
rect 11152 24157 11162 24191
rect 11162 24157 11196 24191
rect 11196 24157 11204 24191
rect 11152 24148 11204 24157
rect 12808 24216 12860 24268
rect 12900 24216 12952 24268
rect 12624 24191 12676 24200
rect 12624 24157 12633 24191
rect 12633 24157 12667 24191
rect 12667 24157 12676 24191
rect 12624 24148 12676 24157
rect 13268 24191 13320 24200
rect 13268 24157 13277 24191
rect 13277 24157 13311 24191
rect 13311 24157 13320 24191
rect 13268 24148 13320 24157
rect 13360 24191 13412 24200
rect 13360 24157 13369 24191
rect 13369 24157 13403 24191
rect 13403 24157 13412 24191
rect 13360 24148 13412 24157
rect 13544 24191 13596 24200
rect 13544 24157 13553 24191
rect 13553 24157 13587 24191
rect 13587 24157 13596 24191
rect 13544 24148 13596 24157
rect 14464 24216 14516 24268
rect 15384 24191 15436 24200
rect 15384 24157 15393 24191
rect 15393 24157 15427 24191
rect 15427 24157 15436 24191
rect 15384 24148 15436 24157
rect 16856 24216 16908 24268
rect 17132 24148 17184 24200
rect 11060 24012 11112 24064
rect 11796 24012 11848 24064
rect 12716 24012 12768 24064
rect 15016 24080 15068 24132
rect 17592 24191 17644 24200
rect 17592 24157 17601 24191
rect 17601 24157 17635 24191
rect 17635 24157 17644 24191
rect 17592 24148 17644 24157
rect 17684 24080 17736 24132
rect 13728 24012 13780 24064
rect 16580 24012 16632 24064
rect 17776 24012 17828 24064
rect 19156 24284 19208 24336
rect 19800 24352 19852 24404
rect 21088 24395 21140 24404
rect 21088 24361 21097 24395
rect 21097 24361 21131 24395
rect 21131 24361 21140 24395
rect 21088 24352 21140 24361
rect 22376 24352 22428 24404
rect 19248 24259 19300 24268
rect 19248 24225 19257 24259
rect 19257 24225 19291 24259
rect 19291 24225 19300 24259
rect 19248 24216 19300 24225
rect 18972 24148 19024 24200
rect 19892 24216 19944 24268
rect 20996 24284 21048 24336
rect 17960 24080 18012 24132
rect 19708 24191 19760 24200
rect 19708 24157 19717 24191
rect 19717 24157 19751 24191
rect 19751 24157 19760 24191
rect 19708 24148 19760 24157
rect 20076 24148 20128 24200
rect 20628 24216 20680 24268
rect 22928 24216 22980 24268
rect 20904 24191 20956 24200
rect 20904 24157 20913 24191
rect 20913 24157 20947 24191
rect 20947 24157 20956 24191
rect 20904 24148 20956 24157
rect 21272 24148 21324 24200
rect 21548 24148 21600 24200
rect 18604 24012 18656 24064
rect 23020 24123 23072 24132
rect 23020 24089 23029 24123
rect 23029 24089 23063 24123
rect 23063 24089 23072 24123
rect 23020 24080 23072 24089
rect 19616 24012 19668 24064
rect 19892 24012 19944 24064
rect 20168 24012 20220 24064
rect 21088 24012 21140 24064
rect 22744 24012 22796 24064
rect 4874 23910 4926 23962
rect 4938 23910 4990 23962
rect 5002 23910 5054 23962
rect 5066 23910 5118 23962
rect 5130 23910 5182 23962
rect 1768 23808 1820 23860
rect 3240 23808 3292 23860
rect 3332 23740 3384 23792
rect 7196 23808 7248 23860
rect 2872 23672 2924 23724
rect 4528 23740 4580 23792
rect 3700 23715 3752 23724
rect 3700 23681 3709 23715
rect 3709 23681 3743 23715
rect 3743 23681 3752 23715
rect 3700 23672 3752 23681
rect 3884 23715 3936 23724
rect 3884 23681 3893 23715
rect 3893 23681 3927 23715
rect 3927 23681 3936 23715
rect 3884 23672 3936 23681
rect 4160 23672 4212 23724
rect 3424 23647 3476 23656
rect 3424 23613 3433 23647
rect 3433 23613 3467 23647
rect 3467 23613 3476 23647
rect 3424 23604 3476 23613
rect 4252 23604 4304 23656
rect 4620 23604 4672 23656
rect 5172 23672 5224 23724
rect 6920 23783 6972 23792
rect 6920 23749 6929 23783
rect 6929 23749 6963 23783
rect 6963 23749 6972 23783
rect 6920 23740 6972 23749
rect 5264 23604 5316 23656
rect 6000 23672 6052 23724
rect 7104 23715 7156 23724
rect 7104 23681 7113 23715
rect 7113 23681 7147 23715
rect 7147 23681 7156 23715
rect 7104 23672 7156 23681
rect 11244 23851 11296 23860
rect 11244 23817 11253 23851
rect 11253 23817 11287 23851
rect 11287 23817 11296 23851
rect 11244 23808 11296 23817
rect 12164 23808 12216 23860
rect 12624 23808 12676 23860
rect 12900 23808 12952 23860
rect 15752 23808 15804 23860
rect 16580 23808 16632 23860
rect 19248 23808 19300 23860
rect 12992 23740 13044 23792
rect 13360 23740 13412 23792
rect 15108 23740 15160 23792
rect 8392 23715 8444 23724
rect 2412 23468 2464 23520
rect 4804 23536 4856 23588
rect 4344 23468 4396 23520
rect 4712 23468 4764 23520
rect 6092 23604 6144 23656
rect 7380 23604 7432 23656
rect 8392 23681 8401 23715
rect 8401 23681 8435 23715
rect 8435 23681 8444 23715
rect 8392 23672 8444 23681
rect 11060 23715 11112 23724
rect 11060 23681 11069 23715
rect 11069 23681 11103 23715
rect 11103 23681 11112 23715
rect 11060 23672 11112 23681
rect 7656 23604 7708 23656
rect 11796 23715 11848 23724
rect 11796 23681 11805 23715
rect 11805 23681 11839 23715
rect 11839 23681 11848 23715
rect 11796 23672 11848 23681
rect 12440 23672 12492 23724
rect 12900 23672 12952 23724
rect 13084 23715 13136 23724
rect 13084 23681 13093 23715
rect 13093 23681 13127 23715
rect 13127 23681 13136 23715
rect 13084 23672 13136 23681
rect 17776 23740 17828 23792
rect 17868 23783 17920 23792
rect 17868 23749 17877 23783
rect 17877 23749 17911 23783
rect 17911 23749 17920 23783
rect 17868 23740 17920 23749
rect 19156 23783 19208 23792
rect 19156 23749 19165 23783
rect 19165 23749 19199 23783
rect 19199 23749 19208 23783
rect 19156 23740 19208 23749
rect 16948 23715 17000 23724
rect 16948 23681 16957 23715
rect 16957 23681 16991 23715
rect 16991 23681 17000 23715
rect 16948 23672 17000 23681
rect 19064 23672 19116 23724
rect 20812 23808 20864 23860
rect 21088 23808 21140 23860
rect 19616 23783 19668 23792
rect 19616 23749 19625 23783
rect 19625 23749 19659 23783
rect 19659 23749 19668 23783
rect 19616 23740 19668 23749
rect 19892 23783 19944 23792
rect 19892 23749 19901 23783
rect 19901 23749 19935 23783
rect 19935 23749 19944 23783
rect 19892 23740 19944 23749
rect 20168 23740 20220 23792
rect 20996 23740 21048 23792
rect 21364 23740 21416 23792
rect 22376 23808 22428 23860
rect 22652 23808 22704 23860
rect 19708 23672 19760 23724
rect 7840 23536 7892 23588
rect 8760 23579 8812 23588
rect 8760 23545 8769 23579
rect 8769 23545 8803 23579
rect 8803 23545 8812 23579
rect 8760 23536 8812 23545
rect 11060 23536 11112 23588
rect 11152 23536 11204 23588
rect 12164 23579 12216 23588
rect 12164 23545 12173 23579
rect 12173 23545 12207 23579
rect 12207 23545 12216 23579
rect 12164 23536 12216 23545
rect 7288 23511 7340 23520
rect 7288 23477 7297 23511
rect 7297 23477 7331 23511
rect 7331 23477 7340 23511
rect 7288 23468 7340 23477
rect 7380 23511 7432 23520
rect 7380 23477 7389 23511
rect 7389 23477 7423 23511
rect 7423 23477 7432 23511
rect 7380 23468 7432 23477
rect 9036 23468 9088 23520
rect 10692 23511 10744 23520
rect 10692 23477 10701 23511
rect 10701 23477 10735 23511
rect 10735 23477 10744 23511
rect 10692 23468 10744 23477
rect 11244 23468 11296 23520
rect 14096 23604 14148 23656
rect 15292 23604 15344 23656
rect 18512 23604 18564 23656
rect 18880 23604 18932 23656
rect 19800 23604 19852 23656
rect 19892 23604 19944 23656
rect 20628 23604 20680 23656
rect 12348 23536 12400 23588
rect 12532 23468 12584 23520
rect 17684 23536 17736 23588
rect 17776 23536 17828 23588
rect 13268 23468 13320 23520
rect 15108 23468 15160 23520
rect 18420 23536 18472 23588
rect 18972 23536 19024 23588
rect 18328 23511 18380 23520
rect 18328 23477 18337 23511
rect 18337 23477 18371 23511
rect 18371 23477 18380 23511
rect 18328 23468 18380 23477
rect 19340 23468 19392 23520
rect 19800 23468 19852 23520
rect 21180 23672 21232 23724
rect 22284 23672 22336 23724
rect 20904 23604 20956 23656
rect 21088 23536 21140 23588
rect 22928 23604 22980 23656
rect 23204 23604 23256 23656
rect 20812 23511 20864 23520
rect 20812 23477 20821 23511
rect 20821 23477 20855 23511
rect 20855 23477 20864 23511
rect 20812 23468 20864 23477
rect 21272 23468 21324 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 3884 23264 3936 23316
rect 5172 23264 5224 23316
rect 7288 23264 7340 23316
rect 9588 23264 9640 23316
rect 2780 23196 2832 23248
rect 8392 23196 8444 23248
rect 7104 23128 7156 23180
rect 9772 23196 9824 23248
rect 11060 23307 11112 23316
rect 11060 23273 11069 23307
rect 11069 23273 11103 23307
rect 11103 23273 11112 23307
rect 11060 23264 11112 23273
rect 11244 23307 11296 23316
rect 11244 23273 11253 23307
rect 11253 23273 11287 23307
rect 11287 23273 11296 23307
rect 11244 23264 11296 23273
rect 12164 23264 12216 23316
rect 12532 23264 12584 23316
rect 14096 23264 14148 23316
rect 14924 23264 14976 23316
rect 15936 23264 15988 23316
rect 16672 23264 16724 23316
rect 16948 23264 17000 23316
rect 20812 23264 20864 23316
rect 10324 23128 10376 23180
rect 11060 23128 11112 23180
rect 1400 23103 1452 23112
rect 1400 23069 1409 23103
rect 1409 23069 1443 23103
rect 1443 23069 1452 23103
rect 1400 23060 1452 23069
rect 2780 23060 2832 23112
rect 4160 23103 4212 23112
rect 4160 23069 4169 23103
rect 4169 23069 4203 23103
rect 4203 23069 4212 23103
rect 4160 23060 4212 23069
rect 4620 23060 4672 23112
rect 7380 23103 7432 23112
rect 7380 23069 7389 23103
rect 7389 23069 7423 23103
rect 7423 23069 7432 23103
rect 7380 23060 7432 23069
rect 2964 22992 3016 23044
rect 3516 22992 3568 23044
rect 8668 23060 8720 23112
rect 10692 23060 10744 23112
rect 3608 22924 3660 22976
rect 8760 22992 8812 23044
rect 9312 22992 9364 23044
rect 9496 23035 9548 23044
rect 9496 23001 9505 23035
rect 9505 23001 9539 23035
rect 9539 23001 9548 23035
rect 9496 22992 9548 23001
rect 9680 22992 9732 23044
rect 8392 22924 8444 22976
rect 9128 22924 9180 22976
rect 9864 22967 9916 22976
rect 9864 22933 9873 22967
rect 9873 22933 9907 22967
rect 9907 22933 9916 22967
rect 9864 22924 9916 22933
rect 10048 22967 10100 22976
rect 10048 22933 10057 22967
rect 10057 22933 10091 22967
rect 10091 22933 10100 22967
rect 10048 22924 10100 22933
rect 10692 22924 10744 22976
rect 12808 23196 12860 23248
rect 12992 23239 13044 23248
rect 12992 23205 13001 23239
rect 13001 23205 13035 23239
rect 13035 23205 13044 23239
rect 12992 23196 13044 23205
rect 16764 23239 16816 23248
rect 16764 23205 16773 23239
rect 16773 23205 16807 23239
rect 16807 23205 16816 23239
rect 16764 23196 16816 23205
rect 11428 23060 11480 23112
rect 12440 23060 12492 23112
rect 12900 23060 12952 23112
rect 14188 23128 14240 23180
rect 14832 23128 14884 23180
rect 15476 23128 15528 23180
rect 18880 23128 18932 23180
rect 13544 23060 13596 23112
rect 14464 23060 14516 23112
rect 15936 23103 15988 23112
rect 15936 23069 15945 23103
rect 15945 23069 15979 23103
rect 15979 23069 15988 23103
rect 15936 23060 15988 23069
rect 17408 23103 17460 23112
rect 17408 23069 17417 23103
rect 17417 23069 17451 23103
rect 17451 23069 17460 23103
rect 17408 23060 17460 23069
rect 17684 23060 17736 23112
rect 17868 23060 17920 23112
rect 14280 22992 14332 23044
rect 13452 22924 13504 22976
rect 16488 23035 16540 23044
rect 16488 23001 16497 23035
rect 16497 23001 16531 23035
rect 16531 23001 16540 23035
rect 16488 22992 16540 23001
rect 17132 22924 17184 22976
rect 17960 22924 18012 22976
rect 4874 22822 4926 22874
rect 4938 22822 4990 22874
rect 5002 22822 5054 22874
rect 5066 22822 5118 22874
rect 5130 22822 5182 22874
rect 3884 22720 3936 22772
rect 7104 22720 7156 22772
rect 9496 22720 9548 22772
rect 2412 22652 2464 22704
rect 3148 22652 3200 22704
rect 6184 22652 6236 22704
rect 9680 22652 9732 22704
rect 10048 22720 10100 22772
rect 12532 22720 12584 22772
rect 12992 22720 13044 22772
rect 13176 22720 13228 22772
rect 13728 22720 13780 22772
rect 16028 22720 16080 22772
rect 16304 22720 16356 22772
rect 17408 22763 17460 22772
rect 17408 22729 17417 22763
rect 17417 22729 17451 22763
rect 17451 22729 17460 22763
rect 17408 22720 17460 22729
rect 23112 22720 23164 22772
rect 11888 22652 11940 22704
rect 12900 22652 12952 22704
rect 13820 22652 13872 22704
rect 8116 22627 8168 22636
rect 8116 22593 8125 22627
rect 8125 22593 8159 22627
rect 8159 22593 8168 22627
rect 8116 22584 8168 22593
rect 8760 22627 8812 22636
rect 8760 22593 8769 22627
rect 8769 22593 8803 22627
rect 8803 22593 8812 22627
rect 8760 22584 8812 22593
rect 8852 22627 8904 22636
rect 8852 22593 8861 22627
rect 8861 22593 8895 22627
rect 8895 22593 8904 22627
rect 8852 22584 8904 22593
rect 9036 22627 9088 22636
rect 9036 22593 9045 22627
rect 9045 22593 9079 22627
rect 9079 22593 9088 22627
rect 9036 22584 9088 22593
rect 9128 22627 9180 22636
rect 9128 22593 9137 22627
rect 9137 22593 9171 22627
rect 9171 22593 9180 22627
rect 9128 22584 9180 22593
rect 9404 22627 9456 22636
rect 9404 22593 9413 22627
rect 9413 22593 9447 22627
rect 9447 22593 9456 22627
rect 9404 22584 9456 22593
rect 9588 22627 9640 22636
rect 9588 22593 9597 22627
rect 9597 22593 9631 22627
rect 9631 22593 9640 22627
rect 9588 22584 9640 22593
rect 9772 22627 9824 22636
rect 9772 22593 9781 22627
rect 9781 22593 9815 22627
rect 9815 22593 9824 22627
rect 9772 22584 9824 22593
rect 1400 22516 1452 22568
rect 8392 22516 8444 22568
rect 9220 22516 9272 22568
rect 10692 22584 10744 22636
rect 12164 22627 12216 22636
rect 12164 22593 12173 22627
rect 12173 22593 12207 22627
rect 12207 22593 12216 22627
rect 12164 22584 12216 22593
rect 12256 22627 12308 22636
rect 12256 22593 12265 22627
rect 12265 22593 12299 22627
rect 12299 22593 12308 22627
rect 12256 22584 12308 22593
rect 12532 22584 12584 22636
rect 13176 22627 13228 22636
rect 13176 22593 13185 22627
rect 13185 22593 13219 22627
rect 13219 22593 13228 22627
rect 13176 22584 13228 22593
rect 10508 22516 10560 22568
rect 12716 22516 12768 22568
rect 8944 22423 8996 22432
rect 8944 22389 8953 22423
rect 8953 22389 8987 22423
rect 8987 22389 8996 22423
rect 8944 22380 8996 22389
rect 9312 22380 9364 22432
rect 11980 22423 12032 22432
rect 11980 22389 11989 22423
rect 11989 22389 12023 22423
rect 12023 22389 12032 22423
rect 11980 22380 12032 22389
rect 12440 22448 12492 22500
rect 14096 22627 14148 22636
rect 14096 22593 14105 22627
rect 14105 22593 14139 22627
rect 14139 22593 14148 22627
rect 14096 22584 14148 22593
rect 14464 22652 14516 22704
rect 14740 22652 14792 22704
rect 15936 22652 15988 22704
rect 17500 22652 17552 22704
rect 20996 22652 21048 22704
rect 16764 22584 16816 22636
rect 21088 22627 21140 22636
rect 21088 22593 21097 22627
rect 21097 22593 21131 22627
rect 21131 22593 21140 22627
rect 21088 22584 21140 22593
rect 21732 22584 21784 22636
rect 23020 22652 23072 22704
rect 14280 22516 14332 22568
rect 16764 22448 16816 22500
rect 17592 22448 17644 22500
rect 22100 22448 22152 22500
rect 22192 22491 22244 22500
rect 22192 22457 22201 22491
rect 22201 22457 22235 22491
rect 22235 22457 22244 22491
rect 22192 22448 22244 22457
rect 12992 22380 13044 22432
rect 13544 22423 13596 22432
rect 13544 22389 13553 22423
rect 13553 22389 13587 22423
rect 13587 22389 13596 22423
rect 13544 22380 13596 22389
rect 14280 22380 14332 22432
rect 14924 22380 14976 22432
rect 15936 22380 15988 22432
rect 22284 22423 22336 22432
rect 22284 22389 22293 22423
rect 22293 22389 22327 22423
rect 22327 22389 22336 22423
rect 22284 22380 22336 22389
rect 22836 22380 22888 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 8944 22176 8996 22228
rect 9956 22176 10008 22228
rect 10508 22176 10560 22228
rect 8392 22108 8444 22160
rect 3608 21972 3660 22024
rect 6000 21972 6052 22024
rect 6368 21972 6420 22024
rect 5816 21904 5868 21956
rect 6552 22015 6604 22024
rect 6552 21981 6561 22015
rect 6561 21981 6595 22015
rect 6595 21981 6604 22015
rect 6552 21972 6604 21981
rect 8668 22040 8720 22092
rect 9220 22083 9272 22092
rect 9220 22049 9229 22083
rect 9229 22049 9263 22083
rect 9263 22049 9272 22083
rect 9220 22040 9272 22049
rect 9956 22040 10008 22092
rect 12072 22108 12124 22160
rect 12164 22040 12216 22092
rect 10324 21972 10376 22024
rect 11520 22015 11572 22024
rect 11520 21981 11529 22015
rect 11529 21981 11563 22015
rect 11563 21981 11572 22015
rect 11520 21972 11572 21981
rect 5632 21836 5684 21888
rect 6920 21836 6972 21888
rect 9864 21904 9916 21956
rect 10600 21904 10652 21956
rect 11888 22015 11940 22024
rect 11888 21981 11897 22015
rect 11897 21981 11931 22015
rect 11931 21981 11940 22015
rect 11888 21972 11940 21981
rect 12072 22015 12124 22024
rect 12072 21981 12081 22015
rect 12081 21981 12115 22015
rect 12115 21981 12124 22015
rect 12072 21972 12124 21981
rect 12716 22108 12768 22160
rect 8576 21836 8628 21888
rect 9680 21879 9732 21888
rect 9680 21845 9689 21879
rect 9689 21845 9723 21879
rect 9723 21845 9732 21879
rect 9680 21836 9732 21845
rect 11520 21836 11572 21888
rect 12532 22040 12584 22092
rect 12992 22176 13044 22228
rect 13084 22219 13136 22228
rect 13084 22185 13093 22219
rect 13093 22185 13127 22219
rect 13127 22185 13136 22219
rect 13084 22176 13136 22185
rect 13176 22176 13228 22228
rect 15568 22176 15620 22228
rect 13452 22108 13504 22160
rect 13636 22108 13688 22160
rect 14924 22108 14976 22160
rect 15016 22108 15068 22160
rect 16212 22151 16264 22160
rect 16212 22117 16221 22151
rect 16221 22117 16255 22151
rect 16255 22117 16264 22151
rect 16212 22108 16264 22117
rect 12992 22040 13044 22092
rect 13084 22040 13136 22092
rect 13268 22040 13320 22092
rect 13360 22040 13412 22092
rect 12624 22015 12676 22024
rect 12624 21981 12633 22015
rect 12633 21981 12667 22015
rect 12667 21981 12676 22015
rect 12624 21972 12676 21981
rect 12532 21904 12584 21956
rect 12716 21836 12768 21888
rect 13360 21904 13412 21956
rect 13544 21904 13596 21956
rect 15016 21972 15068 22024
rect 16028 22015 16080 22024
rect 16028 21981 16037 22015
rect 16037 21981 16071 22015
rect 16071 21981 16080 22015
rect 16028 21972 16080 21981
rect 15016 21879 15068 21888
rect 15016 21845 15025 21879
rect 15025 21845 15059 21879
rect 15059 21845 15068 21879
rect 15016 21836 15068 21845
rect 15660 21947 15712 21956
rect 15660 21913 15669 21947
rect 15669 21913 15703 21947
rect 15703 21913 15712 21947
rect 15660 21904 15712 21913
rect 15752 21904 15804 21956
rect 16304 22015 16356 22024
rect 16304 21981 16313 22015
rect 16313 21981 16347 22015
rect 16347 21981 16356 22015
rect 16304 21972 16356 21981
rect 16488 22015 16540 22024
rect 16488 21981 16497 22015
rect 16497 21981 16531 22015
rect 16531 21981 16540 22015
rect 16488 21972 16540 21981
rect 16396 21904 16448 21956
rect 17132 22219 17184 22228
rect 17132 22185 17141 22219
rect 17141 22185 17175 22219
rect 17175 22185 17184 22219
rect 17132 22176 17184 22185
rect 17960 22219 18012 22228
rect 17960 22185 17969 22219
rect 17969 22185 18003 22219
rect 18003 22185 18012 22219
rect 17960 22176 18012 22185
rect 22376 22219 22428 22228
rect 22376 22185 22385 22219
rect 22385 22185 22419 22219
rect 22419 22185 22428 22219
rect 22376 22176 22428 22185
rect 18236 22108 18288 22160
rect 19800 22108 19852 22160
rect 19984 22151 20036 22160
rect 19984 22117 19993 22151
rect 19993 22117 20027 22151
rect 20027 22117 20036 22151
rect 19984 22108 20036 22117
rect 20444 22083 20496 22092
rect 20444 22049 20453 22083
rect 20453 22049 20487 22083
rect 20487 22049 20496 22083
rect 20444 22040 20496 22049
rect 22836 22176 22888 22228
rect 17960 21972 18012 22024
rect 17776 21904 17828 21956
rect 18420 22015 18472 22024
rect 18420 21981 18429 22015
rect 18429 21981 18463 22015
rect 18463 21981 18472 22015
rect 18420 21972 18472 21981
rect 22928 22040 22980 22092
rect 20168 21904 20220 21956
rect 22284 21972 22336 22024
rect 22836 22015 22888 22024
rect 22836 21981 22845 22015
rect 22845 21981 22879 22015
rect 22879 21981 22888 22015
rect 22836 21972 22888 21981
rect 23112 22015 23164 22024
rect 23112 21981 23121 22015
rect 23121 21981 23155 22015
rect 23155 21981 23164 22015
rect 23112 21972 23164 21981
rect 17500 21836 17552 21888
rect 19064 21836 19116 21888
rect 19248 21879 19300 21888
rect 19248 21845 19257 21879
rect 19257 21845 19291 21879
rect 19291 21845 19300 21879
rect 19248 21836 19300 21845
rect 19432 21836 19484 21888
rect 19892 21836 19944 21888
rect 19984 21836 20036 21888
rect 22468 21904 22520 21956
rect 23204 21904 23256 21956
rect 20996 21836 21048 21888
rect 23020 21879 23072 21888
rect 23020 21845 23029 21879
rect 23029 21845 23063 21879
rect 23063 21845 23072 21879
rect 23020 21836 23072 21845
rect 4874 21734 4926 21786
rect 4938 21734 4990 21786
rect 5002 21734 5054 21786
rect 5066 21734 5118 21786
rect 5130 21734 5182 21786
rect 4988 21632 5040 21684
rect 4160 21564 4212 21616
rect 6092 21564 6144 21616
rect 9404 21632 9456 21684
rect 4620 21496 4672 21548
rect 5632 21539 5684 21548
rect 5632 21505 5641 21539
rect 5641 21505 5675 21539
rect 5675 21505 5684 21539
rect 5632 21496 5684 21505
rect 6000 21539 6052 21548
rect 6000 21505 6009 21539
rect 6009 21505 6043 21539
rect 6043 21505 6052 21539
rect 6000 21496 6052 21505
rect 12072 21632 12124 21684
rect 12256 21675 12308 21684
rect 12256 21641 12265 21675
rect 12265 21641 12299 21675
rect 12299 21641 12308 21675
rect 12256 21632 12308 21641
rect 12440 21632 12492 21684
rect 12624 21632 12676 21684
rect 12992 21632 13044 21684
rect 11888 21564 11940 21616
rect 16028 21632 16080 21684
rect 17960 21675 18012 21684
rect 17960 21641 17969 21675
rect 17969 21641 18003 21675
rect 18003 21641 18012 21675
rect 17960 21632 18012 21641
rect 6920 21539 6972 21548
rect 6920 21505 6929 21539
rect 6929 21505 6963 21539
rect 6963 21505 6972 21539
rect 6920 21496 6972 21505
rect 7656 21496 7708 21548
rect 5816 21471 5868 21480
rect 4712 21360 4764 21412
rect 2964 21292 3016 21344
rect 5816 21437 5825 21471
rect 5825 21437 5859 21471
rect 5859 21437 5868 21471
rect 5816 21428 5868 21437
rect 6460 21428 6512 21480
rect 8024 21471 8076 21480
rect 8024 21437 8033 21471
rect 8033 21437 8067 21471
rect 8067 21437 8076 21471
rect 8024 21428 8076 21437
rect 8392 21539 8444 21548
rect 8392 21505 8401 21539
rect 8401 21505 8435 21539
rect 8435 21505 8444 21539
rect 8392 21496 8444 21505
rect 8576 21539 8628 21548
rect 8576 21505 8589 21539
rect 8589 21505 8628 21539
rect 8576 21496 8628 21505
rect 10784 21496 10836 21548
rect 11520 21539 11572 21548
rect 11520 21505 11529 21539
rect 11529 21505 11563 21539
rect 11563 21505 11572 21539
rect 11520 21496 11572 21505
rect 11704 21539 11756 21548
rect 11704 21505 11713 21539
rect 11713 21505 11747 21539
rect 11747 21505 11756 21539
rect 11704 21496 11756 21505
rect 9772 21428 9824 21480
rect 6552 21360 6604 21412
rect 9864 21360 9916 21412
rect 7288 21335 7340 21344
rect 7288 21301 7297 21335
rect 7297 21301 7331 21335
rect 7331 21301 7340 21335
rect 7288 21292 7340 21301
rect 8760 21292 8812 21344
rect 12164 21496 12216 21548
rect 12532 21539 12584 21548
rect 12532 21505 12538 21539
rect 12538 21505 12572 21539
rect 12572 21505 12584 21539
rect 12532 21496 12584 21505
rect 15660 21564 15712 21616
rect 18052 21564 18104 21616
rect 18420 21632 18472 21684
rect 18512 21632 18564 21684
rect 22192 21632 22244 21684
rect 22836 21632 22888 21684
rect 13268 21496 13320 21548
rect 13360 21539 13412 21548
rect 13360 21505 13369 21539
rect 13369 21505 13403 21539
rect 13403 21505 13412 21539
rect 13360 21496 13412 21505
rect 13452 21539 13504 21548
rect 13452 21505 13461 21539
rect 13461 21505 13495 21539
rect 13495 21505 13504 21539
rect 13452 21496 13504 21505
rect 13636 21539 13688 21548
rect 13636 21505 13645 21539
rect 13645 21505 13679 21539
rect 13679 21505 13688 21539
rect 13636 21496 13688 21505
rect 13728 21539 13780 21548
rect 13728 21505 13737 21539
rect 13737 21505 13771 21539
rect 13771 21505 13780 21539
rect 13728 21496 13780 21505
rect 15016 21496 15068 21548
rect 12900 21428 12952 21480
rect 15108 21471 15160 21480
rect 15108 21437 15117 21471
rect 15117 21437 15151 21471
rect 15151 21437 15160 21471
rect 15108 21428 15160 21437
rect 15476 21496 15528 21548
rect 16304 21496 16356 21548
rect 16672 21539 16724 21548
rect 16672 21505 16681 21539
rect 16681 21505 16715 21539
rect 16715 21505 16724 21539
rect 16672 21496 16724 21505
rect 16764 21539 16816 21548
rect 16764 21505 16773 21539
rect 16773 21505 16807 21539
rect 16807 21505 16816 21539
rect 16764 21496 16816 21505
rect 16948 21539 17000 21548
rect 16948 21505 16957 21539
rect 16957 21505 16991 21539
rect 16991 21505 17000 21539
rect 16948 21496 17000 21505
rect 17040 21539 17092 21548
rect 17040 21505 17049 21539
rect 17049 21505 17083 21539
rect 17083 21505 17092 21539
rect 17040 21496 17092 21505
rect 17132 21539 17184 21548
rect 17132 21505 17141 21539
rect 17141 21505 17175 21539
rect 17175 21505 17184 21539
rect 17132 21496 17184 21505
rect 17776 21496 17828 21548
rect 19248 21564 19300 21616
rect 22928 21607 22980 21616
rect 22928 21573 22937 21607
rect 22937 21573 22971 21607
rect 22971 21573 22980 21607
rect 22928 21564 22980 21573
rect 23204 21564 23256 21616
rect 18328 21539 18380 21548
rect 18328 21505 18337 21539
rect 18337 21505 18371 21539
rect 18371 21505 18380 21539
rect 18328 21496 18380 21505
rect 18880 21496 18932 21548
rect 17500 21428 17552 21480
rect 10048 21360 10100 21412
rect 11980 21360 12032 21412
rect 10600 21292 10652 21344
rect 12992 21292 13044 21344
rect 15568 21360 15620 21412
rect 20720 21496 20772 21548
rect 21548 21496 21600 21548
rect 19892 21428 19944 21480
rect 20076 21471 20128 21480
rect 20076 21437 20085 21471
rect 20085 21437 20119 21471
rect 20119 21437 20128 21471
rect 20076 21428 20128 21437
rect 19248 21292 19300 21344
rect 21916 21471 21968 21480
rect 21916 21437 21925 21471
rect 21925 21437 21959 21471
rect 21959 21437 21968 21471
rect 21916 21428 21968 21437
rect 22100 21539 22152 21548
rect 22100 21505 22109 21539
rect 22109 21505 22143 21539
rect 22143 21505 22152 21539
rect 22100 21496 22152 21505
rect 22376 21539 22428 21548
rect 22376 21505 22385 21539
rect 22385 21505 22419 21539
rect 22419 21505 22428 21539
rect 22376 21496 22428 21505
rect 21180 21335 21232 21344
rect 21180 21301 21189 21335
rect 21189 21301 21223 21335
rect 21223 21301 21232 21335
rect 21180 21292 21232 21301
rect 21732 21292 21784 21344
rect 22468 21360 22520 21412
rect 22100 21292 22152 21344
rect 22652 21471 22704 21480
rect 22652 21437 22661 21471
rect 22661 21437 22695 21471
rect 22695 21437 22704 21471
rect 22652 21428 22704 21437
rect 23020 21292 23072 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 4988 21131 5040 21140
rect 4988 21097 4997 21131
rect 4997 21097 5031 21131
rect 5031 21097 5040 21131
rect 4988 21088 5040 21097
rect 8300 21131 8352 21140
rect 8300 21097 8309 21131
rect 8309 21097 8343 21131
rect 8343 21097 8352 21131
rect 8300 21088 8352 21097
rect 9680 21088 9732 21140
rect 10416 21088 10468 21140
rect 2780 21020 2832 21072
rect 4528 21020 4580 21072
rect 7288 21020 7340 21072
rect 1400 20995 1452 21004
rect 1400 20961 1409 20995
rect 1409 20961 1443 20995
rect 1443 20961 1452 20995
rect 1400 20952 1452 20961
rect 3056 20884 3108 20936
rect 1676 20859 1728 20868
rect 1676 20825 1685 20859
rect 1685 20825 1719 20859
rect 1719 20825 1728 20859
rect 1676 20816 1728 20825
rect 3608 20927 3660 20936
rect 3608 20893 3617 20927
rect 3617 20893 3651 20927
rect 3651 20893 3660 20927
rect 3608 20884 3660 20893
rect 4712 20952 4764 21004
rect 6368 20952 6420 21004
rect 8116 20952 8168 21004
rect 13728 21088 13780 21140
rect 18236 21131 18288 21140
rect 18236 21097 18245 21131
rect 18245 21097 18279 21131
rect 18279 21097 18288 21131
rect 18236 21088 18288 21097
rect 21640 21088 21692 21140
rect 22652 21088 22704 21140
rect 16948 21020 17000 21072
rect 17960 21020 18012 21072
rect 21916 21020 21968 21072
rect 23112 21020 23164 21072
rect 23480 21020 23532 21072
rect 9864 20952 9916 21004
rect 10232 20952 10284 21004
rect 4160 20927 4212 20936
rect 4160 20893 4169 20927
rect 4169 20893 4203 20927
rect 4203 20893 4212 20927
rect 4160 20884 4212 20893
rect 4620 20927 4672 20936
rect 4620 20893 4629 20927
rect 4629 20893 4663 20927
rect 4663 20893 4672 20927
rect 4620 20884 4672 20893
rect 8576 20927 8628 20936
rect 8576 20893 8585 20927
rect 8585 20893 8619 20927
rect 8619 20893 8628 20927
rect 8576 20884 8628 20893
rect 9588 20927 9640 20936
rect 9588 20893 9597 20927
rect 9597 20893 9631 20927
rect 9631 20893 9640 20927
rect 9588 20884 9640 20893
rect 4068 20816 4120 20868
rect 3240 20791 3292 20800
rect 3240 20757 3249 20791
rect 3249 20757 3283 20791
rect 3283 20757 3292 20791
rect 3240 20748 3292 20757
rect 3608 20748 3660 20800
rect 4528 20748 4580 20800
rect 4804 20748 4856 20800
rect 6184 20816 6236 20868
rect 6460 20859 6512 20868
rect 6460 20825 6469 20859
rect 6469 20825 6503 20859
rect 6503 20825 6512 20859
rect 6460 20816 6512 20825
rect 8300 20859 8352 20868
rect 8300 20825 8309 20859
rect 8309 20825 8343 20859
rect 8343 20825 8352 20859
rect 8300 20816 8352 20825
rect 10048 20859 10100 20868
rect 10048 20825 10057 20859
rect 10057 20825 10091 20859
rect 10091 20825 10100 20859
rect 10048 20816 10100 20825
rect 13360 20995 13412 21004
rect 13360 20961 13369 20995
rect 13369 20961 13403 20995
rect 13403 20961 13412 20995
rect 13360 20952 13412 20961
rect 10508 20927 10560 20936
rect 10508 20893 10517 20927
rect 10517 20893 10551 20927
rect 10551 20893 10560 20927
rect 10508 20884 10560 20893
rect 12992 20884 13044 20936
rect 13820 20884 13872 20936
rect 16396 20952 16448 21004
rect 19064 20952 19116 21004
rect 15752 20884 15804 20936
rect 16028 20884 16080 20936
rect 16764 20884 16816 20936
rect 10784 20816 10836 20868
rect 13912 20816 13964 20868
rect 15844 20816 15896 20868
rect 17500 20816 17552 20868
rect 17868 20816 17920 20868
rect 16304 20748 16356 20800
rect 18696 20791 18748 20800
rect 18696 20757 18705 20791
rect 18705 20757 18739 20791
rect 18739 20757 18748 20791
rect 18696 20748 18748 20757
rect 19064 20859 19116 20868
rect 19064 20825 19073 20859
rect 19073 20825 19107 20859
rect 19107 20825 19116 20859
rect 19064 20816 19116 20825
rect 19248 20927 19300 20936
rect 19248 20893 19257 20927
rect 19257 20893 19291 20927
rect 19291 20893 19300 20927
rect 19248 20884 19300 20893
rect 22376 20952 22428 21004
rect 19708 20927 19760 20936
rect 19708 20893 19717 20927
rect 19717 20893 19751 20927
rect 19751 20893 19760 20927
rect 19708 20884 19760 20893
rect 19800 20884 19852 20936
rect 20168 20927 20220 20936
rect 20168 20893 20181 20927
rect 20181 20893 20220 20927
rect 20168 20884 20220 20893
rect 23020 20927 23072 20936
rect 23020 20893 23029 20927
rect 23029 20893 23063 20927
rect 23063 20893 23072 20927
rect 23020 20884 23072 20893
rect 23388 20927 23440 20936
rect 23388 20893 23397 20927
rect 23397 20893 23431 20927
rect 23431 20893 23440 20927
rect 23388 20884 23440 20893
rect 23480 20927 23532 20936
rect 23480 20893 23489 20927
rect 23489 20893 23523 20927
rect 23523 20893 23532 20927
rect 23480 20884 23532 20893
rect 23664 20927 23716 20936
rect 23664 20893 23673 20927
rect 23673 20893 23707 20927
rect 23707 20893 23716 20927
rect 23664 20884 23716 20893
rect 19248 20748 19300 20800
rect 19432 20748 19484 20800
rect 21640 20748 21692 20800
rect 22744 20791 22796 20800
rect 22744 20757 22753 20791
rect 22753 20757 22787 20791
rect 22787 20757 22796 20791
rect 22744 20748 22796 20757
rect 4874 20646 4926 20698
rect 4938 20646 4990 20698
rect 5002 20646 5054 20698
rect 5066 20646 5118 20698
rect 5130 20646 5182 20698
rect 1676 20544 1728 20596
rect 3608 20544 3660 20596
rect 4068 20544 4120 20596
rect 2964 20476 3016 20528
rect 3240 20519 3292 20528
rect 3240 20485 3249 20519
rect 3249 20485 3283 20519
rect 3283 20485 3292 20519
rect 3240 20476 3292 20485
rect 4528 20476 4580 20528
rect 2780 20451 2832 20460
rect 2780 20417 2789 20451
rect 2789 20417 2823 20451
rect 2823 20417 2832 20451
rect 2780 20408 2832 20417
rect 2872 20451 2924 20460
rect 2872 20417 2881 20451
rect 2881 20417 2915 20451
rect 2915 20417 2924 20451
rect 2872 20408 2924 20417
rect 4620 20408 4672 20460
rect 6184 20476 6236 20528
rect 2688 20340 2740 20392
rect 5448 20408 5500 20460
rect 10048 20544 10100 20596
rect 13360 20544 13412 20596
rect 7380 20476 7432 20528
rect 8208 20519 8260 20528
rect 8208 20485 8219 20519
rect 8219 20485 8260 20519
rect 8208 20476 8260 20485
rect 8392 20519 8444 20528
rect 8392 20485 8401 20519
rect 8401 20485 8435 20519
rect 8435 20485 8444 20519
rect 8392 20476 8444 20485
rect 8668 20519 8720 20528
rect 8668 20485 8677 20519
rect 8677 20485 8711 20519
rect 8711 20485 8720 20519
rect 8668 20476 8720 20485
rect 7656 20408 7708 20460
rect 10600 20476 10652 20528
rect 13084 20476 13136 20528
rect 12808 20451 12860 20460
rect 12808 20417 12817 20451
rect 12817 20417 12851 20451
rect 12851 20417 12860 20451
rect 12808 20408 12860 20417
rect 13452 20451 13504 20460
rect 13452 20417 13461 20451
rect 13461 20417 13495 20451
rect 13495 20417 13504 20451
rect 13452 20408 13504 20417
rect 15568 20544 15620 20596
rect 15936 20544 15988 20596
rect 16212 20544 16264 20596
rect 17040 20544 17092 20596
rect 14648 20476 14700 20528
rect 15568 20451 15620 20460
rect 15568 20417 15577 20451
rect 15577 20417 15611 20451
rect 15611 20417 15620 20451
rect 15568 20408 15620 20417
rect 15844 20476 15896 20528
rect 19708 20544 19760 20596
rect 20076 20544 20128 20596
rect 22008 20544 22060 20596
rect 23664 20544 23716 20596
rect 4620 20272 4672 20324
rect 3608 20204 3660 20256
rect 5356 20315 5408 20324
rect 5356 20281 5365 20315
rect 5365 20281 5399 20315
rect 5399 20281 5408 20315
rect 5356 20272 5408 20281
rect 5264 20204 5316 20256
rect 7104 20340 7156 20392
rect 8576 20340 8628 20392
rect 10600 20340 10652 20392
rect 12900 20383 12952 20392
rect 12900 20349 12909 20383
rect 12909 20349 12943 20383
rect 12943 20349 12952 20383
rect 12900 20340 12952 20349
rect 13636 20340 13688 20392
rect 15660 20383 15712 20392
rect 15660 20349 15669 20383
rect 15669 20349 15703 20383
rect 15703 20349 15712 20383
rect 15660 20340 15712 20349
rect 15936 20408 15988 20460
rect 17500 20451 17552 20460
rect 17500 20417 17508 20451
rect 17508 20417 17542 20451
rect 17542 20417 17552 20451
rect 17500 20408 17552 20417
rect 17960 20408 18012 20460
rect 18696 20476 18748 20528
rect 18788 20451 18840 20460
rect 18788 20417 18797 20451
rect 18797 20417 18831 20451
rect 18831 20417 18840 20451
rect 18788 20408 18840 20417
rect 22192 20476 22244 20528
rect 23204 20476 23256 20528
rect 19800 20408 19852 20460
rect 20996 20451 21048 20460
rect 20996 20417 21005 20451
rect 21005 20417 21039 20451
rect 21039 20417 21048 20451
rect 20996 20408 21048 20417
rect 22100 20408 22152 20460
rect 22468 20451 22520 20460
rect 22468 20417 22477 20451
rect 22477 20417 22511 20451
rect 22511 20417 22520 20451
rect 22468 20408 22520 20417
rect 22652 20408 22704 20460
rect 7380 20272 7432 20324
rect 7656 20204 7708 20256
rect 8116 20204 8168 20256
rect 15108 20272 15160 20324
rect 16672 20272 16724 20324
rect 18144 20383 18196 20392
rect 18144 20349 18153 20383
rect 18153 20349 18187 20383
rect 18187 20349 18196 20383
rect 18144 20340 18196 20349
rect 20720 20340 20772 20392
rect 21180 20340 21232 20392
rect 22744 20340 22796 20392
rect 9312 20204 9364 20256
rect 13820 20247 13872 20256
rect 13820 20213 13829 20247
rect 13829 20213 13863 20247
rect 13863 20213 13872 20247
rect 13820 20204 13872 20213
rect 15936 20247 15988 20256
rect 15936 20213 15945 20247
rect 15945 20213 15979 20247
rect 15979 20213 15988 20247
rect 15936 20204 15988 20213
rect 18420 20247 18472 20256
rect 18420 20213 18429 20247
rect 18429 20213 18463 20247
rect 18463 20213 18472 20247
rect 18420 20204 18472 20213
rect 19984 20247 20036 20256
rect 19984 20213 19993 20247
rect 19993 20213 20027 20247
rect 20027 20213 20036 20247
rect 19984 20204 20036 20213
rect 20996 20204 21048 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 13452 20000 13504 20052
rect 13820 20000 13872 20052
rect 18788 20000 18840 20052
rect 19984 20000 20036 20052
rect 2780 19932 2832 19984
rect 3424 19932 3476 19984
rect 8392 19932 8444 19984
rect 1400 19907 1452 19916
rect 1400 19873 1409 19907
rect 1409 19873 1443 19907
rect 1443 19873 1452 19907
rect 1400 19864 1452 19873
rect 2688 19864 2740 19916
rect 3332 19796 3384 19848
rect 3424 19839 3476 19848
rect 3424 19805 3433 19839
rect 3433 19805 3467 19839
rect 3467 19805 3476 19839
rect 3424 19796 3476 19805
rect 3608 19839 3660 19848
rect 3608 19805 3617 19839
rect 3617 19805 3651 19839
rect 3651 19805 3660 19839
rect 3608 19796 3660 19805
rect 5448 19864 5500 19916
rect 6368 19907 6420 19916
rect 6368 19873 6377 19907
rect 6377 19873 6411 19907
rect 6411 19873 6420 19907
rect 6368 19864 6420 19873
rect 7104 19864 7156 19916
rect 7288 19864 7340 19916
rect 11520 19932 11572 19984
rect 12072 19932 12124 19984
rect 4160 19796 4212 19848
rect 5356 19839 5408 19848
rect 4712 19728 4764 19780
rect 3148 19703 3200 19712
rect 3148 19669 3157 19703
rect 3157 19669 3191 19703
rect 3191 19669 3200 19703
rect 3148 19660 3200 19669
rect 4068 19660 4120 19712
rect 5356 19805 5365 19839
rect 5365 19805 5399 19839
rect 5399 19805 5408 19839
rect 5356 19796 5408 19805
rect 7932 19796 7984 19848
rect 5264 19728 5316 19780
rect 5816 19728 5868 19780
rect 7104 19728 7156 19780
rect 8208 19728 8260 19780
rect 9772 19839 9824 19848
rect 9772 19805 9781 19839
rect 9781 19805 9815 19839
rect 9815 19805 9824 19839
rect 9772 19796 9824 19805
rect 9312 19728 9364 19780
rect 12532 19932 12584 19984
rect 15936 19932 15988 19984
rect 15844 19864 15896 19916
rect 6000 19660 6052 19712
rect 7288 19660 7340 19712
rect 7472 19660 7524 19712
rect 8116 19703 8168 19712
rect 8116 19669 8125 19703
rect 8125 19669 8159 19703
rect 8159 19669 8168 19703
rect 8116 19660 8168 19669
rect 8668 19660 8720 19712
rect 9680 19660 9732 19712
rect 13912 19839 13964 19848
rect 13912 19805 13921 19839
rect 13921 19805 13955 19839
rect 13955 19805 13964 19839
rect 13912 19796 13964 19805
rect 17132 19864 17184 19916
rect 18420 19864 18472 19916
rect 14004 19728 14056 19780
rect 14832 19728 14884 19780
rect 19616 19796 19668 19848
rect 20444 19796 20496 19848
rect 16672 19728 16724 19780
rect 19432 19728 19484 19780
rect 22008 19728 22060 19780
rect 12716 19660 12768 19712
rect 19892 19660 19944 19712
rect 4874 19558 4926 19610
rect 4938 19558 4990 19610
rect 5002 19558 5054 19610
rect 5066 19558 5118 19610
rect 5130 19558 5182 19610
rect 2780 19499 2832 19508
rect 2780 19465 2789 19499
rect 2789 19465 2823 19499
rect 2823 19465 2832 19499
rect 2780 19456 2832 19465
rect 2872 19499 2924 19508
rect 2872 19465 2881 19499
rect 2881 19465 2915 19499
rect 2915 19465 2924 19499
rect 2872 19456 2924 19465
rect 3148 19456 3200 19508
rect 7196 19456 7248 19508
rect 9312 19456 9364 19508
rect 10876 19456 10928 19508
rect 12164 19456 12216 19508
rect 13084 19456 13136 19508
rect 16212 19499 16264 19508
rect 16212 19465 16221 19499
rect 16221 19465 16255 19499
rect 16255 19465 16264 19499
rect 16212 19456 16264 19465
rect 17868 19456 17920 19508
rect 17960 19456 18012 19508
rect 18236 19456 18288 19508
rect 19524 19499 19576 19508
rect 19524 19465 19533 19499
rect 19533 19465 19567 19499
rect 19567 19465 19576 19499
rect 19524 19456 19576 19465
rect 3424 19388 3476 19440
rect 2228 19227 2280 19236
rect 2228 19193 2237 19227
rect 2237 19193 2271 19227
rect 2271 19193 2280 19227
rect 2228 19184 2280 19193
rect 3148 19295 3200 19304
rect 3148 19261 3157 19295
rect 3157 19261 3191 19295
rect 3191 19261 3200 19295
rect 3148 19252 3200 19261
rect 5448 19320 5500 19372
rect 5816 19363 5868 19372
rect 5816 19329 5825 19363
rect 5825 19329 5859 19363
rect 5859 19329 5868 19363
rect 5816 19320 5868 19329
rect 6000 19363 6052 19372
rect 6000 19329 6009 19363
rect 6009 19329 6043 19363
rect 6043 19329 6052 19363
rect 6000 19320 6052 19329
rect 6184 19363 6236 19372
rect 6184 19329 6193 19363
rect 6193 19329 6227 19363
rect 6227 19329 6236 19363
rect 6184 19320 6236 19329
rect 6368 19320 6420 19372
rect 11428 19388 11480 19440
rect 11888 19388 11940 19440
rect 12532 19431 12584 19440
rect 12532 19397 12541 19431
rect 12541 19397 12575 19431
rect 12575 19397 12584 19431
rect 12532 19388 12584 19397
rect 8944 19320 8996 19372
rect 9772 19320 9824 19372
rect 14648 19320 14700 19372
rect 15108 19320 15160 19372
rect 16672 19388 16724 19440
rect 20812 19456 20864 19508
rect 22284 19456 22336 19508
rect 20168 19388 20220 19440
rect 8668 19252 8720 19304
rect 3240 19184 3292 19236
rect 4160 19184 4212 19236
rect 4620 19184 4672 19236
rect 6828 19184 6880 19236
rect 7380 19116 7432 19168
rect 7656 19227 7708 19236
rect 7656 19193 7665 19227
rect 7665 19193 7699 19227
rect 7699 19193 7708 19227
rect 7656 19184 7708 19193
rect 10508 19252 10560 19304
rect 12440 19252 12492 19304
rect 12716 19252 12768 19304
rect 13084 19252 13136 19304
rect 15200 19252 15252 19304
rect 16396 19363 16448 19372
rect 16396 19329 16405 19363
rect 16405 19329 16439 19363
rect 16439 19329 16448 19363
rect 16396 19320 16448 19329
rect 19892 19363 19944 19372
rect 19892 19329 19901 19363
rect 19901 19329 19935 19363
rect 19935 19329 19944 19363
rect 19892 19320 19944 19329
rect 20628 19363 20680 19372
rect 20628 19329 20637 19363
rect 20637 19329 20671 19363
rect 20671 19329 20680 19363
rect 20628 19320 20680 19329
rect 22008 19431 22060 19440
rect 22008 19397 22017 19431
rect 22017 19397 22051 19431
rect 22051 19397 22060 19431
rect 22008 19388 22060 19397
rect 21272 19363 21324 19372
rect 21272 19329 21281 19363
rect 21281 19329 21315 19363
rect 21315 19329 21324 19363
rect 21272 19320 21324 19329
rect 22100 19320 22152 19372
rect 20996 19252 21048 19304
rect 12072 19116 12124 19168
rect 12808 19116 12860 19168
rect 15844 19116 15896 19168
rect 19708 19159 19760 19168
rect 19708 19125 19717 19159
rect 19717 19125 19751 19159
rect 19751 19125 19760 19159
rect 19708 19116 19760 19125
rect 20904 19116 20956 19168
rect 22376 19227 22428 19236
rect 22376 19193 22385 19227
rect 22385 19193 22419 19227
rect 22419 19193 22428 19227
rect 22376 19184 22428 19193
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 3148 18912 3200 18964
rect 4804 18912 4856 18964
rect 6092 18912 6144 18964
rect 7564 18912 7616 18964
rect 9864 18912 9916 18964
rect 3332 18844 3384 18896
rect 3608 18776 3660 18828
rect 8300 18844 8352 18896
rect 4804 18776 4856 18828
rect 6368 18776 6420 18828
rect 6828 18819 6880 18828
rect 6828 18785 6837 18819
rect 6837 18785 6871 18819
rect 6871 18785 6880 18819
rect 6828 18776 6880 18785
rect 9312 18844 9364 18896
rect 9220 18819 9272 18828
rect 9220 18785 9229 18819
rect 9229 18785 9263 18819
rect 9263 18785 9272 18819
rect 11888 18887 11940 18896
rect 11888 18853 11897 18887
rect 11897 18853 11931 18887
rect 11931 18853 11940 18887
rect 12440 18955 12492 18964
rect 12440 18921 12449 18955
rect 12449 18921 12483 18955
rect 12483 18921 12492 18955
rect 12440 18912 12492 18921
rect 12716 18955 12768 18964
rect 12716 18921 12725 18955
rect 12725 18921 12759 18955
rect 12759 18921 12768 18955
rect 12716 18912 12768 18921
rect 15200 18955 15252 18964
rect 15200 18921 15209 18955
rect 15209 18921 15243 18955
rect 15243 18921 15252 18955
rect 15200 18912 15252 18921
rect 15752 18912 15804 18964
rect 15936 18912 15988 18964
rect 18788 18912 18840 18964
rect 18880 18955 18932 18964
rect 18880 18921 18898 18955
rect 18898 18921 18932 18955
rect 18880 18912 18932 18921
rect 19064 18912 19116 18964
rect 19708 18955 19760 18964
rect 19708 18921 19717 18955
rect 19717 18921 19751 18955
rect 19751 18921 19760 18955
rect 19708 18912 19760 18921
rect 20168 18912 20220 18964
rect 20904 18955 20956 18964
rect 20904 18921 20913 18955
rect 20913 18921 20947 18955
rect 20947 18921 20956 18955
rect 20904 18912 20956 18921
rect 22376 18912 22428 18964
rect 11888 18844 11940 18853
rect 15660 18844 15712 18896
rect 9220 18776 9272 18785
rect 3056 18708 3108 18760
rect 3148 18751 3200 18760
rect 3148 18717 3157 18751
rect 3157 18717 3191 18751
rect 3191 18717 3200 18751
rect 3148 18708 3200 18717
rect 3240 18751 3292 18760
rect 3240 18717 3249 18751
rect 3249 18717 3283 18751
rect 3283 18717 3292 18751
rect 3240 18708 3292 18717
rect 2228 18640 2280 18692
rect 3700 18572 3752 18624
rect 5356 18751 5408 18760
rect 5356 18717 5365 18751
rect 5365 18717 5399 18751
rect 5399 18717 5408 18751
rect 5356 18708 5408 18717
rect 8760 18708 8812 18760
rect 8852 18708 8904 18760
rect 4804 18640 4856 18692
rect 8116 18640 8168 18692
rect 9680 18708 9732 18760
rect 5264 18572 5316 18624
rect 7104 18572 7156 18624
rect 8392 18572 8444 18624
rect 12072 18751 12124 18760
rect 12072 18717 12081 18751
rect 12081 18717 12115 18751
rect 12115 18717 12124 18751
rect 12072 18708 12124 18717
rect 12164 18751 12216 18760
rect 12164 18717 12173 18751
rect 12173 18717 12207 18751
rect 12207 18717 12216 18751
rect 12164 18708 12216 18717
rect 10968 18640 11020 18692
rect 13084 18751 13136 18760
rect 13084 18717 13093 18751
rect 13093 18717 13127 18751
rect 13127 18717 13136 18751
rect 13084 18708 13136 18717
rect 16120 18776 16172 18828
rect 17408 18819 17460 18828
rect 17408 18785 17417 18819
rect 17417 18785 17451 18819
rect 17451 18785 17460 18819
rect 17408 18776 17460 18785
rect 13636 18708 13688 18760
rect 15752 18708 15804 18760
rect 13452 18640 13504 18692
rect 12808 18572 12860 18624
rect 12900 18572 12952 18624
rect 15108 18640 15160 18692
rect 15844 18683 15896 18692
rect 15844 18649 15853 18683
rect 15853 18649 15887 18683
rect 15887 18649 15896 18683
rect 15844 18640 15896 18649
rect 16028 18708 16080 18760
rect 17776 18708 17828 18760
rect 18236 18751 18288 18760
rect 18236 18717 18245 18751
rect 18245 18717 18279 18751
rect 18279 18717 18288 18751
rect 18236 18708 18288 18717
rect 17040 18640 17092 18692
rect 18052 18640 18104 18692
rect 18696 18708 18748 18760
rect 21272 18844 21324 18896
rect 20628 18776 20680 18828
rect 20168 18708 20220 18760
rect 22284 18819 22336 18828
rect 22284 18785 22293 18819
rect 22293 18785 22327 18819
rect 22327 18785 22336 18819
rect 22284 18776 22336 18785
rect 21640 18708 21692 18760
rect 16672 18572 16724 18624
rect 16856 18572 16908 18624
rect 18880 18615 18932 18624
rect 18880 18581 18907 18615
rect 18907 18581 18932 18615
rect 18880 18572 18932 18581
rect 19156 18640 19208 18692
rect 19984 18640 20036 18692
rect 19524 18572 19576 18624
rect 20260 18683 20312 18692
rect 20260 18649 20301 18683
rect 20301 18649 20312 18683
rect 20260 18640 20312 18649
rect 20628 18640 20680 18692
rect 20720 18640 20772 18692
rect 21180 18683 21232 18692
rect 21180 18649 21189 18683
rect 21189 18649 21223 18683
rect 21223 18649 21232 18683
rect 21180 18640 21232 18649
rect 20812 18572 20864 18624
rect 20904 18615 20956 18624
rect 20904 18581 20913 18615
rect 20913 18581 20947 18615
rect 20947 18581 20956 18615
rect 20904 18572 20956 18581
rect 21088 18615 21140 18624
rect 21088 18581 21097 18615
rect 21097 18581 21131 18615
rect 21131 18581 21140 18615
rect 21088 18572 21140 18581
rect 23296 18640 23348 18692
rect 22100 18572 22152 18624
rect 4874 18470 4926 18522
rect 4938 18470 4990 18522
rect 5002 18470 5054 18522
rect 5066 18470 5118 18522
rect 5130 18470 5182 18522
rect 3148 18368 3200 18420
rect 5356 18411 5408 18420
rect 5356 18377 5365 18411
rect 5365 18377 5399 18411
rect 5399 18377 5408 18411
rect 5356 18368 5408 18377
rect 7380 18368 7432 18420
rect 8116 18411 8168 18420
rect 8116 18377 8125 18411
rect 8125 18377 8159 18411
rect 8159 18377 8168 18411
rect 8116 18368 8168 18377
rect 8760 18368 8812 18420
rect 10600 18368 10652 18420
rect 13268 18411 13320 18420
rect 13268 18377 13277 18411
rect 13277 18377 13311 18411
rect 13311 18377 13320 18411
rect 13268 18368 13320 18377
rect 15108 18368 15160 18420
rect 17040 18411 17092 18420
rect 17040 18377 17049 18411
rect 17049 18377 17083 18411
rect 17083 18377 17092 18411
rect 17040 18368 17092 18377
rect 3700 18343 3752 18352
rect 3700 18309 3709 18343
rect 3709 18309 3743 18343
rect 3743 18309 3752 18343
rect 3700 18300 3752 18309
rect 4988 18300 5040 18352
rect 7104 18300 7156 18352
rect 7472 18343 7524 18352
rect 7472 18309 7481 18343
rect 7481 18309 7515 18343
rect 7515 18309 7524 18343
rect 7472 18300 7524 18309
rect 7932 18300 7984 18352
rect 9220 18300 9272 18352
rect 10968 18343 11020 18352
rect 10968 18309 10977 18343
rect 10977 18309 11011 18343
rect 11011 18309 11020 18343
rect 10968 18300 11020 18309
rect 11152 18343 11204 18352
rect 11152 18309 11161 18343
rect 11161 18309 11195 18343
rect 11195 18309 11204 18343
rect 11152 18300 11204 18309
rect 12164 18300 12216 18352
rect 12440 18343 12492 18352
rect 12440 18309 12449 18343
rect 12449 18309 12483 18343
rect 12483 18309 12492 18343
rect 12440 18300 12492 18309
rect 2872 18275 2924 18284
rect 2872 18241 2881 18275
rect 2881 18241 2915 18275
rect 2915 18241 2924 18275
rect 2872 18232 2924 18241
rect 3240 18232 3292 18284
rect 6092 18232 6144 18284
rect 8668 18275 8720 18284
rect 8668 18241 8677 18275
rect 8677 18241 8711 18275
rect 8711 18241 8720 18275
rect 8668 18232 8720 18241
rect 10048 18232 10100 18284
rect 2780 18164 2832 18216
rect 3424 18028 3476 18080
rect 13176 18273 13228 18284
rect 13176 18239 13185 18273
rect 13185 18239 13219 18273
rect 13219 18239 13228 18273
rect 13176 18232 13228 18239
rect 13452 18275 13504 18284
rect 13452 18241 13461 18275
rect 13461 18241 13495 18275
rect 13495 18241 13504 18275
rect 13452 18232 13504 18241
rect 13636 18275 13688 18284
rect 13636 18241 13645 18275
rect 13645 18241 13679 18275
rect 13679 18241 13688 18275
rect 13636 18232 13688 18241
rect 15476 18300 15528 18352
rect 15660 18300 15712 18352
rect 16672 18343 16724 18352
rect 16672 18309 16681 18343
rect 16681 18309 16715 18343
rect 16715 18309 16724 18343
rect 19616 18368 19668 18420
rect 19984 18368 20036 18420
rect 16672 18300 16724 18309
rect 18144 18300 18196 18352
rect 20076 18300 20128 18352
rect 21088 18300 21140 18352
rect 13360 18164 13412 18216
rect 16396 18232 16448 18284
rect 22192 18275 22244 18284
rect 22192 18241 22201 18275
rect 22201 18241 22235 18275
rect 22235 18241 22244 18275
rect 22192 18232 22244 18241
rect 16304 18164 16356 18216
rect 20168 18164 20220 18216
rect 21640 18207 21692 18216
rect 21640 18173 21649 18207
rect 21649 18173 21683 18207
rect 21683 18173 21692 18207
rect 21640 18164 21692 18173
rect 22284 18207 22336 18216
rect 22284 18173 22293 18207
rect 22293 18173 22327 18207
rect 22327 18173 22336 18207
rect 22284 18164 22336 18173
rect 19064 18096 19116 18148
rect 20260 18096 20312 18148
rect 5264 18028 5316 18080
rect 12440 18028 12492 18080
rect 12716 18028 12768 18080
rect 12992 18028 13044 18080
rect 17224 18071 17276 18080
rect 17224 18037 17233 18071
rect 17233 18037 17267 18071
rect 17267 18037 17276 18071
rect 17224 18028 17276 18037
rect 17684 18071 17736 18080
rect 17684 18037 17693 18071
rect 17693 18037 17727 18071
rect 17727 18037 17736 18071
rect 17684 18028 17736 18037
rect 19156 18028 19208 18080
rect 20904 18028 20956 18080
rect 23388 18028 23440 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 12072 17867 12124 17876
rect 12072 17833 12081 17867
rect 12081 17833 12115 17867
rect 12115 17833 12124 17867
rect 12072 17824 12124 17833
rect 13176 17824 13228 17876
rect 13636 17824 13688 17876
rect 14740 17824 14792 17876
rect 15568 17824 15620 17876
rect 16856 17867 16908 17876
rect 16856 17833 16865 17867
rect 16865 17833 16899 17867
rect 16899 17833 16908 17867
rect 16856 17824 16908 17833
rect 18880 17824 18932 17876
rect 18972 17867 19024 17876
rect 18972 17833 18981 17867
rect 18981 17833 19015 17867
rect 19015 17833 19024 17867
rect 18972 17824 19024 17833
rect 20812 17824 20864 17876
rect 17040 17756 17092 17808
rect 17408 17756 17460 17808
rect 1400 17731 1452 17740
rect 1400 17697 1409 17731
rect 1409 17697 1443 17731
rect 1443 17697 1452 17731
rect 1400 17688 1452 17697
rect 2688 17688 2740 17740
rect 10600 17731 10652 17740
rect 10600 17697 10609 17731
rect 10609 17697 10643 17731
rect 10643 17697 10652 17731
rect 10600 17688 10652 17697
rect 13912 17688 13964 17740
rect 16304 17731 16356 17740
rect 16304 17697 16313 17731
rect 16313 17697 16347 17731
rect 16347 17697 16356 17731
rect 16304 17688 16356 17697
rect 18420 17688 18472 17740
rect 21640 17688 21692 17740
rect 22008 17688 22060 17740
rect 1860 17620 1912 17672
rect 9588 17620 9640 17672
rect 17224 17663 17276 17672
rect 17224 17629 17233 17663
rect 17233 17629 17267 17663
rect 17267 17629 17276 17663
rect 17224 17620 17276 17629
rect 17960 17620 18012 17672
rect 19064 17663 19116 17672
rect 19064 17629 19073 17663
rect 19073 17629 19107 17663
rect 19107 17629 19116 17663
rect 19064 17620 19116 17629
rect 3332 17552 3384 17604
rect 11336 17552 11388 17604
rect 12716 17552 12768 17604
rect 14004 17552 14056 17604
rect 14740 17552 14792 17604
rect 15568 17552 15620 17604
rect 4160 17484 4212 17536
rect 15200 17484 15252 17536
rect 16120 17552 16172 17604
rect 16580 17552 16632 17604
rect 16396 17484 16448 17536
rect 18328 17484 18380 17536
rect 19524 17595 19576 17604
rect 19524 17561 19533 17595
rect 19533 17561 19567 17595
rect 19567 17561 19576 17595
rect 19524 17552 19576 17561
rect 20076 17552 20128 17604
rect 4874 17382 4926 17434
rect 4938 17382 4990 17434
rect 5002 17382 5054 17434
rect 5066 17382 5118 17434
rect 5130 17382 5182 17434
rect 2872 17280 2924 17332
rect 3424 17280 3476 17332
rect 11152 17280 11204 17332
rect 17684 17280 17736 17332
rect 18052 17280 18104 17332
rect 3332 17212 3384 17264
rect 9864 17255 9916 17264
rect 9864 17221 9873 17255
rect 9873 17221 9907 17255
rect 9907 17221 9916 17255
rect 9864 17212 9916 17221
rect 15936 17212 15988 17264
rect 16396 17212 16448 17264
rect 17040 17255 17092 17264
rect 17040 17221 17049 17255
rect 17049 17221 17083 17255
rect 17083 17221 17092 17255
rect 17040 17212 17092 17221
rect 17500 17212 17552 17264
rect 18328 17212 18380 17264
rect 19156 17280 19208 17332
rect 4160 17187 4212 17196
rect 4160 17153 4169 17187
rect 4169 17153 4203 17187
rect 4203 17153 4212 17187
rect 4160 17144 4212 17153
rect 4620 17144 4672 17196
rect 8668 17144 8720 17196
rect 9588 17187 9640 17196
rect 9588 17153 9597 17187
rect 9597 17153 9631 17187
rect 9631 17153 9640 17187
rect 9588 17144 9640 17153
rect 11336 17144 11388 17196
rect 16304 17144 16356 17196
rect 19432 17144 19484 17196
rect 1860 17076 1912 17128
rect 2964 17076 3016 17128
rect 3424 17076 3476 17128
rect 16580 17076 16632 17128
rect 17500 17076 17552 17128
rect 16120 17008 16172 17060
rect 1768 16940 1820 16992
rect 16212 16940 16264 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 2872 16736 2924 16788
rect 8852 16736 8904 16788
rect 10048 16736 10100 16788
rect 21088 16668 21140 16720
rect 1400 16643 1452 16652
rect 1400 16609 1409 16643
rect 1409 16609 1443 16643
rect 1443 16609 1452 16643
rect 1400 16600 1452 16609
rect 1768 16643 1820 16652
rect 1768 16609 1777 16643
rect 1777 16609 1811 16643
rect 1811 16609 1820 16643
rect 1768 16600 1820 16609
rect 4620 16600 4672 16652
rect 6920 16600 6972 16652
rect 8208 16643 8260 16652
rect 8208 16609 8217 16643
rect 8217 16609 8251 16643
rect 8251 16609 8260 16643
rect 8208 16600 8260 16609
rect 22928 16600 22980 16652
rect 5724 16575 5776 16584
rect 5724 16541 5733 16575
rect 5733 16541 5767 16575
rect 5767 16541 5776 16575
rect 5724 16532 5776 16541
rect 22284 16532 22336 16584
rect 3332 16464 3384 16516
rect 6092 16464 6144 16516
rect 9312 16507 9364 16516
rect 9312 16473 9321 16507
rect 9321 16473 9355 16507
rect 9355 16473 9364 16507
rect 9312 16464 9364 16473
rect 20076 16464 20128 16516
rect 21640 16464 21692 16516
rect 7840 16396 7892 16448
rect 9036 16396 9088 16448
rect 22192 16464 22244 16516
rect 23204 16396 23256 16448
rect 4874 16294 4926 16346
rect 4938 16294 4990 16346
rect 5002 16294 5054 16346
rect 5066 16294 5118 16346
rect 5130 16294 5182 16346
rect 5724 16192 5776 16244
rect 6920 16192 6972 16244
rect 2872 16124 2924 16176
rect 6828 16099 6880 16108
rect 6828 16065 6837 16099
rect 6837 16065 6871 16099
rect 6871 16065 6880 16099
rect 6828 16056 6880 16065
rect 8668 16192 8720 16244
rect 8852 16124 8904 16176
rect 9036 16124 9088 16176
rect 11980 16124 12032 16176
rect 7840 16099 7892 16108
rect 7840 16065 7849 16099
rect 7849 16065 7883 16099
rect 7883 16065 7892 16099
rect 7840 16056 7892 16065
rect 12256 16056 12308 16108
rect 2780 15988 2832 16040
rect 2964 16031 3016 16040
rect 2964 15997 2973 16031
rect 2973 15997 3007 16031
rect 3007 15997 3016 16031
rect 2964 15988 3016 15997
rect 3148 15988 3200 16040
rect 5908 16031 5960 16040
rect 5908 15997 5917 16031
rect 5917 15997 5951 16031
rect 5951 15997 5960 16031
rect 5908 15988 5960 15997
rect 6000 16031 6052 16040
rect 6000 15997 6009 16031
rect 6009 15997 6043 16031
rect 6043 15997 6052 16031
rect 6000 15988 6052 15997
rect 10600 16031 10652 16040
rect 10600 15997 10609 16031
rect 10609 15997 10643 16031
rect 10643 15997 10652 16031
rect 10600 15988 10652 15997
rect 13728 16056 13780 16108
rect 14096 15988 14148 16040
rect 20076 16124 20128 16176
rect 15476 16056 15528 16108
rect 15660 16099 15712 16108
rect 15660 16065 15669 16099
rect 15669 16065 15703 16099
rect 15703 16065 15712 16099
rect 15660 16056 15712 16065
rect 18420 16099 18472 16108
rect 18420 16065 18429 16099
rect 18429 16065 18463 16099
rect 18463 16065 18472 16099
rect 18420 16056 18472 16065
rect 14280 16031 14332 16040
rect 14280 15997 14289 16031
rect 14289 15997 14323 16031
rect 14323 15997 14332 16031
rect 14280 15988 14332 15997
rect 14740 16031 14792 16040
rect 14740 15997 14749 16031
rect 14749 15997 14783 16031
rect 14783 15997 14792 16031
rect 14740 15988 14792 15997
rect 14832 16031 14884 16040
rect 14832 15997 14841 16031
rect 14841 15997 14875 16031
rect 14875 15997 14884 16031
rect 14832 15988 14884 15997
rect 15384 15988 15436 16040
rect 19892 15988 19944 16040
rect 20812 15988 20864 16040
rect 21364 16099 21416 16108
rect 21364 16065 21373 16099
rect 21373 16065 21407 16099
rect 21407 16065 21416 16099
rect 21364 16056 21416 16065
rect 23204 16124 23256 16176
rect 23388 16124 23440 16176
rect 22100 16056 22152 16108
rect 22652 15988 22704 16040
rect 23112 16031 23164 16040
rect 23112 15997 23121 16031
rect 23121 15997 23155 16031
rect 23155 15997 23164 16031
rect 23112 15988 23164 15997
rect 2044 15852 2096 15904
rect 5356 15852 5408 15904
rect 10140 15852 10192 15904
rect 12808 15852 12860 15904
rect 13728 15852 13780 15904
rect 14096 15895 14148 15904
rect 14096 15861 14105 15895
rect 14105 15861 14139 15895
rect 14139 15861 14148 15895
rect 14096 15852 14148 15861
rect 16028 15920 16080 15972
rect 20352 15920 20404 15972
rect 22284 15920 22336 15972
rect 15568 15852 15620 15904
rect 17776 15852 17828 15904
rect 20628 15852 20680 15904
rect 21180 15852 21232 15904
rect 22008 15852 22060 15904
rect 23204 15852 23256 15904
rect 23296 15852 23348 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 6092 15648 6144 15700
rect 7748 15648 7800 15700
rect 8208 15648 8260 15700
rect 1400 15580 1452 15632
rect 2596 15512 2648 15564
rect 4712 15580 4764 15632
rect 4620 15512 4672 15564
rect 5356 15555 5408 15564
rect 5356 15521 5365 15555
rect 5365 15521 5399 15555
rect 5399 15521 5408 15555
rect 5356 15512 5408 15521
rect 6828 15512 6880 15564
rect 10600 15648 10652 15700
rect 14832 15648 14884 15700
rect 12440 15580 12492 15632
rect 13728 15580 13780 15632
rect 14096 15580 14148 15632
rect 15384 15623 15436 15632
rect 15384 15589 15393 15623
rect 15393 15589 15427 15623
rect 15427 15589 15436 15623
rect 15384 15580 15436 15589
rect 15752 15623 15804 15632
rect 15752 15589 15761 15623
rect 15761 15589 15795 15623
rect 15795 15589 15804 15623
rect 15752 15580 15804 15589
rect 9588 15512 9640 15564
rect 10140 15555 10192 15564
rect 10140 15521 10149 15555
rect 10149 15521 10183 15555
rect 10183 15521 10192 15555
rect 10140 15512 10192 15521
rect 1400 15487 1452 15496
rect 1400 15453 1409 15487
rect 1409 15453 1443 15487
rect 1443 15453 1452 15487
rect 1400 15444 1452 15453
rect 2044 15487 2096 15496
rect 2044 15453 2053 15487
rect 2053 15453 2087 15487
rect 2087 15453 2096 15487
rect 2044 15444 2096 15453
rect 2872 15444 2924 15496
rect 8852 15444 8904 15496
rect 9312 15444 9364 15496
rect 12256 15512 12308 15564
rect 10968 15444 11020 15496
rect 12900 15487 12952 15496
rect 12900 15453 12909 15487
rect 12909 15453 12943 15487
rect 12943 15453 12952 15487
rect 12900 15444 12952 15453
rect 13728 15487 13780 15496
rect 13728 15453 13742 15487
rect 13742 15453 13776 15487
rect 13776 15453 13780 15487
rect 13728 15444 13780 15453
rect 14096 15487 14148 15496
rect 14096 15453 14105 15487
rect 14105 15453 14139 15487
rect 14139 15453 14148 15487
rect 14096 15444 14148 15453
rect 19800 15691 19852 15700
rect 19800 15657 19809 15691
rect 19809 15657 19843 15691
rect 19843 15657 19852 15691
rect 19800 15648 19852 15657
rect 21364 15648 21416 15700
rect 20352 15580 20404 15632
rect 22652 15623 22704 15632
rect 22652 15589 22661 15623
rect 22661 15589 22695 15623
rect 22695 15589 22704 15623
rect 22652 15580 22704 15589
rect 16580 15512 16632 15564
rect 3332 15376 3384 15428
rect 3976 15376 4028 15428
rect 6092 15376 6144 15428
rect 2964 15308 3016 15360
rect 3608 15308 3660 15360
rect 4436 15308 4488 15360
rect 7840 15308 7892 15360
rect 9220 15351 9272 15360
rect 9220 15317 9229 15351
rect 9229 15317 9263 15351
rect 9263 15317 9272 15351
rect 9220 15308 9272 15317
rect 9680 15351 9732 15360
rect 9680 15317 9689 15351
rect 9689 15317 9723 15351
rect 9723 15317 9732 15351
rect 9680 15308 9732 15317
rect 10692 15308 10744 15360
rect 10784 15308 10836 15360
rect 11336 15376 11388 15428
rect 12256 15308 12308 15360
rect 12532 15308 12584 15360
rect 13176 15308 13228 15360
rect 13360 15419 13412 15428
rect 13360 15385 13369 15419
rect 13369 15385 13403 15419
rect 13403 15385 13412 15419
rect 13360 15376 13412 15385
rect 13452 15308 13504 15360
rect 13820 15376 13872 15428
rect 15476 15487 15528 15496
rect 15476 15453 15485 15487
rect 15485 15453 15519 15487
rect 15519 15453 15528 15487
rect 15476 15444 15528 15453
rect 15568 15487 15620 15496
rect 15568 15453 15577 15487
rect 15577 15453 15611 15487
rect 15611 15453 15620 15487
rect 15568 15444 15620 15453
rect 15844 15444 15896 15496
rect 16304 15487 16356 15496
rect 16304 15453 16313 15487
rect 16313 15453 16347 15487
rect 16347 15453 16356 15487
rect 16304 15444 16356 15453
rect 20720 15512 20772 15564
rect 20904 15555 20956 15564
rect 20904 15521 20913 15555
rect 20913 15521 20947 15555
rect 20947 15521 20956 15555
rect 20904 15512 20956 15521
rect 21824 15512 21876 15564
rect 23112 15648 23164 15700
rect 23388 15648 23440 15700
rect 23204 15580 23256 15632
rect 20352 15487 20404 15496
rect 20352 15453 20369 15487
rect 20369 15453 20404 15487
rect 17500 15376 17552 15428
rect 19340 15419 19392 15428
rect 19340 15385 19349 15419
rect 19349 15385 19383 15419
rect 19383 15385 19392 15419
rect 20352 15444 20404 15453
rect 20628 15487 20680 15496
rect 20628 15453 20637 15487
rect 20637 15453 20671 15487
rect 20671 15453 20680 15487
rect 20628 15444 20680 15453
rect 23296 15444 23348 15496
rect 19340 15376 19392 15385
rect 14740 15308 14792 15360
rect 16212 15308 16264 15360
rect 17224 15308 17276 15360
rect 21088 15376 21140 15428
rect 21180 15419 21232 15428
rect 21180 15385 21189 15419
rect 21189 15385 21223 15419
rect 21223 15385 21232 15419
rect 21180 15376 21232 15385
rect 21640 15376 21692 15428
rect 22468 15376 22520 15428
rect 24492 15419 24544 15428
rect 24492 15385 24501 15419
rect 24501 15385 24535 15419
rect 24535 15385 24544 15419
rect 24492 15376 24544 15385
rect 20720 15308 20772 15360
rect 20996 15308 21048 15360
rect 21364 15308 21416 15360
rect 23296 15351 23348 15360
rect 23296 15317 23305 15351
rect 23305 15317 23339 15351
rect 23339 15317 23348 15351
rect 23296 15308 23348 15317
rect 24308 15308 24360 15360
rect 4874 15206 4926 15258
rect 4938 15206 4990 15258
rect 5002 15206 5054 15258
rect 5066 15206 5118 15258
rect 5130 15206 5182 15258
rect 112 15104 164 15156
rect 2596 15036 2648 15088
rect 2780 15011 2832 15020
rect 2780 14977 2789 15011
rect 2789 14977 2823 15011
rect 2823 14977 2832 15011
rect 2780 14968 2832 14977
rect 2872 15011 2924 15020
rect 2872 14977 2881 15011
rect 2881 14977 2915 15011
rect 2915 14977 2924 15011
rect 2872 14968 2924 14977
rect 3976 15036 4028 15088
rect 6000 15036 6052 15088
rect 6828 15036 6880 15088
rect 8852 15036 8904 15088
rect 10784 15036 10836 15088
rect 12532 15079 12584 15088
rect 3608 15011 3660 15020
rect 3608 14977 3617 15011
rect 3617 14977 3651 15011
rect 3651 14977 3660 15011
rect 3608 14968 3660 14977
rect 6644 14968 6696 15020
rect 12532 15045 12541 15079
rect 12541 15045 12575 15079
rect 12575 15045 12584 15079
rect 12532 15036 12584 15045
rect 12808 15079 12860 15088
rect 12808 15045 12817 15079
rect 12817 15045 12851 15079
rect 12851 15045 12860 15079
rect 12808 15036 12860 15045
rect 15660 15104 15712 15156
rect 16304 15104 16356 15156
rect 18880 15104 18932 15156
rect 3148 14900 3200 14952
rect 6552 14900 6604 14952
rect 7840 14943 7892 14952
rect 7840 14909 7849 14943
rect 7849 14909 7883 14943
rect 7883 14909 7892 14943
rect 7840 14900 7892 14909
rect 9680 14968 9732 15020
rect 10692 14968 10744 15020
rect 11520 14968 11572 15020
rect 12256 15011 12308 15020
rect 12256 14977 12265 15011
rect 12265 14977 12299 15011
rect 12299 14977 12308 15011
rect 12256 14968 12308 14977
rect 12440 15011 12492 15020
rect 12440 14977 12449 15011
rect 12449 14977 12483 15011
rect 12483 14977 12492 15011
rect 12440 14968 12492 14977
rect 12992 14968 13044 15020
rect 13360 14968 13412 15020
rect 8668 14900 8720 14952
rect 11704 14943 11756 14952
rect 11704 14909 11713 14943
rect 11713 14909 11747 14943
rect 11747 14909 11756 14943
rect 11704 14900 11756 14909
rect 16764 15036 16816 15088
rect 18512 15036 18564 15088
rect 20812 15036 20864 15088
rect 22192 15036 22244 15088
rect 14924 15011 14976 15020
rect 14924 14977 14933 15011
rect 14933 14977 14967 15011
rect 14967 14977 14976 15011
rect 14924 14968 14976 14977
rect 15292 14968 15344 15020
rect 15476 15011 15528 15020
rect 15476 14977 15485 15011
rect 15485 14977 15519 15011
rect 15519 14977 15528 15011
rect 15476 14968 15528 14977
rect 15752 14968 15804 15020
rect 16028 15011 16080 15020
rect 16028 14977 16037 15011
rect 16037 14977 16071 15011
rect 16071 14977 16080 15011
rect 16028 14968 16080 14977
rect 16212 14968 16264 15020
rect 17224 14968 17276 15020
rect 4436 14832 4488 14884
rect 1768 14764 1820 14816
rect 4712 14764 4764 14816
rect 5356 14764 5408 14816
rect 6460 14764 6512 14816
rect 8944 14832 8996 14884
rect 16580 14900 16632 14952
rect 17316 14943 17368 14952
rect 17316 14909 17325 14943
rect 17325 14909 17359 14943
rect 17359 14909 17368 14943
rect 17316 14900 17368 14909
rect 7656 14764 7708 14816
rect 9220 14764 9272 14816
rect 12072 14875 12124 14884
rect 12072 14841 12081 14875
rect 12081 14841 12115 14875
rect 12115 14841 12124 14875
rect 12072 14832 12124 14841
rect 12440 14764 12492 14816
rect 12624 14764 12676 14816
rect 13176 14764 13228 14816
rect 13268 14764 13320 14816
rect 18052 14764 18104 14816
rect 19524 14943 19576 14952
rect 19524 14909 19533 14943
rect 19533 14909 19567 14943
rect 19567 14909 19576 14943
rect 19524 14900 19576 14909
rect 21272 14943 21324 14952
rect 21272 14909 21281 14943
rect 21281 14909 21315 14943
rect 21315 14909 21324 14943
rect 21272 14900 21324 14909
rect 22192 14900 22244 14952
rect 22560 14968 22612 15020
rect 23204 15036 23256 15088
rect 24308 15036 24360 15088
rect 22928 15011 22980 15020
rect 22928 14977 22937 15011
rect 22937 14977 22971 15011
rect 22971 14977 22980 15011
rect 22928 14968 22980 14977
rect 23480 14968 23532 15020
rect 22560 14832 22612 14884
rect 24860 14943 24912 14952
rect 24860 14909 24869 14943
rect 24869 14909 24903 14943
rect 24903 14909 24912 14943
rect 24860 14900 24912 14909
rect 20904 14764 20956 14816
rect 21732 14764 21784 14816
rect 21916 14807 21968 14816
rect 21916 14773 21925 14807
rect 21925 14773 21959 14807
rect 21959 14773 21968 14807
rect 21916 14764 21968 14773
rect 22284 14764 22336 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 2780 14560 2832 14612
rect 3240 14560 3292 14612
rect 5908 14560 5960 14612
rect 6644 14560 6696 14612
rect 6828 14492 6880 14544
rect 1768 14467 1820 14476
rect 1768 14433 1777 14467
rect 1777 14433 1811 14467
rect 1811 14433 1820 14467
rect 1768 14424 1820 14433
rect 3148 14424 3200 14476
rect 6000 14424 6052 14476
rect 6460 14467 6512 14476
rect 6460 14433 6469 14467
rect 6469 14433 6503 14467
rect 6503 14433 6512 14467
rect 6460 14424 6512 14433
rect 6920 14424 6972 14476
rect 1676 14356 1728 14408
rect 3332 14356 3384 14408
rect 5632 14356 5684 14408
rect 6552 14356 6604 14408
rect 6092 14288 6144 14340
rect 6828 14399 6880 14408
rect 6828 14365 6837 14399
rect 6837 14365 6871 14399
rect 6871 14365 6880 14399
rect 6828 14356 6880 14365
rect 8116 14356 8168 14408
rect 9680 14356 9732 14408
rect 12348 14560 12400 14612
rect 13820 14560 13872 14612
rect 14924 14560 14976 14612
rect 15844 14560 15896 14612
rect 17316 14603 17368 14612
rect 17316 14569 17325 14603
rect 17325 14569 17359 14603
rect 17359 14569 17368 14603
rect 17316 14560 17368 14569
rect 19524 14560 19576 14612
rect 21364 14560 21416 14612
rect 22008 14560 22060 14612
rect 22376 14560 22428 14612
rect 12072 14535 12124 14544
rect 12072 14501 12081 14535
rect 12081 14501 12115 14535
rect 12115 14501 12124 14535
rect 12072 14492 12124 14501
rect 14096 14492 14148 14544
rect 12440 14467 12492 14476
rect 12440 14433 12449 14467
rect 12449 14433 12483 14467
rect 12483 14433 12492 14467
rect 12440 14424 12492 14433
rect 11520 14399 11572 14408
rect 11520 14365 11529 14399
rect 11529 14365 11563 14399
rect 11563 14365 11572 14399
rect 11520 14356 11572 14365
rect 11612 14356 11664 14408
rect 9312 14288 9364 14340
rect 10140 14288 10192 14340
rect 11428 14288 11480 14340
rect 11796 14331 11848 14340
rect 11796 14297 11805 14331
rect 11805 14297 11839 14331
rect 11839 14297 11848 14331
rect 11796 14288 11848 14297
rect 12256 14288 12308 14340
rect 14188 14424 14240 14476
rect 12992 14399 13044 14408
rect 12992 14365 13001 14399
rect 13001 14365 13035 14399
rect 13035 14365 13044 14399
rect 12992 14356 13044 14365
rect 13084 14399 13136 14408
rect 13084 14365 13093 14399
rect 13093 14365 13127 14399
rect 13127 14365 13136 14399
rect 13084 14356 13136 14365
rect 13176 14356 13228 14408
rect 13360 14399 13412 14408
rect 13360 14365 13369 14399
rect 13369 14365 13403 14399
rect 13403 14365 13412 14399
rect 13360 14356 13412 14365
rect 13452 14399 13504 14408
rect 13452 14365 13461 14399
rect 13461 14365 13495 14399
rect 13495 14365 13504 14399
rect 13452 14356 13504 14365
rect 4436 14220 4488 14272
rect 4528 14263 4580 14272
rect 4528 14229 4537 14263
rect 4537 14229 4571 14263
rect 4571 14229 4580 14263
rect 4528 14220 4580 14229
rect 4712 14220 4764 14272
rect 5540 14220 5592 14272
rect 7380 14263 7432 14272
rect 7380 14229 7389 14263
rect 7389 14229 7423 14263
rect 7423 14229 7432 14263
rect 7380 14220 7432 14229
rect 10416 14220 10468 14272
rect 12624 14220 12676 14272
rect 12716 14263 12768 14272
rect 12716 14229 12725 14263
rect 12725 14229 12759 14263
rect 12759 14229 12768 14263
rect 12716 14220 12768 14229
rect 12808 14220 12860 14272
rect 17776 14467 17828 14476
rect 17776 14433 17785 14467
rect 17785 14433 17819 14467
rect 17819 14433 17828 14467
rect 17776 14424 17828 14433
rect 21088 14492 21140 14544
rect 21272 14492 21324 14544
rect 23296 14603 23348 14612
rect 23296 14569 23305 14603
rect 23305 14569 23339 14603
rect 23339 14569 23348 14603
rect 23296 14560 23348 14569
rect 20996 14467 21048 14476
rect 20996 14433 21005 14467
rect 21005 14433 21039 14467
rect 21039 14433 21048 14467
rect 20996 14424 21048 14433
rect 18052 14356 18104 14408
rect 21640 14356 21692 14408
rect 21732 14399 21784 14408
rect 21732 14365 21741 14399
rect 21741 14365 21775 14399
rect 21775 14365 21784 14399
rect 21732 14356 21784 14365
rect 21916 14399 21968 14408
rect 21916 14365 21925 14399
rect 21925 14365 21959 14399
rect 21959 14365 21968 14399
rect 21916 14356 21968 14365
rect 22192 14399 22244 14408
rect 22192 14365 22201 14399
rect 22201 14365 22235 14399
rect 22235 14365 22244 14399
rect 22192 14356 22244 14365
rect 22284 14356 22336 14408
rect 13728 14288 13780 14340
rect 14096 14331 14148 14340
rect 14096 14297 14105 14331
rect 14105 14297 14139 14331
rect 14139 14297 14148 14331
rect 14096 14288 14148 14297
rect 14280 14263 14332 14272
rect 14280 14229 14305 14263
rect 14305 14229 14332 14263
rect 15292 14331 15344 14340
rect 15292 14297 15301 14331
rect 15301 14297 15335 14331
rect 15335 14297 15344 14331
rect 15292 14288 15344 14297
rect 20996 14288 21048 14340
rect 23020 14356 23072 14408
rect 23388 14399 23440 14408
rect 23388 14365 23397 14399
rect 23397 14365 23431 14399
rect 23431 14365 23440 14399
rect 23388 14356 23440 14365
rect 23112 14331 23164 14340
rect 23112 14297 23121 14331
rect 23121 14297 23155 14331
rect 23155 14297 23164 14331
rect 23112 14288 23164 14297
rect 14280 14220 14332 14229
rect 15752 14220 15804 14272
rect 4874 14118 4926 14170
rect 4938 14118 4990 14170
rect 5002 14118 5054 14170
rect 5066 14118 5118 14170
rect 5130 14118 5182 14170
rect 1768 14016 1820 14068
rect 4528 14016 4580 14068
rect 7380 14016 7432 14068
rect 8208 14016 8260 14068
rect 3332 13948 3384 14000
rect 848 13880 900 13932
rect 1676 13880 1728 13932
rect 2320 13855 2372 13864
rect 2320 13821 2329 13855
rect 2329 13821 2363 13855
rect 2363 13821 2372 13855
rect 2320 13812 2372 13821
rect 4436 13923 4488 13932
rect 4436 13889 4445 13923
rect 4445 13889 4479 13923
rect 4479 13889 4488 13923
rect 4436 13880 4488 13889
rect 6644 13948 6696 14000
rect 9680 14016 9732 14068
rect 10416 14059 10468 14068
rect 10416 14025 10425 14059
rect 10425 14025 10459 14059
rect 10459 14025 10468 14059
rect 10416 14016 10468 14025
rect 12072 13948 12124 14000
rect 5632 13880 5684 13932
rect 7472 13880 7524 13932
rect 4712 13812 4764 13864
rect 6644 13812 6696 13864
rect 7748 13855 7800 13864
rect 5356 13744 5408 13796
rect 6920 13744 6972 13796
rect 7748 13821 7757 13855
rect 7757 13821 7791 13855
rect 7791 13821 7800 13855
rect 7748 13812 7800 13821
rect 8116 13923 8168 13932
rect 8116 13889 8125 13923
rect 8125 13889 8159 13923
rect 8159 13889 8168 13923
rect 8116 13880 8168 13889
rect 11704 13880 11756 13932
rect 8392 13812 8444 13864
rect 8484 13855 8536 13864
rect 8484 13821 8493 13855
rect 8493 13821 8527 13855
rect 8527 13821 8536 13855
rect 8484 13812 8536 13821
rect 10508 13855 10560 13864
rect 4896 13676 4948 13728
rect 6736 13676 6788 13728
rect 7196 13719 7248 13728
rect 7196 13685 7205 13719
rect 7205 13685 7239 13719
rect 7239 13685 7248 13719
rect 7196 13676 7248 13685
rect 7472 13676 7524 13728
rect 10508 13821 10517 13855
rect 10517 13821 10551 13855
rect 10551 13821 10560 13855
rect 10508 13812 10560 13821
rect 10600 13744 10652 13796
rect 11336 13744 11388 13796
rect 12072 13855 12124 13864
rect 12072 13821 12081 13855
rect 12081 13821 12115 13855
rect 12115 13821 12124 13855
rect 12992 14016 13044 14068
rect 15476 14016 15528 14068
rect 18696 14016 18748 14068
rect 21456 14016 21508 14068
rect 22928 14016 22980 14068
rect 23480 14016 23532 14068
rect 12716 13948 12768 14000
rect 14280 13948 14332 14000
rect 20996 13948 21048 14000
rect 12072 13812 12124 13821
rect 13268 13812 13320 13864
rect 12808 13744 12860 13796
rect 13360 13744 13412 13796
rect 13636 13923 13688 13932
rect 13636 13889 13645 13923
rect 13645 13889 13679 13923
rect 13679 13889 13688 13923
rect 13636 13880 13688 13889
rect 17040 13880 17092 13932
rect 17500 13923 17552 13932
rect 17500 13889 17509 13923
rect 17509 13889 17543 13923
rect 17543 13889 17552 13923
rect 17500 13880 17552 13889
rect 21916 13880 21968 13932
rect 22192 13923 22244 13932
rect 22192 13889 22201 13923
rect 22201 13889 22235 13923
rect 22235 13889 22244 13923
rect 22192 13880 22244 13889
rect 23388 13948 23440 14000
rect 22652 13880 22704 13932
rect 23296 13880 23348 13932
rect 17868 13855 17920 13864
rect 17868 13821 17877 13855
rect 17877 13821 17911 13855
rect 17911 13821 17920 13855
rect 17868 13812 17920 13821
rect 22744 13855 22796 13864
rect 22744 13821 22753 13855
rect 22753 13821 22787 13855
rect 22787 13821 22796 13855
rect 22744 13812 22796 13821
rect 22928 13812 22980 13864
rect 23664 13812 23716 13864
rect 13820 13744 13872 13796
rect 18052 13744 18104 13796
rect 22468 13744 22520 13796
rect 9864 13676 9916 13728
rect 18328 13719 18380 13728
rect 18328 13685 18337 13719
rect 18337 13685 18371 13719
rect 18371 13685 18380 13719
rect 18328 13676 18380 13685
rect 22284 13676 22336 13728
rect 22560 13676 22612 13728
rect 22836 13676 22888 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 2320 13472 2372 13524
rect 8484 13472 8536 13524
rect 11704 13472 11756 13524
rect 14096 13472 14148 13524
rect 16304 13472 16356 13524
rect 18512 13472 18564 13524
rect 21916 13472 21968 13524
rect 22284 13472 22336 13524
rect 22468 13472 22520 13524
rect 3148 13404 3200 13456
rect 3240 13379 3292 13388
rect 3240 13345 3249 13379
rect 3249 13345 3283 13379
rect 3283 13345 3292 13379
rect 3240 13336 3292 13345
rect 8392 13404 8444 13456
rect 11796 13404 11848 13456
rect 17408 13404 17460 13456
rect 17776 13404 17828 13456
rect 4620 13336 4672 13388
rect 4896 13379 4948 13388
rect 4896 13345 4905 13379
rect 4905 13345 4939 13379
rect 4939 13345 4948 13379
rect 4896 13336 4948 13345
rect 5540 13336 5592 13388
rect 6828 13379 6880 13388
rect 6828 13345 6837 13379
rect 6837 13345 6871 13379
rect 6871 13345 6880 13379
rect 6828 13336 6880 13345
rect 7196 13379 7248 13388
rect 7196 13345 7205 13379
rect 7205 13345 7239 13379
rect 7239 13345 7248 13379
rect 7196 13336 7248 13345
rect 9404 13379 9456 13388
rect 9404 13345 9413 13379
rect 9413 13345 9447 13379
rect 9447 13345 9456 13379
rect 9404 13336 9456 13345
rect 9772 13336 9824 13388
rect 10600 13336 10652 13388
rect 4712 13268 4764 13320
rect 6644 13268 6696 13320
rect 11428 13268 11480 13320
rect 8208 13200 8260 13252
rect 11520 13200 11572 13252
rect 13084 13200 13136 13252
rect 15292 13268 15344 13320
rect 15752 13311 15804 13320
rect 15752 13277 15761 13311
rect 15761 13277 15795 13311
rect 15795 13277 15804 13311
rect 15752 13268 15804 13277
rect 16028 13311 16080 13320
rect 16028 13277 16037 13311
rect 16037 13277 16071 13311
rect 16071 13277 16080 13311
rect 16028 13268 16080 13277
rect 16212 13268 16264 13320
rect 16764 13311 16816 13320
rect 16764 13277 16773 13311
rect 16773 13277 16807 13311
rect 16807 13277 16816 13311
rect 16764 13268 16816 13277
rect 17684 13311 17736 13320
rect 17684 13277 17693 13311
rect 17693 13277 17727 13311
rect 17727 13277 17736 13311
rect 17684 13268 17736 13277
rect 17776 13311 17828 13320
rect 17776 13277 17785 13311
rect 17785 13277 17819 13311
rect 17819 13277 17828 13311
rect 17776 13268 17828 13277
rect 18052 13336 18104 13388
rect 21272 13447 21324 13456
rect 21272 13413 21281 13447
rect 21281 13413 21315 13447
rect 21315 13413 21324 13447
rect 21272 13404 21324 13413
rect 22100 13404 22152 13456
rect 23020 13472 23072 13524
rect 23204 13472 23256 13524
rect 23664 13515 23716 13524
rect 23664 13481 23673 13515
rect 23673 13481 23707 13515
rect 23707 13481 23716 13515
rect 23664 13472 23716 13481
rect 6552 13132 6604 13184
rect 9864 13132 9916 13184
rect 11612 13132 11664 13184
rect 17224 13200 17276 13252
rect 17592 13200 17644 13252
rect 20996 13311 21048 13320
rect 20996 13277 21005 13311
rect 21005 13277 21039 13311
rect 21039 13277 21048 13311
rect 20996 13268 21048 13277
rect 21088 13311 21140 13320
rect 21088 13277 21097 13311
rect 21097 13277 21131 13311
rect 21131 13277 21140 13311
rect 21088 13268 21140 13277
rect 21456 13268 21508 13320
rect 21548 13311 21600 13320
rect 21548 13277 21557 13311
rect 21557 13277 21591 13311
rect 21591 13277 21600 13311
rect 21548 13268 21600 13277
rect 22008 13268 22060 13320
rect 22376 13268 22428 13320
rect 23112 13336 23164 13388
rect 23204 13268 23256 13320
rect 23296 13311 23348 13320
rect 23296 13277 23305 13311
rect 23305 13277 23339 13311
rect 23339 13277 23348 13311
rect 23296 13268 23348 13277
rect 23480 13311 23532 13320
rect 23480 13277 23489 13311
rect 23489 13277 23523 13311
rect 23523 13277 23532 13311
rect 24492 13336 24544 13388
rect 23480 13268 23532 13277
rect 15016 13132 15068 13184
rect 16948 13175 17000 13184
rect 16948 13141 16957 13175
rect 16957 13141 16991 13175
rect 16991 13141 17000 13175
rect 16948 13132 17000 13141
rect 17040 13132 17092 13184
rect 18144 13175 18196 13184
rect 18144 13141 18153 13175
rect 18153 13141 18187 13175
rect 18187 13141 18196 13175
rect 18144 13132 18196 13141
rect 18420 13132 18472 13184
rect 20628 13132 20680 13184
rect 21180 13132 21232 13184
rect 22100 13132 22152 13184
rect 22652 13200 22704 13252
rect 23572 13200 23624 13252
rect 24032 13268 24084 13320
rect 24584 13311 24636 13320
rect 24584 13277 24593 13311
rect 24593 13277 24627 13311
rect 24627 13277 24636 13311
rect 24584 13268 24636 13277
rect 24308 13132 24360 13184
rect 24768 13175 24820 13184
rect 24768 13141 24777 13175
rect 24777 13141 24811 13175
rect 24811 13141 24820 13175
rect 24768 13132 24820 13141
rect 4874 13030 4926 13082
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 3240 12928 3292 12980
rect 6644 12928 6696 12980
rect 7472 12928 7524 12980
rect 16764 12928 16816 12980
rect 4620 12860 4672 12912
rect 6276 12792 6328 12844
rect 7104 12860 7156 12912
rect 16304 12860 16356 12912
rect 17132 12903 17184 12912
rect 17132 12869 17141 12903
rect 17141 12869 17175 12903
rect 17175 12869 17184 12903
rect 17132 12860 17184 12869
rect 17500 12860 17552 12912
rect 18696 12928 18748 12980
rect 6736 12835 6788 12844
rect 6736 12801 6745 12835
rect 6745 12801 6779 12835
rect 6779 12801 6788 12835
rect 6736 12792 6788 12801
rect 10692 12792 10744 12844
rect 12072 12835 12124 12844
rect 12072 12801 12081 12835
rect 12081 12801 12115 12835
rect 12115 12801 12124 12835
rect 12072 12792 12124 12801
rect 13820 12792 13872 12844
rect 15016 12835 15068 12844
rect 15016 12801 15025 12835
rect 15025 12801 15059 12835
rect 15059 12801 15068 12835
rect 15016 12792 15068 12801
rect 16764 12792 16816 12844
rect 2320 12656 2372 12708
rect 4712 12724 4764 12776
rect 5356 12767 5408 12776
rect 5356 12733 5365 12767
rect 5365 12733 5399 12767
rect 5399 12733 5408 12767
rect 5356 12724 5408 12733
rect 9588 12767 9640 12776
rect 9588 12733 9597 12767
rect 9597 12733 9631 12767
rect 9631 12733 9640 12767
rect 9588 12724 9640 12733
rect 9772 12767 9824 12776
rect 9772 12733 9781 12767
rect 9781 12733 9815 12767
rect 9815 12733 9824 12767
rect 9772 12724 9824 12733
rect 14648 12767 14700 12776
rect 14648 12733 14657 12767
rect 14657 12733 14691 12767
rect 14691 12733 14700 12767
rect 14648 12724 14700 12733
rect 17040 12792 17092 12844
rect 17224 12835 17276 12844
rect 17224 12801 17233 12835
rect 17233 12801 17267 12835
rect 17267 12801 17276 12835
rect 17224 12792 17276 12801
rect 17684 12860 17736 12912
rect 21364 12971 21416 12980
rect 21364 12937 21373 12971
rect 21373 12937 21407 12971
rect 21407 12937 21416 12971
rect 21364 12928 21416 12937
rect 21456 12928 21508 12980
rect 21640 12928 21692 12980
rect 18328 12767 18380 12776
rect 18328 12733 18337 12767
rect 18337 12733 18371 12767
rect 18371 12733 18380 12767
rect 18328 12724 18380 12733
rect 22468 12971 22520 12980
rect 22468 12937 22477 12971
rect 22477 12937 22511 12971
rect 22511 12937 22520 12971
rect 22468 12928 22520 12937
rect 18696 12792 18748 12844
rect 18788 12767 18840 12776
rect 18788 12733 18797 12767
rect 18797 12733 18831 12767
rect 18831 12733 18840 12767
rect 18788 12724 18840 12733
rect 19708 12835 19760 12844
rect 19708 12801 19717 12835
rect 19717 12801 19751 12835
rect 19751 12801 19760 12835
rect 19708 12792 19760 12801
rect 20904 12724 20956 12776
rect 21088 12724 21140 12776
rect 18236 12656 18288 12708
rect 22560 12835 22612 12844
rect 22560 12801 22569 12835
rect 22569 12801 22603 12835
rect 22603 12801 22612 12835
rect 23480 12860 23532 12912
rect 24032 12860 24084 12912
rect 22560 12792 22612 12801
rect 22836 12792 22888 12844
rect 23020 12835 23072 12844
rect 23020 12801 23029 12835
rect 23029 12801 23063 12835
rect 23063 12801 23072 12835
rect 23020 12792 23072 12801
rect 23112 12835 23164 12844
rect 23112 12801 23121 12835
rect 23121 12801 23155 12835
rect 23155 12801 23164 12835
rect 23112 12792 23164 12801
rect 21916 12724 21968 12776
rect 23388 12792 23440 12844
rect 24308 12835 24360 12844
rect 24308 12801 24317 12835
rect 24317 12801 24351 12835
rect 24351 12801 24360 12835
rect 24308 12792 24360 12801
rect 24492 12835 24544 12844
rect 24492 12801 24501 12835
rect 24501 12801 24535 12835
rect 24535 12801 24544 12835
rect 24492 12792 24544 12801
rect 22376 12656 22428 12708
rect 4068 12588 4120 12640
rect 4804 12631 4856 12640
rect 4804 12597 4813 12631
rect 4813 12597 4847 12631
rect 4847 12597 4856 12631
rect 4804 12588 4856 12597
rect 9128 12631 9180 12640
rect 9128 12597 9137 12631
rect 9137 12597 9171 12631
rect 9171 12597 9180 12631
rect 9128 12588 9180 12597
rect 12164 12631 12216 12640
rect 12164 12597 12173 12631
rect 12173 12597 12207 12631
rect 12207 12597 12216 12631
rect 12164 12588 12216 12597
rect 17408 12588 17460 12640
rect 18420 12588 18472 12640
rect 19984 12588 20036 12640
rect 20996 12631 21048 12640
rect 20996 12597 21005 12631
rect 21005 12597 21039 12631
rect 21039 12597 21048 12631
rect 20996 12588 21048 12597
rect 21180 12588 21232 12640
rect 22468 12588 22520 12640
rect 22836 12631 22888 12640
rect 22836 12597 22845 12631
rect 22845 12597 22879 12631
rect 22879 12597 22888 12631
rect 22836 12588 22888 12597
rect 23388 12631 23440 12640
rect 23388 12597 23397 12631
rect 23397 12597 23431 12631
rect 23431 12597 23440 12631
rect 23388 12588 23440 12597
rect 23572 12631 23624 12640
rect 23572 12597 23581 12631
rect 23581 12597 23615 12631
rect 23615 12597 23624 12631
rect 23572 12588 23624 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 6644 12384 6696 12436
rect 9588 12384 9640 12436
rect 10692 12384 10744 12436
rect 17040 12384 17092 12436
rect 17500 12384 17552 12436
rect 17868 12384 17920 12436
rect 18788 12384 18840 12436
rect 22100 12384 22152 12436
rect 22376 12427 22428 12436
rect 22376 12393 22385 12427
rect 22385 12393 22419 12427
rect 22419 12393 22428 12427
rect 22376 12384 22428 12393
rect 22468 12384 22520 12436
rect 24032 12384 24084 12436
rect 12348 12316 12400 12368
rect 19708 12316 19760 12368
rect 4620 12248 4672 12300
rect 9128 12248 9180 12300
rect 3424 12223 3476 12232
rect 3424 12189 3433 12223
rect 3433 12189 3467 12223
rect 3467 12189 3476 12223
rect 3424 12180 3476 12189
rect 4160 12223 4212 12232
rect 4160 12189 4169 12223
rect 4169 12189 4203 12223
rect 4203 12189 4212 12223
rect 4160 12180 4212 12189
rect 6828 12180 6880 12232
rect 9220 12180 9272 12232
rect 1676 12155 1728 12164
rect 1676 12121 1685 12155
rect 1685 12121 1719 12155
rect 1719 12121 1728 12155
rect 1676 12112 1728 12121
rect 3148 12087 3200 12096
rect 3148 12053 3157 12087
rect 3157 12053 3191 12087
rect 3191 12053 3200 12087
rect 3148 12044 3200 12053
rect 3332 12087 3384 12096
rect 3332 12053 3341 12087
rect 3341 12053 3375 12087
rect 3375 12053 3384 12087
rect 3332 12044 3384 12053
rect 5724 12112 5776 12164
rect 7104 12112 7156 12164
rect 9680 12112 9732 12164
rect 6276 12044 6328 12096
rect 8668 12044 8720 12096
rect 11612 12248 11664 12300
rect 12256 12291 12308 12300
rect 12256 12257 12265 12291
rect 12265 12257 12299 12291
rect 12299 12257 12308 12291
rect 12256 12248 12308 12257
rect 16948 12248 17000 12300
rect 17500 12248 17552 12300
rect 11336 12223 11388 12232
rect 11336 12189 11345 12223
rect 11345 12189 11379 12223
rect 11379 12189 11388 12223
rect 11336 12180 11388 12189
rect 11428 12223 11480 12232
rect 11428 12189 11437 12223
rect 11437 12189 11471 12223
rect 11471 12189 11480 12223
rect 11428 12180 11480 12189
rect 11520 12223 11572 12232
rect 11520 12189 11529 12223
rect 11529 12189 11563 12223
rect 11563 12189 11572 12223
rect 11520 12180 11572 12189
rect 12164 12223 12216 12232
rect 12164 12189 12173 12223
rect 12173 12189 12207 12223
rect 12207 12189 12216 12223
rect 12164 12180 12216 12189
rect 12808 12223 12860 12232
rect 12808 12189 12817 12223
rect 12817 12189 12851 12223
rect 12851 12189 12860 12223
rect 12808 12180 12860 12189
rect 13360 12223 13412 12232
rect 13360 12189 13369 12223
rect 13369 12189 13403 12223
rect 13403 12189 13412 12223
rect 13360 12180 13412 12189
rect 14832 12223 14884 12232
rect 14832 12189 14841 12223
rect 14841 12189 14875 12223
rect 14875 12189 14884 12223
rect 14832 12180 14884 12189
rect 12072 12112 12124 12164
rect 13176 12112 13228 12164
rect 16396 12112 16448 12164
rect 17592 12180 17644 12232
rect 17408 12155 17460 12164
rect 17408 12121 17433 12155
rect 17433 12121 17460 12155
rect 17408 12112 17460 12121
rect 12716 12044 12768 12096
rect 13912 12044 13964 12096
rect 17132 12044 17184 12096
rect 17684 12044 17736 12096
rect 18236 12223 18288 12232
rect 18236 12189 18245 12223
rect 18245 12189 18279 12223
rect 18279 12189 18288 12223
rect 18236 12180 18288 12189
rect 18420 12223 18472 12232
rect 18420 12189 18429 12223
rect 18429 12189 18463 12223
rect 18463 12189 18472 12223
rect 18420 12180 18472 12189
rect 18512 12223 18564 12232
rect 18512 12189 18521 12223
rect 18521 12189 18555 12223
rect 18555 12189 18564 12223
rect 18512 12180 18564 12189
rect 18788 12180 18840 12232
rect 19064 12180 19116 12232
rect 19616 12223 19668 12232
rect 19616 12189 19625 12223
rect 19625 12189 19659 12223
rect 19659 12189 19668 12223
rect 19616 12180 19668 12189
rect 19892 12223 19944 12232
rect 19892 12189 19901 12223
rect 19901 12189 19935 12223
rect 19935 12189 19944 12223
rect 19892 12180 19944 12189
rect 21456 12316 21508 12368
rect 20720 12248 20772 12300
rect 21088 12248 21140 12300
rect 20628 12223 20680 12232
rect 20628 12189 20637 12223
rect 20637 12189 20671 12223
rect 20671 12189 20680 12223
rect 20628 12180 20680 12189
rect 20904 12223 20956 12232
rect 20904 12189 20913 12223
rect 20913 12189 20947 12223
rect 20947 12189 20956 12223
rect 20904 12180 20956 12189
rect 21640 12248 21692 12300
rect 20076 12112 20128 12164
rect 21456 12223 21508 12232
rect 21456 12189 21465 12223
rect 21465 12189 21499 12223
rect 21499 12189 21508 12223
rect 21456 12180 21508 12189
rect 22192 12316 22244 12368
rect 22008 12291 22060 12300
rect 22008 12257 22017 12291
rect 22017 12257 22051 12291
rect 22051 12257 22060 12291
rect 22008 12248 22060 12257
rect 22376 12248 22428 12300
rect 22468 12291 22520 12300
rect 22468 12257 22477 12291
rect 22477 12257 22511 12291
rect 22511 12257 22520 12291
rect 22468 12248 22520 12257
rect 24860 12248 24912 12300
rect 21916 12223 21968 12232
rect 21916 12189 21925 12223
rect 21925 12189 21959 12223
rect 21959 12189 21968 12223
rect 21916 12180 21968 12189
rect 20444 12087 20496 12096
rect 20444 12053 20453 12087
rect 20453 12053 20487 12087
rect 20487 12053 20496 12087
rect 20444 12044 20496 12053
rect 21088 12044 21140 12096
rect 21272 12044 21324 12096
rect 21916 12044 21968 12096
rect 22836 12112 22888 12164
rect 23204 12112 23256 12164
rect 22284 12044 22336 12096
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 1676 11840 1728 11892
rect 6552 11840 6604 11892
rect 8300 11840 8352 11892
rect 9680 11840 9732 11892
rect 5724 11772 5776 11824
rect 6644 11772 6696 11824
rect 10140 11840 10192 11892
rect 11520 11840 11572 11892
rect 11428 11772 11480 11824
rect 12256 11883 12308 11892
rect 12256 11849 12265 11883
rect 12265 11849 12299 11883
rect 12299 11849 12308 11883
rect 12256 11840 12308 11849
rect 18052 11840 18104 11892
rect 18512 11840 18564 11892
rect 18788 11840 18840 11892
rect 1676 11747 1728 11756
rect 1676 11713 1685 11747
rect 1685 11713 1719 11747
rect 1719 11713 1728 11747
rect 1676 11704 1728 11713
rect 2320 11747 2372 11756
rect 2320 11713 2329 11747
rect 2329 11713 2363 11747
rect 2363 11713 2372 11747
rect 2320 11704 2372 11713
rect 3332 11704 3384 11756
rect 4804 11704 4856 11756
rect 6736 11747 6788 11756
rect 6736 11713 6745 11747
rect 6745 11713 6779 11747
rect 6779 11713 6788 11747
rect 6736 11704 6788 11713
rect 8668 11704 8720 11756
rect 9220 11747 9272 11756
rect 9220 11713 9229 11747
rect 9229 11713 9263 11747
rect 9263 11713 9272 11747
rect 9220 11704 9272 11713
rect 11612 11747 11664 11756
rect 11612 11713 11621 11747
rect 11621 11713 11655 11747
rect 11655 11713 11664 11747
rect 11612 11704 11664 11713
rect 12072 11772 12124 11824
rect 12808 11772 12860 11824
rect 17960 11772 18012 11824
rect 3148 11636 3200 11688
rect 4068 11636 4120 11688
rect 4620 11636 4672 11688
rect 6920 11679 6972 11688
rect 6920 11645 6929 11679
rect 6929 11645 6963 11679
rect 6963 11645 6972 11679
rect 6920 11636 6972 11645
rect 7840 11636 7892 11688
rect 9772 11636 9824 11688
rect 12348 11747 12400 11756
rect 12348 11713 12357 11747
rect 12357 11713 12391 11747
rect 12391 11713 12400 11747
rect 12348 11704 12400 11713
rect 12716 11679 12768 11688
rect 12716 11645 12725 11679
rect 12725 11645 12759 11679
rect 12759 11645 12768 11679
rect 12716 11636 12768 11645
rect 13176 11747 13228 11756
rect 13176 11713 13185 11747
rect 13185 11713 13219 11747
rect 13219 11713 13228 11747
rect 13176 11704 13228 11713
rect 13360 11747 13412 11756
rect 13360 11713 13369 11747
rect 13369 11713 13403 11747
rect 13403 11713 13412 11747
rect 13360 11704 13412 11713
rect 13912 11747 13964 11756
rect 13912 11713 13921 11747
rect 13921 11713 13955 11747
rect 13955 11713 13964 11747
rect 13912 11704 13964 11713
rect 18144 11747 18196 11756
rect 18144 11713 18153 11747
rect 18153 11713 18187 11747
rect 18187 11713 18196 11747
rect 18144 11704 18196 11713
rect 19064 11883 19116 11892
rect 19064 11849 19073 11883
rect 19073 11849 19107 11883
rect 19107 11849 19116 11883
rect 19064 11840 19116 11849
rect 19892 11840 19944 11892
rect 19984 11747 20036 11756
rect 19984 11713 19993 11747
rect 19993 11713 20027 11747
rect 20027 11713 20036 11747
rect 19984 11704 20036 11713
rect 20996 11840 21048 11892
rect 24584 11840 24636 11892
rect 20260 11747 20312 11756
rect 20260 11713 20269 11747
rect 20269 11713 20303 11747
rect 20303 11713 20312 11747
rect 20260 11704 20312 11713
rect 19616 11636 19668 11688
rect 20168 11636 20220 11688
rect 21916 11747 21968 11756
rect 21916 11713 21925 11747
rect 21925 11713 21959 11747
rect 21959 11713 21968 11747
rect 21916 11704 21968 11713
rect 21364 11636 21416 11688
rect 22192 11747 22244 11756
rect 22192 11713 22201 11747
rect 22201 11713 22235 11747
rect 22235 11713 22244 11747
rect 22192 11704 22244 11713
rect 22376 11636 22428 11688
rect 23112 11636 23164 11688
rect 848 11500 900 11552
rect 1584 11500 1636 11552
rect 4712 11500 4764 11552
rect 6368 11543 6420 11552
rect 6368 11509 6377 11543
rect 6377 11509 6411 11543
rect 6411 11509 6420 11543
rect 6368 11500 6420 11509
rect 7288 11500 7340 11552
rect 13452 11568 13504 11620
rect 21824 11568 21876 11620
rect 22468 11568 22520 11620
rect 9864 11500 9916 11552
rect 10324 11500 10376 11552
rect 17960 11500 18012 11552
rect 18052 11500 18104 11552
rect 21364 11500 21416 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 1676 11296 1728 11348
rect 3424 11296 3476 11348
rect 6736 11296 6788 11348
rect 8484 11296 8536 11348
rect 8668 11339 8720 11348
rect 8668 11305 8677 11339
rect 8677 11305 8711 11339
rect 8711 11305 8720 11339
rect 8668 11296 8720 11305
rect 9772 11339 9824 11348
rect 9772 11305 9781 11339
rect 9781 11305 9815 11339
rect 9815 11305 9824 11339
rect 9772 11296 9824 11305
rect 15568 11296 15620 11348
rect 17132 11296 17184 11348
rect 20168 11296 20220 11348
rect 20260 11296 20312 11348
rect 21916 11339 21968 11348
rect 21916 11305 21925 11339
rect 21925 11305 21959 11339
rect 21959 11305 21968 11339
rect 21916 11296 21968 11305
rect 22100 11296 22152 11348
rect 10140 11228 10192 11280
rect 11612 11228 11664 11280
rect 1584 11135 1636 11144
rect 1584 11101 1593 11135
rect 1593 11101 1627 11135
rect 1627 11101 1636 11135
rect 1584 11092 1636 11101
rect 3240 11092 3292 11144
rect 4620 11160 4672 11212
rect 6368 11160 6420 11212
rect 6828 11160 6880 11212
rect 7288 11203 7340 11212
rect 7288 11169 7297 11203
rect 7297 11169 7331 11203
rect 7331 11169 7340 11203
rect 7288 11160 7340 11169
rect 4160 11092 4212 11144
rect 6276 11092 6328 11144
rect 4528 11024 4580 11076
rect 3240 10956 3292 11008
rect 4068 10956 4120 11008
rect 4252 10956 4304 11008
rect 5724 11024 5776 11076
rect 8300 11024 8352 11076
rect 10324 11203 10376 11212
rect 10324 11169 10333 11203
rect 10333 11169 10367 11203
rect 10367 11169 10376 11203
rect 10324 11160 10376 11169
rect 12072 11160 12124 11212
rect 13360 11092 13412 11144
rect 20352 11228 20404 11280
rect 22192 11228 22244 11280
rect 14832 11160 14884 11212
rect 15936 11160 15988 11212
rect 16580 11160 16632 11212
rect 20076 11160 20128 11212
rect 13636 11135 13688 11144
rect 13636 11101 13645 11135
rect 13645 11101 13679 11135
rect 13679 11101 13688 11135
rect 13636 11092 13688 11101
rect 13820 11092 13872 11144
rect 15568 11135 15620 11144
rect 15568 11101 15577 11135
rect 15577 11101 15611 11135
rect 15611 11101 15620 11135
rect 15568 11092 15620 11101
rect 19892 11092 19944 11144
rect 20260 11135 20312 11144
rect 20260 11101 20269 11135
rect 20269 11101 20303 11135
rect 20303 11101 20312 11135
rect 20260 11092 20312 11101
rect 21364 11203 21416 11212
rect 21364 11169 21373 11203
rect 21373 11169 21407 11203
rect 21407 11169 21416 11203
rect 21364 11160 21416 11169
rect 22284 11160 22336 11212
rect 20444 11135 20496 11144
rect 20444 11101 20453 11135
rect 20453 11101 20487 11135
rect 20487 11101 20496 11135
rect 20444 11092 20496 11101
rect 20904 11135 20956 11144
rect 20904 11101 20913 11135
rect 20913 11101 20947 11135
rect 20947 11101 20956 11135
rect 20904 11092 20956 11101
rect 10324 11024 10376 11076
rect 10692 11024 10744 11076
rect 11428 11024 11480 11076
rect 16396 11024 16448 11076
rect 17224 11024 17276 11076
rect 17592 11024 17644 11076
rect 18880 11067 18932 11076
rect 18880 11033 18889 11067
rect 18889 11033 18923 11067
rect 18923 11033 18932 11067
rect 21548 11135 21600 11144
rect 21548 11101 21557 11135
rect 21557 11101 21591 11135
rect 21591 11101 21600 11135
rect 21548 11092 21600 11101
rect 22100 11135 22152 11144
rect 22100 11101 22109 11135
rect 22109 11101 22143 11135
rect 22143 11101 22152 11135
rect 22100 11092 22152 11101
rect 22376 11135 22428 11144
rect 22376 11101 22385 11135
rect 22385 11101 22419 11135
rect 22419 11101 22428 11135
rect 22376 11092 22428 11101
rect 18880 11024 18932 11033
rect 10876 10956 10928 11008
rect 12900 10999 12952 11008
rect 12900 10965 12909 10999
rect 12909 10965 12943 10999
rect 12943 10965 12952 10999
rect 12900 10956 12952 10965
rect 13268 10956 13320 11008
rect 13912 10956 13964 11008
rect 19340 10956 19392 11008
rect 20444 10956 20496 11008
rect 22560 11024 22612 11076
rect 23020 11024 23072 11076
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 8944 10752 8996 10804
rect 9036 10752 9088 10804
rect 10876 10752 10928 10804
rect 12900 10752 12952 10804
rect 13820 10752 13872 10804
rect 17132 10795 17184 10804
rect 17132 10761 17141 10795
rect 17141 10761 17175 10795
rect 17175 10761 17184 10795
rect 17132 10752 17184 10761
rect 17592 10795 17644 10804
rect 17592 10761 17601 10795
rect 17601 10761 17635 10795
rect 17635 10761 17644 10795
rect 17592 10752 17644 10761
rect 19892 10752 19944 10804
rect 20904 10752 20956 10804
rect 21548 10795 21600 10804
rect 21548 10761 21557 10795
rect 21557 10761 21591 10795
rect 21591 10761 21600 10795
rect 21548 10752 21600 10761
rect 22376 10752 22428 10804
rect 8300 10684 8352 10736
rect 2780 10659 2832 10668
rect 2780 10625 2789 10659
rect 2789 10625 2823 10659
rect 2823 10625 2832 10659
rect 2780 10616 2832 10625
rect 3148 10616 3200 10668
rect 6920 10616 6972 10668
rect 13268 10659 13320 10668
rect 13268 10625 13276 10659
rect 13276 10625 13310 10659
rect 13310 10625 13320 10659
rect 13268 10616 13320 10625
rect 13360 10659 13412 10668
rect 13360 10625 13369 10659
rect 13369 10625 13403 10659
rect 13403 10625 13412 10659
rect 13360 10616 13412 10625
rect 13452 10659 13504 10668
rect 13452 10625 13461 10659
rect 13461 10625 13495 10659
rect 13495 10625 13504 10659
rect 13452 10616 13504 10625
rect 13728 10659 13780 10668
rect 13728 10625 13737 10659
rect 13737 10625 13771 10659
rect 13771 10625 13780 10659
rect 13728 10616 13780 10625
rect 13820 10659 13872 10668
rect 13820 10625 13829 10659
rect 13829 10625 13863 10659
rect 13863 10625 13872 10659
rect 13820 10616 13872 10625
rect 3424 10548 3476 10600
rect 3976 10548 4028 10600
rect 4252 10548 4304 10600
rect 7748 10591 7800 10600
rect 7748 10557 7757 10591
rect 7757 10557 7791 10591
rect 7791 10557 7800 10591
rect 7748 10548 7800 10557
rect 15936 10659 15988 10668
rect 15936 10625 15945 10659
rect 15945 10625 15979 10659
rect 15979 10625 15988 10659
rect 15936 10616 15988 10625
rect 16764 10616 16816 10668
rect 21824 10684 21876 10736
rect 21272 10659 21324 10668
rect 21272 10625 21281 10659
rect 21281 10625 21315 10659
rect 21315 10625 21324 10659
rect 21272 10616 21324 10625
rect 22468 10659 22520 10668
rect 22468 10625 22477 10659
rect 22477 10625 22511 10659
rect 22511 10625 22520 10659
rect 22468 10616 22520 10625
rect 23388 10616 23440 10668
rect 3516 10480 3568 10532
rect 3148 10412 3200 10464
rect 3332 10412 3384 10464
rect 4160 10455 4212 10464
rect 4160 10421 4169 10455
rect 4169 10421 4203 10455
rect 4203 10421 4212 10455
rect 4160 10412 4212 10421
rect 4620 10412 4672 10464
rect 5356 10412 5408 10464
rect 13544 10412 13596 10464
rect 13728 10480 13780 10532
rect 17316 10548 17368 10600
rect 21548 10591 21600 10600
rect 21548 10557 21557 10591
rect 21557 10557 21591 10591
rect 21591 10557 21600 10591
rect 21548 10548 21600 10557
rect 13912 10412 13964 10464
rect 14004 10455 14056 10464
rect 14004 10421 14013 10455
rect 14013 10421 14047 10455
rect 14047 10421 14056 10455
rect 14004 10412 14056 10421
rect 14372 10455 14424 10464
rect 14372 10421 14381 10455
rect 14381 10421 14415 10455
rect 14415 10421 14424 10455
rect 14372 10412 14424 10421
rect 15200 10412 15252 10464
rect 21180 10412 21232 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 3424 10208 3476 10260
rect 4528 10251 4580 10260
rect 4528 10217 4537 10251
rect 4537 10217 4571 10251
rect 4571 10217 4580 10251
rect 4528 10208 4580 10217
rect 5264 10208 5316 10260
rect 17684 10208 17736 10260
rect 19892 10251 19944 10260
rect 19892 10217 19901 10251
rect 19901 10217 19935 10251
rect 19935 10217 19944 10251
rect 19892 10208 19944 10217
rect 21824 10208 21876 10260
rect 2964 10140 3016 10192
rect 3516 10140 3568 10192
rect 3976 10183 4028 10192
rect 3976 10149 3985 10183
rect 3985 10149 4019 10183
rect 4019 10149 4028 10183
rect 3976 10140 4028 10149
rect 1768 10072 1820 10124
rect 4344 10115 4396 10124
rect 4344 10081 4353 10115
rect 4353 10081 4387 10115
rect 4387 10081 4396 10115
rect 4344 10072 4396 10081
rect 2872 10004 2924 10056
rect 3148 10004 3200 10056
rect 3332 10047 3384 10056
rect 3332 10013 3341 10047
rect 3341 10013 3375 10047
rect 3375 10013 3384 10047
rect 3332 10004 3384 10013
rect 4160 10047 4212 10056
rect 4160 10013 4169 10047
rect 4169 10013 4203 10047
rect 4203 10013 4212 10047
rect 4160 10004 4212 10013
rect 4804 10140 4856 10192
rect 6092 10183 6144 10192
rect 6092 10149 6101 10183
rect 6101 10149 6135 10183
rect 6135 10149 6144 10183
rect 6092 10140 6144 10149
rect 6920 10072 6972 10124
rect 9312 10072 9364 10124
rect 5448 10004 5500 10056
rect 6552 10004 6604 10056
rect 8944 10004 8996 10056
rect 9680 10004 9732 10056
rect 10508 10072 10560 10124
rect 10784 10004 10836 10056
rect 16028 10140 16080 10192
rect 13452 10115 13504 10124
rect 13452 10081 13461 10115
rect 13461 10081 13495 10115
rect 13495 10081 13504 10115
rect 13452 10072 13504 10081
rect 14004 10072 14056 10124
rect 6644 9936 6696 9988
rect 2136 9911 2188 9920
rect 2136 9877 2145 9911
rect 2145 9877 2179 9911
rect 2179 9877 2188 9911
rect 2136 9868 2188 9877
rect 3240 9868 3292 9920
rect 4160 9868 4212 9920
rect 4712 9868 4764 9920
rect 4896 9868 4948 9920
rect 7012 9868 7064 9920
rect 9312 9868 9364 9920
rect 10140 9868 10192 9920
rect 10416 9911 10468 9920
rect 10416 9877 10425 9911
rect 10425 9877 10459 9911
rect 10459 9877 10468 9911
rect 10416 9868 10468 9877
rect 11888 9868 11940 9920
rect 13360 10004 13412 10056
rect 13544 10047 13596 10056
rect 13544 10013 13553 10047
rect 13553 10013 13587 10047
rect 13587 10013 13596 10047
rect 13544 10004 13596 10013
rect 13912 10004 13964 10056
rect 14188 10004 14240 10056
rect 14372 10047 14424 10056
rect 14372 10013 14381 10047
rect 14381 10013 14415 10047
rect 14415 10013 14424 10047
rect 14372 10004 14424 10013
rect 15936 10072 15988 10124
rect 16672 10072 16724 10124
rect 17960 10072 18012 10124
rect 18604 10115 18656 10124
rect 18604 10081 18613 10115
rect 18613 10081 18647 10115
rect 18647 10081 18656 10115
rect 18604 10072 18656 10081
rect 15752 10047 15804 10056
rect 15752 10013 15761 10047
rect 15761 10013 15795 10047
rect 15795 10013 15804 10047
rect 15752 10004 15804 10013
rect 16580 10004 16632 10056
rect 19524 10140 19576 10192
rect 20352 10183 20404 10192
rect 20352 10149 20361 10183
rect 20361 10149 20395 10183
rect 20395 10149 20404 10183
rect 20352 10140 20404 10149
rect 22100 10140 22152 10192
rect 20260 10072 20312 10124
rect 15844 9936 15896 9988
rect 15292 9868 15344 9920
rect 16396 9868 16448 9920
rect 17960 9868 18012 9920
rect 19524 10047 19576 10056
rect 19524 10013 19533 10047
rect 19533 10013 19567 10047
rect 19567 10013 19576 10047
rect 19524 10004 19576 10013
rect 20076 10047 20128 10056
rect 20076 10013 20085 10047
rect 20085 10013 20119 10047
rect 20119 10013 20128 10047
rect 20076 10004 20128 10013
rect 20720 10072 20772 10124
rect 20444 10047 20496 10056
rect 20444 10013 20453 10047
rect 20453 10013 20487 10047
rect 20487 10013 20496 10047
rect 20444 10004 20496 10013
rect 22652 10047 22704 10056
rect 22652 10013 22661 10047
rect 22661 10013 22695 10047
rect 22695 10013 22704 10047
rect 22652 10004 22704 10013
rect 19800 9936 19852 9988
rect 18788 9868 18840 9920
rect 20168 9911 20220 9920
rect 20168 9877 20177 9911
rect 20177 9877 20211 9911
rect 20211 9877 20220 9911
rect 20168 9868 20220 9877
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 4344 9664 4396 9716
rect 4896 9664 4948 9716
rect 5356 9664 5408 9716
rect 6552 9664 6604 9716
rect 9036 9664 9088 9716
rect 10784 9664 10836 9716
rect 2780 9596 2832 9648
rect 3332 9571 3384 9580
rect 3332 9537 3341 9571
rect 3341 9537 3375 9571
rect 3375 9537 3384 9571
rect 3332 9528 3384 9537
rect 4160 9528 4212 9580
rect 5540 9596 5592 9648
rect 6460 9596 6512 9648
rect 3976 9460 4028 9512
rect 4804 9528 4856 9580
rect 5172 9571 5224 9580
rect 5172 9537 5181 9571
rect 5181 9537 5215 9571
rect 5215 9537 5224 9571
rect 5172 9528 5224 9537
rect 5264 9528 5316 9580
rect 6368 9528 6420 9580
rect 6920 9596 6972 9648
rect 8024 9596 8076 9648
rect 10232 9596 10284 9648
rect 14188 9664 14240 9716
rect 4804 9392 4856 9444
rect 5448 9392 5500 9444
rect 6276 9460 6328 9512
rect 6644 9460 6696 9512
rect 7748 9392 7800 9444
rect 3240 9367 3292 9376
rect 3240 9333 3249 9367
rect 3249 9333 3283 9367
rect 3283 9333 3292 9367
rect 3240 9324 3292 9333
rect 3332 9324 3384 9376
rect 4528 9324 4580 9376
rect 5908 9324 5960 9376
rect 7932 9324 7984 9376
rect 8484 9503 8536 9512
rect 8484 9469 8493 9503
rect 8493 9469 8527 9503
rect 8527 9469 8536 9503
rect 8484 9460 8536 9469
rect 11980 9639 12032 9648
rect 11980 9605 11989 9639
rect 11989 9605 12023 9639
rect 12023 9605 12032 9639
rect 11980 9596 12032 9605
rect 12164 9528 12216 9580
rect 12164 9392 12216 9444
rect 13636 9596 13688 9648
rect 16580 9664 16632 9716
rect 17592 9664 17644 9716
rect 20168 9664 20220 9716
rect 13912 9503 13964 9512
rect 13912 9469 13921 9503
rect 13921 9469 13955 9503
rect 13955 9469 13964 9503
rect 13912 9460 13964 9469
rect 15108 9528 15160 9580
rect 15200 9528 15252 9580
rect 14280 9460 14332 9512
rect 15752 9460 15804 9512
rect 16120 9503 16172 9512
rect 16120 9469 16129 9503
rect 16129 9469 16163 9503
rect 16163 9469 16172 9503
rect 16120 9460 16172 9469
rect 17500 9571 17552 9580
rect 17500 9537 17509 9571
rect 17509 9537 17543 9571
rect 17543 9537 17552 9571
rect 17500 9528 17552 9537
rect 18788 9596 18840 9648
rect 21272 9664 21324 9716
rect 17224 9503 17276 9512
rect 17224 9469 17233 9503
rect 17233 9469 17267 9503
rect 17267 9469 17276 9503
rect 17224 9460 17276 9469
rect 12900 9324 12952 9376
rect 15476 9367 15528 9376
rect 15476 9333 15485 9367
rect 15485 9333 15519 9367
rect 15519 9333 15528 9367
rect 15476 9324 15528 9333
rect 15936 9324 15988 9376
rect 19524 9528 19576 9580
rect 19800 9571 19852 9580
rect 19800 9537 19809 9571
rect 19809 9537 19843 9571
rect 19843 9537 19852 9571
rect 19800 9528 19852 9537
rect 19892 9571 19944 9580
rect 19892 9537 19901 9571
rect 19901 9537 19935 9571
rect 19935 9537 19944 9571
rect 19892 9528 19944 9537
rect 20076 9571 20128 9580
rect 20076 9537 20085 9571
rect 20085 9537 20119 9571
rect 20119 9537 20128 9571
rect 20076 9528 20128 9537
rect 20260 9528 20312 9580
rect 20628 9503 20680 9512
rect 20628 9469 20637 9503
rect 20637 9469 20671 9503
rect 20671 9469 20680 9503
rect 20628 9460 20680 9469
rect 21180 9571 21232 9580
rect 21180 9537 21189 9571
rect 21189 9537 21223 9571
rect 21223 9537 21232 9571
rect 21180 9528 21232 9537
rect 22652 9596 22704 9648
rect 21548 9460 21600 9512
rect 20352 9392 20404 9444
rect 20996 9392 21048 9444
rect 21180 9392 21232 9444
rect 22284 9392 22336 9444
rect 17868 9324 17920 9376
rect 18052 9324 18104 9376
rect 19892 9324 19944 9376
rect 21548 9324 21600 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 4436 9120 4488 9172
rect 4804 9120 4856 9172
rect 6092 9163 6144 9172
rect 6092 9129 6101 9163
rect 6101 9129 6135 9163
rect 6135 9129 6144 9163
rect 6092 9120 6144 9129
rect 6276 9163 6328 9172
rect 6276 9129 6285 9163
rect 6285 9129 6319 9163
rect 6319 9129 6328 9163
rect 6276 9120 6328 9129
rect 10232 9120 10284 9172
rect 10968 9120 11020 9172
rect 11888 9120 11940 9172
rect 12348 9120 12400 9172
rect 13636 9120 13688 9172
rect 15384 9120 15436 9172
rect 15936 9120 15988 9172
rect 16120 9120 16172 9172
rect 3056 8984 3108 9036
rect 2780 8916 2832 8968
rect 4068 8984 4120 9036
rect 4344 8984 4396 9036
rect 4804 8984 4856 9036
rect 2504 8780 2556 8832
rect 3608 8959 3660 8968
rect 3608 8925 3617 8959
rect 3617 8925 3651 8959
rect 3651 8925 3660 8959
rect 3608 8916 3660 8925
rect 4712 8916 4764 8968
rect 5540 9052 5592 9104
rect 6644 9052 6696 9104
rect 5632 8984 5684 9036
rect 5724 8984 5776 9036
rect 8024 8984 8076 9036
rect 9588 9052 9640 9104
rect 5264 8916 5316 8968
rect 5356 8959 5408 8968
rect 5356 8925 5365 8959
rect 5365 8925 5399 8959
rect 5399 8925 5408 8959
rect 5356 8916 5408 8925
rect 3516 8848 3568 8900
rect 3424 8780 3476 8832
rect 3792 8823 3844 8832
rect 3792 8789 3801 8823
rect 3801 8789 3835 8823
rect 3835 8789 3844 8823
rect 3792 8780 3844 8789
rect 4068 8823 4120 8832
rect 4068 8789 4077 8823
rect 4077 8789 4111 8823
rect 4111 8789 4120 8823
rect 4068 8780 4120 8789
rect 4252 8891 4304 8900
rect 4252 8857 4261 8891
rect 4261 8857 4295 8891
rect 4295 8857 4304 8891
rect 4252 8848 4304 8857
rect 4436 8891 4488 8900
rect 4436 8857 4445 8891
rect 4445 8857 4479 8891
rect 4479 8857 4488 8891
rect 4436 8848 4488 8857
rect 4804 8848 4856 8900
rect 5540 8959 5592 8968
rect 5540 8925 5549 8959
rect 5549 8925 5583 8959
rect 5583 8925 5592 8959
rect 5540 8916 5592 8925
rect 9680 8984 9732 9036
rect 10416 8984 10468 9036
rect 10784 8984 10836 9036
rect 11796 8984 11848 9036
rect 12164 8916 12216 8968
rect 12348 8916 12400 8968
rect 12532 8959 12584 8968
rect 12532 8925 12541 8959
rect 12541 8925 12575 8959
rect 12575 8925 12584 8959
rect 12532 8916 12584 8925
rect 14280 8984 14332 9036
rect 5908 8891 5960 8900
rect 5908 8857 5917 8891
rect 5917 8857 5951 8891
rect 5951 8857 5960 8891
rect 5908 8848 5960 8857
rect 6736 8848 6788 8900
rect 7288 8848 7340 8900
rect 7932 8848 7984 8900
rect 8852 8848 8904 8900
rect 7380 8780 7432 8832
rect 10968 8848 11020 8900
rect 11888 8780 11940 8832
rect 12900 8891 12952 8900
rect 12900 8857 12909 8891
rect 12909 8857 12943 8891
rect 12943 8857 12952 8891
rect 12900 8848 12952 8857
rect 15476 8916 15528 8968
rect 16672 8916 16724 8968
rect 17500 8984 17552 9036
rect 20628 9120 20680 9172
rect 19892 9027 19944 9036
rect 19892 8993 19901 9027
rect 19901 8993 19935 9027
rect 19935 8993 19944 9027
rect 19892 8984 19944 8993
rect 20628 8984 20680 9036
rect 22468 9052 22520 9104
rect 17040 8916 17092 8968
rect 16396 8848 16448 8900
rect 18788 8916 18840 8968
rect 19064 8916 19116 8968
rect 20076 8959 20128 8968
rect 20076 8925 20085 8959
rect 20085 8925 20119 8959
rect 20119 8925 20128 8959
rect 20076 8916 20128 8925
rect 20720 8916 20772 8968
rect 13176 8823 13228 8832
rect 13176 8789 13185 8823
rect 13185 8789 13219 8823
rect 13219 8789 13228 8823
rect 13176 8780 13228 8789
rect 16764 8780 16816 8832
rect 17408 8780 17460 8832
rect 20444 8848 20496 8900
rect 20996 8959 21048 8968
rect 20996 8925 21005 8959
rect 21005 8925 21039 8959
rect 21039 8925 21048 8959
rect 20996 8916 21048 8925
rect 21456 8959 21508 8968
rect 21456 8925 21465 8959
rect 21465 8925 21499 8959
rect 21499 8925 21508 8959
rect 21456 8916 21508 8925
rect 21180 8780 21232 8832
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 3240 8576 3292 8628
rect 2504 8483 2556 8492
rect 2504 8449 2513 8483
rect 2513 8449 2547 8483
rect 2547 8449 2556 8483
rect 2504 8440 2556 8449
rect 2964 8508 3016 8560
rect 4068 8576 4120 8628
rect 4160 8576 4212 8628
rect 4804 8576 4856 8628
rect 5264 8619 5316 8628
rect 5264 8585 5273 8619
rect 5273 8585 5307 8619
rect 5307 8585 5316 8619
rect 5264 8576 5316 8585
rect 8024 8576 8076 8628
rect 2872 8483 2924 8492
rect 2872 8449 2881 8483
rect 2881 8449 2915 8483
rect 2915 8449 2924 8483
rect 2872 8440 2924 8449
rect 3056 8483 3108 8492
rect 3056 8449 3065 8483
rect 3065 8449 3099 8483
rect 3099 8449 3108 8483
rect 3056 8440 3108 8449
rect 3148 8483 3200 8492
rect 3148 8449 3157 8483
rect 3157 8449 3191 8483
rect 3191 8449 3200 8483
rect 3148 8440 3200 8449
rect 3240 8483 3292 8492
rect 3240 8449 3249 8483
rect 3249 8449 3283 8483
rect 3283 8449 3292 8483
rect 3240 8440 3292 8449
rect 3976 8440 4028 8492
rect 4160 8440 4212 8492
rect 4344 8483 4396 8492
rect 4344 8449 4353 8483
rect 4353 8449 4387 8483
rect 4387 8449 4396 8483
rect 4344 8440 4396 8449
rect 4804 8483 4856 8492
rect 4804 8449 4813 8483
rect 4813 8449 4847 8483
rect 4847 8449 4856 8483
rect 4804 8440 4856 8449
rect 5172 8483 5224 8492
rect 5172 8449 5181 8483
rect 5181 8449 5215 8483
rect 5215 8449 5224 8483
rect 5172 8440 5224 8449
rect 5264 8440 5316 8492
rect 5540 8440 5592 8492
rect 5724 8440 5776 8492
rect 6920 8440 6972 8492
rect 8208 8508 8260 8560
rect 8852 8551 8904 8560
rect 8852 8517 8861 8551
rect 8861 8517 8895 8551
rect 8895 8517 8904 8551
rect 8852 8508 8904 8517
rect 7288 8440 7340 8492
rect 7380 8483 7432 8492
rect 7380 8449 7389 8483
rect 7389 8449 7423 8483
rect 7423 8449 7432 8483
rect 7380 8440 7432 8449
rect 2228 8347 2280 8356
rect 2228 8313 2237 8347
rect 2237 8313 2271 8347
rect 2271 8313 2280 8347
rect 2228 8304 2280 8313
rect 3240 8304 3292 8356
rect 4712 8415 4764 8424
rect 4712 8381 4721 8415
rect 4721 8381 4755 8415
rect 4755 8381 4764 8415
rect 4712 8372 4764 8381
rect 12900 8576 12952 8628
rect 17040 8619 17092 8628
rect 17040 8585 17049 8619
rect 17049 8585 17083 8619
rect 17083 8585 17092 8619
rect 17040 8576 17092 8585
rect 17408 8619 17460 8628
rect 17408 8585 17417 8619
rect 17417 8585 17451 8619
rect 17451 8585 17460 8619
rect 17408 8576 17460 8585
rect 20260 8619 20312 8628
rect 20260 8585 20269 8619
rect 20269 8585 20303 8619
rect 20303 8585 20312 8619
rect 20260 8576 20312 8585
rect 21456 8576 21508 8628
rect 9312 8483 9364 8492
rect 9312 8449 9321 8483
rect 9321 8449 9355 8483
rect 9355 8449 9364 8483
rect 9312 8440 9364 8449
rect 16028 8508 16080 8560
rect 10140 8440 10192 8492
rect 10784 8483 10836 8492
rect 10784 8449 10793 8483
rect 10793 8449 10827 8483
rect 10827 8449 10836 8483
rect 10784 8440 10836 8449
rect 12532 8483 12584 8492
rect 12532 8449 12541 8483
rect 12541 8449 12575 8483
rect 12575 8449 12584 8483
rect 12532 8440 12584 8449
rect 12808 8440 12860 8492
rect 13360 8440 13412 8492
rect 17224 8440 17276 8492
rect 20444 8483 20496 8492
rect 20444 8449 20453 8483
rect 20453 8449 20487 8483
rect 20487 8449 20496 8483
rect 20444 8440 20496 8449
rect 20720 8440 20772 8492
rect 10232 8372 10284 8424
rect 12164 8372 12216 8424
rect 15936 8372 15988 8424
rect 18604 8372 18656 8424
rect 3976 8236 4028 8288
rect 4896 8304 4948 8356
rect 6368 8304 6420 8356
rect 5172 8236 5224 8288
rect 5632 8236 5684 8288
rect 7196 8236 7248 8288
rect 12992 8236 13044 8288
rect 13636 8279 13688 8288
rect 13636 8245 13645 8279
rect 13645 8245 13679 8279
rect 13679 8245 13688 8279
rect 13636 8236 13688 8245
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 3056 8032 3108 8084
rect 3332 8075 3384 8084
rect 3332 8041 3341 8075
rect 3341 8041 3375 8075
rect 3375 8041 3384 8075
rect 3332 8032 3384 8041
rect 3608 8075 3660 8084
rect 3608 8041 3617 8075
rect 3617 8041 3651 8075
rect 3651 8041 3660 8075
rect 3608 8032 3660 8041
rect 12256 8032 12308 8084
rect 16580 8032 16632 8084
rect 17776 8032 17828 8084
rect 2964 8007 3016 8016
rect 2964 7973 2973 8007
rect 2973 7973 3007 8007
rect 3007 7973 3016 8007
rect 2964 7964 3016 7973
rect 5264 7964 5316 8016
rect 6368 7964 6420 8016
rect 6920 7964 6972 8016
rect 3148 7896 3200 7948
rect 3240 7939 3292 7948
rect 3240 7905 3249 7939
rect 3249 7905 3283 7939
rect 3283 7905 3292 7939
rect 3240 7896 3292 7905
rect 3700 7896 3752 7948
rect 3424 7871 3476 7880
rect 3424 7837 3433 7871
rect 3433 7837 3467 7871
rect 3467 7837 3476 7871
rect 3424 7828 3476 7837
rect 3976 7871 4028 7880
rect 3976 7837 3985 7871
rect 3985 7837 4019 7871
rect 4019 7837 4028 7871
rect 3976 7828 4028 7837
rect 2872 7692 2924 7744
rect 3884 7760 3936 7812
rect 4896 7896 4948 7948
rect 5724 7896 5776 7948
rect 4344 7871 4396 7880
rect 4344 7837 4353 7871
rect 4353 7837 4387 7871
rect 4387 7837 4396 7871
rect 4344 7828 4396 7837
rect 5448 7828 5500 7880
rect 12992 7939 13044 7948
rect 12992 7905 13001 7939
rect 13001 7905 13035 7939
rect 13035 7905 13044 7939
rect 12992 7896 13044 7905
rect 13820 8007 13872 8016
rect 13820 7973 13829 8007
rect 13829 7973 13863 8007
rect 13863 7973 13872 8007
rect 13820 7964 13872 7973
rect 4712 7760 4764 7812
rect 6736 7828 6788 7880
rect 6920 7871 6972 7880
rect 6920 7837 6929 7871
rect 6929 7837 6963 7871
rect 6963 7837 6972 7871
rect 6920 7828 6972 7837
rect 7196 7828 7248 7880
rect 7288 7828 7340 7880
rect 9680 7828 9732 7880
rect 12348 7871 12400 7880
rect 12348 7837 12357 7871
rect 12357 7837 12391 7871
rect 12391 7837 12400 7871
rect 12348 7828 12400 7837
rect 12440 7871 12492 7880
rect 12440 7837 12449 7871
rect 12449 7837 12483 7871
rect 12483 7837 12492 7871
rect 12440 7828 12492 7837
rect 13268 7871 13320 7880
rect 13268 7837 13277 7871
rect 13277 7837 13311 7871
rect 13311 7837 13320 7871
rect 14280 7939 14332 7948
rect 14280 7905 14289 7939
rect 14289 7905 14323 7939
rect 14323 7905 14332 7939
rect 14280 7896 14332 7905
rect 13268 7828 13320 7837
rect 14648 7871 14700 7880
rect 14648 7837 14657 7871
rect 14657 7837 14691 7871
rect 14691 7837 14700 7871
rect 14648 7828 14700 7837
rect 18512 7871 18564 7880
rect 18512 7837 18521 7871
rect 18521 7837 18555 7871
rect 18555 7837 18564 7871
rect 18512 7828 18564 7837
rect 4252 7692 4304 7744
rect 13176 7760 13228 7812
rect 16396 7760 16448 7812
rect 5448 7735 5500 7744
rect 5448 7701 5457 7735
rect 5457 7701 5491 7735
rect 5491 7701 5500 7735
rect 5448 7692 5500 7701
rect 5908 7692 5960 7744
rect 6736 7692 6788 7744
rect 7380 7692 7432 7744
rect 13360 7692 13412 7744
rect 13452 7735 13504 7744
rect 13452 7701 13461 7735
rect 13461 7701 13495 7735
rect 13495 7701 13504 7735
rect 13452 7692 13504 7701
rect 18788 7735 18840 7744
rect 18788 7701 18797 7735
rect 18797 7701 18831 7735
rect 18831 7701 18840 7735
rect 18788 7692 18840 7701
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 2872 7531 2924 7540
rect 2872 7497 2881 7531
rect 2881 7497 2915 7531
rect 2915 7497 2924 7531
rect 2872 7488 2924 7497
rect 4068 7488 4120 7540
rect 4160 7531 4212 7540
rect 4160 7497 4169 7531
rect 4169 7497 4203 7531
rect 4203 7497 4212 7531
rect 4160 7488 4212 7497
rect 4344 7488 4396 7540
rect 5264 7488 5316 7540
rect 5356 7488 5408 7540
rect 7380 7488 7432 7540
rect 9404 7488 9456 7540
rect 10324 7488 10376 7540
rect 13268 7488 13320 7540
rect 14648 7488 14700 7540
rect 3608 7420 3660 7472
rect 3148 7395 3200 7404
rect 3148 7361 3156 7395
rect 3156 7361 3190 7395
rect 3190 7361 3200 7395
rect 3148 7352 3200 7361
rect 3516 7352 3568 7404
rect 3884 7352 3936 7404
rect 4252 7395 4304 7404
rect 4252 7361 4261 7395
rect 4261 7361 4295 7395
rect 4295 7361 4304 7395
rect 4252 7352 4304 7361
rect 5172 7420 5224 7472
rect 5356 7352 5408 7404
rect 6736 7463 6788 7472
rect 6736 7429 6745 7463
rect 6745 7429 6779 7463
rect 6779 7429 6788 7463
rect 6736 7420 6788 7429
rect 4896 7284 4948 7336
rect 4988 7216 5040 7268
rect 5908 7395 5960 7404
rect 5908 7361 5917 7395
rect 5917 7361 5951 7395
rect 5951 7361 5960 7395
rect 5908 7352 5960 7361
rect 6552 7395 6604 7404
rect 6552 7361 6561 7395
rect 6561 7361 6595 7395
rect 6595 7361 6604 7395
rect 6552 7352 6604 7361
rect 9864 7352 9916 7404
rect 10140 7395 10192 7404
rect 10140 7361 10149 7395
rect 10149 7361 10183 7395
rect 10183 7361 10192 7395
rect 10140 7352 10192 7361
rect 9680 7284 9732 7336
rect 11704 7395 11756 7404
rect 11704 7361 11713 7395
rect 11713 7361 11747 7395
rect 11747 7361 11756 7395
rect 11704 7352 11756 7361
rect 13636 7420 13688 7472
rect 12256 7395 12308 7404
rect 12256 7361 12265 7395
rect 12265 7361 12299 7395
rect 12299 7361 12308 7395
rect 12256 7352 12308 7361
rect 12348 7352 12400 7404
rect 12900 7352 12952 7404
rect 12440 7284 12492 7336
rect 13452 7352 13504 7404
rect 13820 7284 13872 7336
rect 16580 7420 16632 7472
rect 19616 7488 19668 7540
rect 18604 7420 18656 7472
rect 16948 7395 17000 7404
rect 16948 7361 16957 7395
rect 16957 7361 16991 7395
rect 16991 7361 17000 7395
rect 16948 7352 17000 7361
rect 17132 7395 17184 7404
rect 17132 7361 17141 7395
rect 17141 7361 17175 7395
rect 17175 7361 17184 7395
rect 17132 7352 17184 7361
rect 17224 7284 17276 7336
rect 3240 7148 3292 7200
rect 6000 7191 6052 7200
rect 6000 7157 6009 7191
rect 6009 7157 6043 7191
rect 6043 7157 6052 7191
rect 6000 7148 6052 7157
rect 8300 7148 8352 7200
rect 9772 7191 9824 7200
rect 9772 7157 9781 7191
rect 9781 7157 9815 7191
rect 9815 7157 9824 7191
rect 9772 7148 9824 7157
rect 10324 7148 10376 7200
rect 10692 7191 10744 7200
rect 10692 7157 10701 7191
rect 10701 7157 10735 7191
rect 10735 7157 10744 7191
rect 10692 7148 10744 7157
rect 13728 7216 13780 7268
rect 18144 7284 18196 7336
rect 21364 7216 21416 7268
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 3608 6987 3660 6996
rect 3608 6953 3617 6987
rect 3617 6953 3651 6987
rect 3651 6953 3660 6987
rect 3608 6944 3660 6953
rect 3884 6876 3936 6928
rect 2136 6808 2188 6860
rect 2504 6851 2556 6860
rect 2504 6817 2513 6851
rect 2513 6817 2547 6851
rect 2547 6817 2556 6851
rect 2504 6808 2556 6817
rect 4712 6944 4764 6996
rect 4896 6987 4948 6996
rect 4896 6953 4905 6987
rect 4905 6953 4939 6987
rect 4939 6953 4948 6987
rect 4896 6944 4948 6953
rect 5080 6944 5132 6996
rect 9588 6944 9640 6996
rect 10140 6944 10192 6996
rect 11060 6944 11112 6996
rect 11612 6944 11664 6996
rect 11704 6944 11756 6996
rect 12256 6944 12308 6996
rect 12532 6944 12584 6996
rect 16948 6944 17000 6996
rect 18604 6944 18656 6996
rect 19984 6944 20036 6996
rect 20720 6944 20772 6996
rect 2228 6740 2280 6792
rect 3148 6672 3200 6724
rect 3516 6740 3568 6792
rect 4896 6808 4948 6860
rect 5264 6851 5316 6860
rect 5264 6817 5273 6851
rect 5273 6817 5307 6851
rect 5307 6817 5316 6851
rect 5264 6808 5316 6817
rect 1676 6604 1728 6656
rect 3884 6647 3936 6656
rect 3884 6613 3893 6647
rect 3893 6613 3927 6647
rect 3927 6613 3936 6647
rect 3884 6604 3936 6613
rect 4160 6740 4212 6792
rect 4252 6715 4304 6724
rect 4252 6681 4261 6715
rect 4261 6681 4295 6715
rect 4295 6681 4304 6715
rect 4252 6672 4304 6681
rect 5356 6740 5408 6792
rect 7012 6808 7064 6860
rect 8484 6851 8536 6860
rect 8484 6817 8493 6851
rect 8493 6817 8527 6851
rect 8527 6817 8536 6851
rect 8484 6808 8536 6817
rect 9772 6808 9824 6860
rect 7840 6740 7892 6792
rect 8024 6740 8076 6792
rect 6828 6672 6880 6724
rect 10140 6672 10192 6724
rect 11152 6672 11204 6724
rect 12164 6876 12216 6928
rect 11612 6808 11664 6860
rect 12900 6876 12952 6928
rect 17132 6808 17184 6860
rect 18052 6851 18104 6860
rect 18052 6817 18061 6851
rect 18061 6817 18095 6851
rect 18095 6817 18104 6851
rect 18052 6808 18104 6817
rect 18144 6808 18196 6860
rect 20812 6808 20864 6860
rect 12440 6783 12492 6792
rect 12440 6749 12449 6783
rect 12449 6749 12483 6783
rect 12483 6749 12492 6783
rect 12440 6740 12492 6749
rect 12624 6783 12676 6792
rect 12624 6749 12633 6783
rect 12633 6749 12667 6783
rect 12667 6749 12676 6783
rect 12624 6740 12676 6749
rect 12900 6783 12952 6792
rect 12900 6749 12909 6783
rect 12909 6749 12943 6783
rect 12943 6749 12952 6783
rect 12900 6740 12952 6749
rect 11612 6672 11664 6724
rect 11796 6715 11848 6724
rect 11796 6681 11805 6715
rect 11805 6681 11839 6715
rect 11839 6681 11848 6715
rect 11796 6672 11848 6681
rect 11888 6715 11940 6724
rect 11888 6681 11897 6715
rect 11897 6681 11931 6715
rect 11931 6681 11940 6715
rect 11888 6672 11940 6681
rect 12808 6672 12860 6724
rect 15660 6715 15712 6724
rect 15660 6681 15669 6715
rect 15669 6681 15703 6715
rect 15703 6681 15712 6715
rect 15660 6672 15712 6681
rect 6552 6604 6604 6656
rect 7288 6604 7340 6656
rect 7564 6647 7616 6656
rect 7564 6613 7573 6647
rect 7573 6613 7607 6647
rect 7607 6613 7616 6647
rect 7564 6604 7616 6613
rect 8116 6604 8168 6656
rect 9588 6604 9640 6656
rect 12256 6604 12308 6656
rect 13728 6604 13780 6656
rect 16580 6672 16632 6724
rect 17224 6672 17276 6724
rect 19064 6783 19116 6792
rect 19064 6749 19073 6783
rect 19073 6749 19107 6783
rect 19107 6749 19116 6783
rect 19064 6740 19116 6749
rect 19616 6783 19668 6792
rect 19616 6749 19625 6783
rect 19625 6749 19659 6783
rect 19659 6749 19668 6783
rect 19616 6740 19668 6749
rect 19984 6672 20036 6724
rect 17316 6647 17368 6656
rect 17316 6613 17325 6647
rect 17325 6613 17359 6647
rect 17359 6613 17368 6647
rect 17316 6604 17368 6613
rect 17500 6647 17552 6656
rect 17500 6613 17509 6647
rect 17509 6613 17543 6647
rect 17543 6613 17552 6647
rect 17500 6604 17552 6613
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 2504 6400 2556 6452
rect 1676 6375 1728 6384
rect 1676 6341 1685 6375
rect 1685 6341 1719 6375
rect 1719 6341 1728 6375
rect 1676 6332 1728 6341
rect 3148 6443 3200 6452
rect 3148 6409 3157 6443
rect 3157 6409 3191 6443
rect 3191 6409 3200 6443
rect 3148 6400 3200 6409
rect 3792 6400 3844 6452
rect 4252 6400 4304 6452
rect 5448 6400 5500 6452
rect 6000 6400 6052 6452
rect 6828 6443 6880 6452
rect 6828 6409 6837 6443
rect 6837 6409 6871 6443
rect 6871 6409 6880 6443
rect 6828 6400 6880 6409
rect 10140 6400 10192 6452
rect 10876 6400 10928 6452
rect 11796 6400 11848 6452
rect 1400 6239 1452 6248
rect 1400 6205 1409 6239
rect 1409 6205 1443 6239
rect 1443 6205 1452 6239
rect 1400 6196 1452 6205
rect 2872 6196 2924 6248
rect 3608 6196 3660 6248
rect 8024 6264 8076 6316
rect 8116 6307 8168 6316
rect 8116 6273 8125 6307
rect 8125 6273 8159 6307
rect 8159 6273 8168 6307
rect 8116 6264 8168 6273
rect 9036 6264 9088 6316
rect 9588 6375 9640 6384
rect 9588 6341 9597 6375
rect 9597 6341 9631 6375
rect 9631 6341 9640 6375
rect 9588 6332 9640 6341
rect 10140 6264 10192 6316
rect 10324 6264 10376 6316
rect 6460 6196 6512 6248
rect 11704 6307 11756 6316
rect 11704 6273 11713 6307
rect 11713 6273 11747 6307
rect 11747 6273 11756 6307
rect 11704 6264 11756 6273
rect 12808 6375 12860 6384
rect 12808 6341 12817 6375
rect 12817 6341 12851 6375
rect 12851 6341 12860 6375
rect 12808 6332 12860 6341
rect 11888 6196 11940 6248
rect 3240 6103 3292 6112
rect 3240 6069 3249 6103
rect 3249 6069 3283 6103
rect 3283 6069 3292 6103
rect 3240 6060 3292 6069
rect 6552 6060 6604 6112
rect 11704 6060 11756 6112
rect 12716 6307 12768 6316
rect 12716 6273 12725 6307
rect 12725 6273 12759 6307
rect 12759 6273 12768 6307
rect 15660 6400 15712 6452
rect 16488 6400 16540 6452
rect 14740 6332 14792 6384
rect 12716 6264 12768 6273
rect 13636 6307 13688 6316
rect 13636 6273 13645 6307
rect 13645 6273 13679 6307
rect 13679 6273 13688 6307
rect 13636 6264 13688 6273
rect 13728 6307 13780 6316
rect 13728 6273 13737 6307
rect 13737 6273 13771 6307
rect 13771 6273 13780 6307
rect 13728 6264 13780 6273
rect 14556 6264 14608 6316
rect 14924 6307 14976 6316
rect 14924 6273 14933 6307
rect 14933 6273 14967 6307
rect 14967 6273 14976 6307
rect 14924 6264 14976 6273
rect 15660 6264 15712 6316
rect 15476 6196 15528 6248
rect 16120 6307 16172 6316
rect 16120 6273 16129 6307
rect 16129 6273 16163 6307
rect 16163 6273 16172 6307
rect 16120 6264 16172 6273
rect 16212 6307 16264 6316
rect 16212 6273 16221 6307
rect 16221 6273 16255 6307
rect 16255 6273 16264 6307
rect 16212 6264 16264 6273
rect 17500 6400 17552 6452
rect 19616 6400 19668 6452
rect 20720 6400 20772 6452
rect 21548 6443 21600 6452
rect 21548 6409 21557 6443
rect 21557 6409 21591 6443
rect 21591 6409 21600 6443
rect 21548 6400 21600 6409
rect 18788 6332 18840 6384
rect 16672 6307 16724 6316
rect 16672 6273 16681 6307
rect 16681 6273 16715 6307
rect 16715 6273 16724 6307
rect 16672 6264 16724 6273
rect 14648 6171 14700 6180
rect 14648 6137 14657 6171
rect 14657 6137 14691 6171
rect 14691 6137 14700 6171
rect 14648 6128 14700 6137
rect 16396 6196 16448 6248
rect 17500 6196 17552 6248
rect 20812 6196 20864 6248
rect 18052 6128 18104 6180
rect 18972 6128 19024 6180
rect 13084 6060 13136 6112
rect 13268 6103 13320 6112
rect 13268 6069 13277 6103
rect 13277 6069 13311 6103
rect 13311 6069 13320 6103
rect 13268 6060 13320 6069
rect 18788 6060 18840 6112
rect 21364 6307 21416 6316
rect 21364 6273 21373 6307
rect 21373 6273 21407 6307
rect 21407 6273 21416 6307
rect 21364 6264 21416 6273
rect 24676 6264 24728 6316
rect 21088 6239 21140 6248
rect 21088 6205 21097 6239
rect 21097 6205 21131 6239
rect 21131 6205 21140 6239
rect 21088 6196 21140 6205
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 3240 5856 3292 5908
rect 5356 5856 5408 5908
rect 7564 5856 7616 5908
rect 1400 5720 1452 5772
rect 3700 5720 3752 5772
rect 4620 5720 4672 5772
rect 6552 5763 6604 5772
rect 6552 5729 6561 5763
rect 6561 5729 6595 5763
rect 6595 5729 6604 5763
rect 6552 5720 6604 5729
rect 8024 5720 8076 5772
rect 2872 5652 2924 5704
rect 7288 5695 7340 5704
rect 7288 5661 7297 5695
rect 7297 5661 7331 5695
rect 7331 5661 7340 5695
rect 7288 5652 7340 5661
rect 10416 5856 10468 5908
rect 10876 5856 10928 5908
rect 10508 5788 10560 5840
rect 11060 5788 11112 5840
rect 11336 5856 11388 5908
rect 13636 5856 13688 5908
rect 16212 5856 16264 5908
rect 17500 5856 17552 5908
rect 11888 5788 11940 5840
rect 15476 5788 15528 5840
rect 6092 5584 6144 5636
rect 7012 5584 7064 5636
rect 9036 5584 9088 5636
rect 10416 5627 10468 5636
rect 10416 5593 10425 5627
rect 10425 5593 10459 5627
rect 10459 5593 10468 5627
rect 10416 5584 10468 5593
rect 10508 5627 10560 5636
rect 10508 5593 10517 5627
rect 10517 5593 10551 5627
rect 10551 5593 10560 5627
rect 10508 5584 10560 5593
rect 3608 5516 3660 5568
rect 10876 5695 10928 5704
rect 10876 5661 10885 5695
rect 10885 5661 10919 5695
rect 10919 5661 10928 5695
rect 10876 5652 10928 5661
rect 11152 5695 11204 5704
rect 11152 5661 11161 5695
rect 11161 5661 11195 5695
rect 11195 5661 11204 5695
rect 11152 5652 11204 5661
rect 11060 5627 11112 5636
rect 11060 5593 11069 5627
rect 11069 5593 11103 5627
rect 11103 5593 11112 5627
rect 11060 5584 11112 5593
rect 11704 5695 11756 5704
rect 11704 5661 11713 5695
rect 11713 5661 11747 5695
rect 11747 5661 11756 5695
rect 11704 5652 11756 5661
rect 11336 5584 11388 5636
rect 12808 5652 12860 5704
rect 14556 5695 14608 5704
rect 11244 5516 11296 5568
rect 11888 5516 11940 5568
rect 12716 5516 12768 5568
rect 13084 5584 13136 5636
rect 14556 5661 14565 5695
rect 14565 5661 14599 5695
rect 14599 5661 14608 5695
rect 14556 5652 14608 5661
rect 14740 5695 14792 5704
rect 14740 5661 14749 5695
rect 14749 5661 14783 5695
rect 14783 5661 14792 5695
rect 14740 5652 14792 5661
rect 14924 5695 14976 5704
rect 14924 5661 14933 5695
rect 14933 5661 14967 5695
rect 14967 5661 14976 5695
rect 14924 5652 14976 5661
rect 13636 5516 13688 5568
rect 14648 5516 14700 5568
rect 15568 5584 15620 5636
rect 15936 5695 15988 5704
rect 15936 5661 15945 5695
rect 15945 5661 15979 5695
rect 15979 5661 15988 5695
rect 15936 5652 15988 5661
rect 16396 5788 16448 5840
rect 16672 5763 16724 5772
rect 16672 5729 16681 5763
rect 16681 5729 16715 5763
rect 16715 5729 16724 5763
rect 16672 5720 16724 5729
rect 16580 5695 16632 5704
rect 16580 5661 16589 5695
rect 16589 5661 16623 5695
rect 16623 5661 16632 5695
rect 16580 5652 16632 5661
rect 17224 5788 17276 5840
rect 17316 5720 17368 5772
rect 21088 5856 21140 5908
rect 20812 5720 20864 5772
rect 21824 5720 21876 5772
rect 19524 5652 19576 5704
rect 15292 5516 15344 5568
rect 15476 5559 15528 5568
rect 15476 5525 15485 5559
rect 15485 5525 15519 5559
rect 15519 5525 15528 5559
rect 15476 5516 15528 5525
rect 16120 5516 16172 5568
rect 18788 5584 18840 5636
rect 19984 5584 20036 5636
rect 18696 5559 18748 5568
rect 18696 5525 18705 5559
rect 18705 5525 18739 5559
rect 18739 5525 18748 5559
rect 18696 5516 18748 5525
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 5264 5312 5316 5364
rect 3884 5244 3936 5296
rect 3700 5219 3752 5228
rect 3700 5185 3709 5219
rect 3709 5185 3743 5219
rect 3743 5185 3752 5219
rect 3700 5176 3752 5185
rect 2872 5108 2924 5160
rect 6092 5244 6144 5296
rect 10324 5312 10376 5364
rect 11060 5312 11112 5364
rect 9036 5244 9088 5296
rect 9864 5244 9916 5296
rect 12256 5244 12308 5296
rect 14740 5312 14792 5364
rect 15292 5312 15344 5364
rect 15936 5312 15988 5364
rect 16672 5312 16724 5364
rect 19984 5312 20036 5364
rect 15568 5244 15620 5296
rect 8024 5176 8076 5228
rect 8300 5219 8352 5228
rect 8300 5185 8309 5219
rect 8309 5185 8343 5219
rect 8343 5185 8352 5219
rect 8300 5176 8352 5185
rect 11336 5176 11388 5228
rect 11704 5219 11756 5228
rect 11704 5185 11713 5219
rect 11713 5185 11747 5219
rect 11747 5185 11756 5219
rect 11704 5176 11756 5185
rect 12624 5176 12676 5228
rect 13084 5219 13136 5228
rect 13084 5185 13093 5219
rect 13093 5185 13127 5219
rect 13127 5185 13136 5219
rect 13084 5176 13136 5185
rect 11888 5151 11940 5160
rect 11888 5117 11897 5151
rect 11897 5117 11931 5151
rect 11931 5117 11940 5151
rect 11888 5108 11940 5117
rect 12992 5108 13044 5160
rect 13636 5176 13688 5228
rect 15660 5219 15712 5228
rect 15660 5185 15669 5219
rect 15669 5185 15703 5219
rect 15703 5185 15712 5219
rect 15660 5176 15712 5185
rect 16580 5244 16632 5296
rect 21548 5176 21600 5228
rect 14924 5108 14976 5160
rect 11244 5040 11296 5092
rect 13636 5040 13688 5092
rect 13912 5040 13964 5092
rect 7104 4972 7156 5024
rect 12900 4972 12952 5024
rect 13360 4972 13412 5024
rect 13820 5015 13872 5024
rect 13820 4981 13829 5015
rect 13829 4981 13863 5015
rect 13863 4981 13872 5015
rect 13820 4972 13872 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 13268 4632 13320 4684
rect 12900 4607 12952 4616
rect 12900 4573 12909 4607
rect 12909 4573 12943 4607
rect 12943 4573 12952 4607
rect 12900 4564 12952 4573
rect 15108 4428 15160 4480
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 15292 4267 15344 4276
rect 15292 4233 15301 4267
rect 15301 4233 15335 4267
rect 15335 4233 15344 4267
rect 15292 4224 15344 4233
rect 15108 4156 15160 4208
rect 13360 4131 13412 4140
rect 13360 4097 13369 4131
rect 13369 4097 13403 4131
rect 13403 4097 13412 4131
rect 13360 4088 13412 4097
rect 13728 4088 13780 4140
rect 13912 4088 13964 4140
rect 14924 4131 14976 4140
rect 14924 4097 14933 4131
rect 14933 4097 14967 4131
rect 14967 4097 14976 4131
rect 14924 4088 14976 4097
rect 14188 4063 14240 4072
rect 14188 4029 14197 4063
rect 14197 4029 14231 4063
rect 14231 4029 14240 4063
rect 14188 4020 14240 4029
rect 15200 3884 15252 3936
rect 18696 4088 18748 4140
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 14188 3680 14240 3732
rect 14924 3680 14976 3732
rect 24676 3723 24728 3732
rect 24676 3689 24685 3723
rect 24685 3689 24719 3723
rect 24719 3689 24728 3723
rect 24676 3680 24728 3689
rect 13912 3544 13964 3596
rect 13820 3476 13872 3528
rect 15108 3544 15160 3596
rect 15200 3476 15252 3528
rect 24860 3519 24912 3528
rect 24860 3485 24869 3519
rect 24869 3485 24903 3519
rect 24903 3485 24912 3519
rect 24860 3476 24912 3485
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
<< metal2 >>
rect 9034 27826 9090 28469
rect 9678 27826 9734 28469
rect 10322 27826 10378 28469
rect 10966 27826 11022 28469
rect 9034 27798 9260 27826
rect 9034 27669 9090 27798
rect 4874 26140 5182 26149
rect 4874 26138 4880 26140
rect 4936 26138 4960 26140
rect 5016 26138 5040 26140
rect 5096 26138 5120 26140
rect 5176 26138 5182 26140
rect 4936 26086 4938 26138
rect 5118 26086 5120 26138
rect 4874 26084 4880 26086
rect 4936 26084 4960 26086
rect 5016 26084 5040 26086
rect 5096 26084 5120 26086
rect 5176 26084 5182 26086
rect 4874 26075 5182 26084
rect 9232 25974 9260 27798
rect 9678 27798 9904 27826
rect 9678 27669 9734 27798
rect 9876 25974 9904 27798
rect 10322 27798 10548 27826
rect 10322 27669 10378 27798
rect 10520 25974 10548 27798
rect 10888 27798 11022 27826
rect 9220 25968 9272 25974
rect 9220 25910 9272 25916
rect 9864 25968 9916 25974
rect 9864 25910 9916 25916
rect 10508 25968 10560 25974
rect 10508 25910 10560 25916
rect 10888 25906 10916 27798
rect 10966 27669 11022 27798
rect 11610 27826 11666 28469
rect 12254 27826 12310 28469
rect 12898 27826 12954 28469
rect 13542 27826 13598 28469
rect 14186 27826 14242 28469
rect 14830 27826 14886 28469
rect 15474 27826 15530 28469
rect 16118 27826 16174 28469
rect 17406 27826 17462 28469
rect 18050 27826 18106 28469
rect 11610 27798 11744 27826
rect 11610 27669 11666 27798
rect 11716 25906 11744 27798
rect 12254 27798 12388 27826
rect 12254 27669 12310 27798
rect 12360 25974 12388 27798
rect 12898 27798 13032 27826
rect 12898 27669 12954 27798
rect 12348 25968 12400 25974
rect 12348 25910 12400 25916
rect 13004 25906 13032 27798
rect 13542 27798 13768 27826
rect 13542 27669 13598 27798
rect 13740 25974 13768 27798
rect 14186 27798 14412 27826
rect 14186 27669 14242 27798
rect 14384 25974 14412 27798
rect 14830 27798 15056 27826
rect 14830 27669 14886 27798
rect 15028 25974 15056 27798
rect 15474 27798 15608 27826
rect 15474 27669 15530 27798
rect 13728 25968 13780 25974
rect 13728 25910 13780 25916
rect 14372 25968 14424 25974
rect 14372 25910 14424 25916
rect 15016 25968 15068 25974
rect 15016 25910 15068 25916
rect 15580 25906 15608 27798
rect 16118 27798 16252 27826
rect 16118 27669 16174 27798
rect 16224 25906 16252 27798
rect 17406 27798 17632 27826
rect 17406 27669 17462 27798
rect 17604 25974 17632 27798
rect 18050 27798 18276 27826
rect 18050 27669 18106 27798
rect 18248 25974 18276 27798
rect 17592 25968 17644 25974
rect 17592 25910 17644 25916
rect 18236 25968 18288 25974
rect 18236 25910 18288 25916
rect 4712 25900 4764 25906
rect 4712 25842 4764 25848
rect 10876 25900 10928 25906
rect 10876 25842 10928 25848
rect 11704 25900 11756 25906
rect 11704 25842 11756 25848
rect 12992 25900 13044 25906
rect 12992 25842 13044 25848
rect 15568 25900 15620 25906
rect 15568 25842 15620 25848
rect 16212 25900 16264 25906
rect 16212 25842 16264 25848
rect 4620 25832 4672 25838
rect 4620 25774 4672 25780
rect 2044 25696 2096 25702
rect 2044 25638 2096 25644
rect 2056 25362 2084 25638
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4632 25498 4660 25774
rect 4724 25498 4752 25842
rect 10600 25832 10652 25838
rect 10600 25774 10652 25780
rect 17500 25832 17552 25838
rect 17500 25774 17552 25780
rect 4804 25696 4856 25702
rect 4804 25638 4856 25644
rect 9312 25696 9364 25702
rect 9312 25638 9364 25644
rect 10140 25696 10192 25702
rect 10140 25638 10192 25644
rect 4620 25492 4672 25498
rect 4620 25434 4672 25440
rect 4712 25492 4764 25498
rect 4712 25434 4764 25440
rect 2044 25356 2096 25362
rect 2044 25298 2096 25304
rect 3700 25356 3752 25362
rect 3700 25298 3752 25304
rect 1400 25288 1452 25294
rect 1400 25230 1452 25236
rect 1412 24750 1440 25230
rect 1400 24744 1452 24750
rect 1400 24686 1452 24692
rect 1768 24744 1820 24750
rect 1768 24686 1820 24692
rect 110 24304 166 24313
rect 110 24239 166 24248
rect 124 15162 152 24239
rect 1412 23118 1440 24686
rect 1780 24342 1808 24686
rect 1768 24336 1820 24342
rect 1768 24278 1820 24284
rect 1780 23866 1808 24278
rect 2056 24138 2084 25298
rect 3056 25220 3108 25226
rect 3056 25162 3108 25168
rect 3068 24954 3096 25162
rect 3056 24948 3108 24954
rect 3056 24890 3108 24896
rect 2044 24132 2096 24138
rect 2044 24074 2096 24080
rect 2780 24064 2832 24070
rect 2780 24006 2832 24012
rect 2872 24064 2924 24070
rect 2872 24006 2924 24012
rect 1768 23860 1820 23866
rect 1768 23802 1820 23808
rect 2412 23520 2464 23526
rect 2412 23462 2464 23468
rect 1400 23112 1452 23118
rect 1400 23054 1452 23060
rect 1412 22574 1440 23054
rect 2424 22710 2452 23462
rect 2792 23254 2820 24006
rect 2884 23730 2912 24006
rect 2872 23724 2924 23730
rect 2872 23666 2924 23672
rect 2780 23248 2832 23254
rect 2780 23190 2832 23196
rect 2780 23112 2832 23118
rect 2780 23054 2832 23060
rect 2412 22704 2464 22710
rect 2412 22646 2464 22652
rect 1400 22568 1452 22574
rect 1400 22510 1452 22516
rect 1412 21010 1440 22510
rect 2792 21078 2820 23054
rect 2964 23044 3016 23050
rect 2964 22986 3016 22992
rect 2976 21350 3004 22986
rect 3068 22692 3096 24890
rect 3332 24608 3384 24614
rect 3332 24550 3384 24556
rect 3240 24200 3292 24206
rect 3240 24142 3292 24148
rect 3252 23866 3280 24142
rect 3240 23860 3292 23866
rect 3240 23802 3292 23808
rect 3344 23798 3372 24550
rect 3712 24274 3740 25298
rect 4816 25294 4844 25638
rect 4160 25288 4212 25294
rect 4160 25230 4212 25236
rect 4712 25288 4764 25294
rect 4712 25230 4764 25236
rect 4804 25288 4856 25294
rect 4804 25230 4856 25236
rect 6000 25288 6052 25294
rect 8484 25288 8536 25294
rect 6000 25230 6052 25236
rect 8312 25236 8484 25242
rect 8312 25230 8536 25236
rect 4172 24834 4200 25230
rect 4080 24806 4200 24834
rect 3884 24744 3936 24750
rect 3884 24686 3936 24692
rect 3896 24410 3924 24686
rect 3884 24404 3936 24410
rect 3884 24346 3936 24352
rect 3700 24268 3752 24274
rect 3700 24210 3752 24216
rect 3424 24200 3476 24206
rect 3424 24142 3476 24148
rect 3608 24200 3660 24206
rect 3608 24142 3660 24148
rect 3332 23792 3384 23798
rect 3332 23734 3384 23740
rect 3436 23662 3464 24142
rect 3620 24070 3648 24142
rect 3608 24064 3660 24070
rect 3608 24006 3660 24012
rect 3424 23656 3476 23662
rect 3424 23598 3476 23604
rect 3516 23044 3568 23050
rect 3516 22986 3568 22992
rect 3148 22704 3200 22710
rect 3068 22664 3148 22692
rect 3148 22646 3200 22652
rect 2964 21344 3016 21350
rect 2964 21286 3016 21292
rect 2780 21072 2832 21078
rect 2780 21014 2832 21020
rect 1400 21004 1452 21010
rect 1400 20946 1452 20952
rect 1412 19922 1440 20946
rect 1676 20868 1728 20874
rect 1676 20810 1728 20816
rect 1688 20602 1716 20810
rect 1676 20596 1728 20602
rect 1676 20538 1728 20544
rect 2976 20534 3004 21286
rect 3056 20936 3108 20942
rect 3056 20878 3108 20884
rect 2964 20528 3016 20534
rect 2964 20470 3016 20476
rect 2780 20460 2832 20466
rect 2780 20402 2832 20408
rect 2872 20460 2924 20466
rect 2872 20402 2924 20408
rect 2688 20392 2740 20398
rect 2688 20334 2740 20340
rect 2700 19922 2728 20334
rect 2792 19990 2820 20402
rect 2780 19984 2832 19990
rect 2780 19926 2832 19932
rect 1400 19916 1452 19922
rect 1400 19858 1452 19864
rect 2688 19916 2740 19922
rect 2688 19858 2740 19864
rect 2228 19236 2280 19242
rect 2228 19178 2280 19184
rect 2240 18698 2268 19178
rect 2228 18692 2280 18698
rect 2228 18634 2280 18640
rect 2700 18170 2728 19858
rect 2792 19514 2820 19926
rect 2884 19514 2912 20402
rect 2780 19508 2832 19514
rect 2780 19450 2832 19456
rect 2872 19508 2924 19514
rect 2872 19450 2924 19456
rect 3068 18766 3096 20878
rect 3240 20800 3292 20806
rect 3240 20742 3292 20748
rect 3252 20534 3280 20742
rect 3240 20528 3292 20534
rect 3240 20470 3292 20476
rect 3424 19984 3476 19990
rect 3424 19926 3476 19932
rect 3436 19854 3464 19926
rect 3332 19848 3384 19854
rect 3332 19790 3384 19796
rect 3424 19848 3476 19854
rect 3424 19790 3476 19796
rect 3148 19712 3200 19718
rect 3148 19654 3200 19660
rect 3160 19514 3188 19654
rect 3148 19508 3200 19514
rect 3148 19450 3200 19456
rect 3160 19394 3188 19450
rect 3160 19366 3280 19394
rect 3148 19304 3200 19310
rect 3148 19246 3200 19252
rect 3160 18970 3188 19246
rect 3252 19242 3280 19366
rect 3240 19236 3292 19242
rect 3240 19178 3292 19184
rect 3148 18964 3200 18970
rect 3148 18906 3200 18912
rect 3344 18902 3372 19790
rect 3424 19440 3476 19446
rect 3424 19382 3476 19388
rect 3332 18896 3384 18902
rect 3332 18838 3384 18844
rect 3056 18760 3108 18766
rect 3056 18702 3108 18708
rect 3148 18760 3200 18766
rect 3148 18702 3200 18708
rect 3240 18760 3292 18766
rect 3240 18702 3292 18708
rect 3160 18426 3188 18702
rect 3148 18420 3200 18426
rect 3148 18362 3200 18368
rect 3252 18290 3280 18702
rect 2872 18284 2924 18290
rect 2872 18226 2924 18232
rect 3240 18284 3292 18290
rect 3240 18226 3292 18232
rect 2780 18216 2832 18222
rect 2700 18164 2780 18170
rect 2700 18158 2832 18164
rect 2700 18142 2820 18158
rect 2700 17746 2728 18142
rect 1400 17740 1452 17746
rect 1400 17682 1452 17688
rect 2688 17740 2740 17746
rect 2688 17682 2740 17688
rect 1412 16658 1440 17682
rect 1860 17672 1912 17678
rect 1860 17614 1912 17620
rect 1872 17134 1900 17614
rect 2884 17338 2912 18226
rect 3344 17610 3372 18838
rect 3436 18086 3464 19382
rect 3424 18080 3476 18086
rect 3424 18022 3476 18028
rect 3332 17604 3384 17610
rect 3332 17546 3384 17552
rect 2872 17332 2924 17338
rect 2872 17274 2924 17280
rect 1860 17128 1912 17134
rect 1860 17070 1912 17076
rect 1768 16992 1820 16998
rect 1768 16934 1820 16940
rect 1780 16658 1808 16934
rect 1400 16652 1452 16658
rect 1400 16594 1452 16600
rect 1768 16652 1820 16658
rect 1768 16594 1820 16600
rect 1412 15638 1440 16594
rect 1400 15632 1452 15638
rect 1400 15574 1452 15580
rect 1400 15496 1452 15502
rect 1400 15438 1452 15444
rect 112 15156 164 15162
rect 112 15098 164 15104
rect 1412 15065 1440 15438
rect 1398 15056 1454 15065
rect 1398 14991 1454 15000
rect 1768 14816 1820 14822
rect 1768 14758 1820 14764
rect 1780 14482 1808 14758
rect 1768 14476 1820 14482
rect 1768 14418 1820 14424
rect 1676 14408 1728 14414
rect 1872 14362 1900 17070
rect 2884 16794 2912 17274
rect 3344 17270 3372 17546
rect 3436 17338 3464 18022
rect 3424 17332 3476 17338
rect 3424 17274 3476 17280
rect 3332 17264 3384 17270
rect 3528 17218 3556 22986
rect 3620 22982 3648 24006
rect 3712 23730 3740 24210
rect 3884 24200 3936 24206
rect 3884 24142 3936 24148
rect 3896 23730 3924 24142
rect 4080 24070 4108 24806
rect 4528 24744 4580 24750
rect 4580 24704 4660 24732
rect 4528 24686 4580 24692
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4252 24404 4304 24410
rect 4252 24346 4304 24352
rect 4344 24404 4396 24410
rect 4344 24346 4396 24352
rect 4160 24200 4212 24206
rect 4160 24142 4212 24148
rect 4068 24064 4120 24070
rect 4068 24006 4120 24012
rect 4172 23730 4200 24142
rect 3700 23724 3752 23730
rect 3700 23666 3752 23672
rect 3884 23724 3936 23730
rect 3884 23666 3936 23672
rect 4160 23724 4212 23730
rect 4160 23666 4212 23672
rect 3896 23322 3924 23666
rect 4172 23508 4200 23666
rect 4264 23662 4292 24346
rect 4252 23656 4304 23662
rect 4252 23598 4304 23604
rect 4356 23526 4384 24346
rect 4632 24342 4660 24704
rect 4620 24336 4672 24342
rect 4620 24278 4672 24284
rect 4724 24070 4752 25230
rect 5356 25220 5408 25226
rect 5356 25162 5408 25168
rect 4804 25152 4856 25158
rect 4804 25094 4856 25100
rect 5264 25152 5316 25158
rect 5264 25094 5316 25100
rect 4816 24410 4844 25094
rect 4874 25052 5182 25061
rect 4874 25050 4880 25052
rect 4936 25050 4960 25052
rect 5016 25050 5040 25052
rect 5096 25050 5120 25052
rect 5176 25050 5182 25052
rect 4936 24998 4938 25050
rect 5118 24998 5120 25050
rect 4874 24996 4880 24998
rect 4936 24996 4960 24998
rect 5016 24996 5040 24998
rect 5096 24996 5120 24998
rect 5176 24996 5182 24998
rect 4874 24987 5182 24996
rect 4804 24404 4856 24410
rect 4804 24346 4856 24352
rect 5276 24206 5304 25094
rect 4804 24200 4856 24206
rect 4804 24142 4856 24148
rect 5264 24200 5316 24206
rect 5264 24142 5316 24148
rect 4528 24064 4580 24070
rect 4528 24006 4580 24012
rect 4712 24064 4764 24070
rect 4712 24006 4764 24012
rect 4540 23798 4568 24006
rect 4528 23792 4580 23798
rect 4528 23734 4580 23740
rect 4620 23656 4672 23662
rect 4620 23598 4672 23604
rect 4080 23480 4200 23508
rect 4344 23520 4396 23526
rect 3884 23316 3936 23322
rect 4080 23304 4108 23480
rect 4344 23462 4396 23468
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4080 23276 4200 23304
rect 3884 23258 3936 23264
rect 3608 22976 3660 22982
rect 3608 22918 3660 22924
rect 3896 22778 3924 23258
rect 4172 23118 4200 23276
rect 4632 23118 4660 23598
rect 4724 23526 4752 24006
rect 4816 23594 4844 24142
rect 5264 24064 5316 24070
rect 5264 24006 5316 24012
rect 4874 23964 5182 23973
rect 4874 23962 4880 23964
rect 4936 23962 4960 23964
rect 5016 23962 5040 23964
rect 5096 23962 5120 23964
rect 5176 23962 5182 23964
rect 4936 23910 4938 23962
rect 5118 23910 5120 23962
rect 4874 23908 4880 23910
rect 4936 23908 4960 23910
rect 5016 23908 5040 23910
rect 5096 23908 5120 23910
rect 5176 23908 5182 23910
rect 4874 23899 5182 23908
rect 5172 23724 5224 23730
rect 5172 23666 5224 23672
rect 4804 23588 4856 23594
rect 4804 23530 4856 23536
rect 4712 23520 4764 23526
rect 4712 23462 4764 23468
rect 5184 23508 5212 23666
rect 5276 23662 5304 24006
rect 5264 23656 5316 23662
rect 5264 23598 5316 23604
rect 5368 23508 5396 25162
rect 6012 24954 6040 25230
rect 7380 25220 7432 25226
rect 7380 25162 7432 25168
rect 8312 25214 8524 25230
rect 6000 24948 6052 24954
rect 6000 24890 6052 24896
rect 6012 23730 6040 24890
rect 7196 24608 7248 24614
rect 7196 24550 7248 24556
rect 7208 24410 7236 24550
rect 7196 24404 7248 24410
rect 7196 24346 7248 24352
rect 6184 24132 6236 24138
rect 6184 24074 6236 24080
rect 6000 23724 6052 23730
rect 6000 23666 6052 23672
rect 6092 23656 6144 23662
rect 6092 23598 6144 23604
rect 5184 23480 5396 23508
rect 5184 23322 5212 23480
rect 5172 23316 5224 23322
rect 5172 23258 5224 23264
rect 4160 23112 4212 23118
rect 4160 23054 4212 23060
rect 4620 23112 4672 23118
rect 4620 23054 4672 23060
rect 4874 22876 5182 22885
rect 4874 22874 4880 22876
rect 4936 22874 4960 22876
rect 5016 22874 5040 22876
rect 5096 22874 5120 22876
rect 5176 22874 5182 22876
rect 4936 22822 4938 22874
rect 5118 22822 5120 22874
rect 4874 22820 4880 22822
rect 4936 22820 4960 22822
rect 5016 22820 5040 22822
rect 5096 22820 5120 22822
rect 5176 22820 5182 22822
rect 4874 22811 5182 22820
rect 3884 22772 3936 22778
rect 3884 22714 3936 22720
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 3608 22024 3660 22030
rect 3608 21966 3660 21972
rect 6000 22024 6052 22030
rect 6000 21966 6052 21972
rect 3620 20942 3648 21966
rect 5816 21956 5868 21962
rect 5816 21898 5868 21904
rect 5632 21888 5684 21894
rect 5632 21830 5684 21836
rect 4874 21788 5182 21797
rect 4874 21786 4880 21788
rect 4936 21786 4960 21788
rect 5016 21786 5040 21788
rect 5096 21786 5120 21788
rect 5176 21786 5182 21788
rect 4936 21734 4938 21786
rect 5118 21734 5120 21786
rect 4874 21732 4880 21734
rect 4936 21732 4960 21734
rect 5016 21732 5040 21734
rect 5096 21732 5120 21734
rect 5176 21732 5182 21734
rect 4874 21723 5182 21732
rect 4988 21684 5040 21690
rect 4988 21626 5040 21632
rect 4160 21616 4212 21622
rect 4160 21558 4212 21564
rect 4172 21434 4200 21558
rect 4620 21548 4672 21554
rect 4620 21490 4672 21496
rect 4080 21406 4200 21434
rect 4080 21026 4108 21406
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4528 21072 4580 21078
rect 4080 20998 4200 21026
rect 4528 21014 4580 21020
rect 4172 20942 4200 20998
rect 3608 20936 3660 20942
rect 3608 20878 3660 20884
rect 4160 20936 4212 20942
rect 4160 20878 4212 20884
rect 3620 20806 3648 20878
rect 4068 20868 4120 20874
rect 4068 20810 4120 20816
rect 3608 20800 3660 20806
rect 3608 20742 3660 20748
rect 3620 20602 3648 20742
rect 4080 20602 4108 20810
rect 3608 20596 3660 20602
rect 3608 20538 3660 20544
rect 4068 20596 4120 20602
rect 4068 20538 4120 20544
rect 4172 20346 4200 20878
rect 4540 20806 4568 21014
rect 4632 20942 4660 21490
rect 4712 21412 4764 21418
rect 4712 21354 4764 21360
rect 4724 21010 4752 21354
rect 5000 21146 5028 21626
rect 5644 21554 5672 21830
rect 5632 21548 5684 21554
rect 5632 21490 5684 21496
rect 5828 21486 5856 21898
rect 6012 21554 6040 21966
rect 6104 21622 6132 23598
rect 6196 22710 6224 24074
rect 6920 24064 6972 24070
rect 6920 24006 6972 24012
rect 6932 23798 6960 24006
rect 7208 23866 7236 24346
rect 7392 24070 7420 25162
rect 7564 25152 7616 25158
rect 7564 25094 7616 25100
rect 7470 24440 7526 24449
rect 7470 24375 7526 24384
rect 7484 24138 7512 24375
rect 7576 24138 7604 25094
rect 8312 24834 8340 25214
rect 8392 25152 8444 25158
rect 8392 25094 8444 25100
rect 8128 24806 8340 24834
rect 8128 24342 8156 24806
rect 8208 24744 8260 24750
rect 8206 24712 8208 24721
rect 8260 24712 8262 24721
rect 8404 24698 8432 25094
rect 8496 24818 8524 25214
rect 9220 25220 9272 25226
rect 9220 25162 9272 25168
rect 8576 25152 8628 25158
rect 8576 25094 8628 25100
rect 8484 24812 8536 24818
rect 8484 24754 8536 24760
rect 8404 24670 8524 24698
rect 8206 24647 8262 24656
rect 8116 24336 8168 24342
rect 8116 24278 8168 24284
rect 7840 24200 7892 24206
rect 7840 24142 7892 24148
rect 7472 24132 7524 24138
rect 7472 24074 7524 24080
rect 7564 24132 7616 24138
rect 7564 24074 7616 24080
rect 7380 24064 7432 24070
rect 7380 24006 7432 24012
rect 7196 23860 7248 23866
rect 7196 23802 7248 23808
rect 6920 23792 6972 23798
rect 6920 23734 6972 23740
rect 7104 23724 7156 23730
rect 7104 23666 7156 23672
rect 7116 23186 7144 23666
rect 7392 23662 7420 24006
rect 7576 23848 7604 24074
rect 7576 23820 7696 23848
rect 7668 23662 7696 23820
rect 7380 23656 7432 23662
rect 7380 23598 7432 23604
rect 7656 23656 7708 23662
rect 7656 23598 7708 23604
rect 7852 23594 7880 24142
rect 7840 23588 7892 23594
rect 7840 23530 7892 23536
rect 7288 23520 7340 23526
rect 7288 23462 7340 23468
rect 7380 23520 7432 23526
rect 7380 23462 7432 23468
rect 7300 23322 7328 23462
rect 7288 23316 7340 23322
rect 7288 23258 7340 23264
rect 7104 23180 7156 23186
rect 7104 23122 7156 23128
rect 7116 22778 7144 23122
rect 7392 23118 7420 23462
rect 7380 23112 7432 23118
rect 7380 23054 7432 23060
rect 7104 22772 7156 22778
rect 7104 22714 7156 22720
rect 6184 22704 6236 22710
rect 6184 22646 6236 22652
rect 6092 21616 6144 21622
rect 6092 21558 6144 21564
rect 6000 21548 6052 21554
rect 6000 21490 6052 21496
rect 5816 21480 5868 21486
rect 5816 21422 5868 21428
rect 4988 21140 5040 21146
rect 4988 21082 5040 21088
rect 4712 21004 4764 21010
rect 4712 20946 4764 20952
rect 4620 20936 4672 20942
rect 4620 20878 4672 20884
rect 4528 20800 4580 20806
rect 4528 20742 4580 20748
rect 4540 20534 4568 20742
rect 4528 20528 4580 20534
rect 4528 20470 4580 20476
rect 4632 20466 4660 20878
rect 4620 20460 4672 20466
rect 4620 20402 4672 20408
rect 4724 20346 4752 20946
rect 6196 20874 6224 22646
rect 6368 22024 6420 22030
rect 6552 22024 6604 22030
rect 6420 21984 6552 22012
rect 6368 21966 6420 21972
rect 6552 21966 6604 21972
rect 6460 21480 6512 21486
rect 6460 21422 6512 21428
rect 6368 21004 6420 21010
rect 6368 20946 6420 20952
rect 6184 20868 6236 20874
rect 6184 20810 6236 20816
rect 4804 20800 4856 20806
rect 4804 20742 4856 20748
rect 4080 20318 4200 20346
rect 4632 20330 4752 20346
rect 4620 20324 4752 20330
rect 3608 20256 3660 20262
rect 3608 20198 3660 20204
rect 3620 19854 3648 20198
rect 3608 19848 3660 19854
rect 3608 19790 3660 19796
rect 3620 18834 3648 19790
rect 4080 19718 4108 20318
rect 4672 20318 4752 20324
rect 4620 20266 4672 20272
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4160 19848 4212 19854
rect 4160 19790 4212 19796
rect 4068 19712 4120 19718
rect 4068 19654 4120 19660
rect 4172 19242 4200 19790
rect 4712 19780 4764 19786
rect 4712 19722 4764 19728
rect 4160 19236 4212 19242
rect 4160 19178 4212 19184
rect 4620 19236 4672 19242
rect 4620 19178 4672 19184
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 3608 18828 3660 18834
rect 3608 18770 3660 18776
rect 3700 18624 3752 18630
rect 3700 18566 3752 18572
rect 3712 18358 3740 18566
rect 3700 18352 3752 18358
rect 3700 18294 3752 18300
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4160 17536 4212 17542
rect 4160 17478 4212 17484
rect 3332 17206 3384 17212
rect 2964 17128 3016 17134
rect 2964 17070 3016 17076
rect 2872 16788 2924 16794
rect 2872 16730 2924 16736
rect 2884 16266 2912 16730
rect 2792 16238 2912 16266
rect 2792 16046 2820 16238
rect 2872 16176 2924 16182
rect 2872 16118 2924 16124
rect 2780 16040 2832 16046
rect 2780 15982 2832 15988
rect 2044 15904 2096 15910
rect 2044 15846 2096 15852
rect 2056 15502 2084 15846
rect 2596 15564 2648 15570
rect 2596 15506 2648 15512
rect 2044 15496 2096 15502
rect 2044 15438 2096 15444
rect 2608 15094 2636 15506
rect 2884 15502 2912 16118
rect 2976 16046 3004 17070
rect 3344 16522 3372 17206
rect 3436 17190 3556 17218
rect 4172 17202 4200 17478
rect 4632 17202 4660 19178
rect 4160 17196 4212 17202
rect 3436 17134 3464 17190
rect 4160 17138 4212 17144
rect 4620 17196 4672 17202
rect 4620 17138 4672 17144
rect 3424 17128 3476 17134
rect 3424 17070 3476 17076
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4632 16658 4660 17138
rect 4620 16652 4672 16658
rect 4620 16594 4672 16600
rect 3332 16516 3384 16522
rect 3332 16458 3384 16464
rect 2964 16040 3016 16046
rect 2964 15982 3016 15988
rect 3148 16040 3200 16046
rect 3148 15982 3200 15988
rect 2872 15496 2924 15502
rect 2872 15438 2924 15444
rect 2596 15088 2648 15094
rect 2596 15030 2648 15036
rect 2884 15026 2912 15438
rect 2964 15360 3016 15366
rect 2964 15302 3016 15308
rect 2780 15020 2832 15026
rect 2780 14962 2832 14968
rect 2872 15020 2924 15026
rect 2872 14962 2924 14968
rect 2792 14618 2820 14962
rect 2780 14612 2832 14618
rect 2780 14554 2832 14560
rect 1676 14350 1728 14356
rect 846 14240 902 14249
rect 846 14175 902 14184
rect 860 13938 888 14175
rect 1688 13938 1716 14350
rect 1780 14334 1900 14362
rect 1780 14074 1808 14334
rect 1768 14068 1820 14074
rect 1768 14010 1820 14016
rect 848 13932 900 13938
rect 848 13874 900 13880
rect 1676 13932 1728 13938
rect 1676 13874 1728 13880
rect 1676 12164 1728 12170
rect 1676 12106 1728 12112
rect 1688 11898 1716 12106
rect 1676 11892 1728 11898
rect 1676 11834 1728 11840
rect 1676 11756 1728 11762
rect 1676 11698 1728 11704
rect 848 11552 900 11558
rect 846 11520 848 11529
rect 1584 11552 1636 11558
rect 900 11520 902 11529
rect 1584 11494 1636 11500
rect 846 11455 902 11464
rect 1596 11150 1624 11494
rect 1688 11354 1716 11698
rect 1676 11348 1728 11354
rect 1676 11290 1728 11296
rect 1584 11144 1636 11150
rect 1584 11086 1636 11092
rect 1780 10130 1808 14010
rect 2320 13864 2372 13870
rect 2320 13806 2372 13812
rect 2332 13530 2360 13806
rect 2320 13524 2372 13530
rect 2320 13466 2372 13472
rect 2320 12708 2372 12714
rect 2320 12650 2372 12656
rect 2332 11762 2360 12650
rect 2320 11756 2372 11762
rect 2320 11698 2372 11704
rect 2780 10668 2832 10674
rect 2780 10610 2832 10616
rect 1768 10124 1820 10130
rect 1768 10066 1820 10072
rect 2136 9920 2188 9926
rect 2136 9862 2188 9868
rect 2148 6866 2176 9862
rect 2792 9654 2820 10610
rect 2976 10198 3004 15302
rect 3160 14958 3188 15982
rect 3344 15434 3372 16458
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4632 15570 4660 16594
rect 4724 15638 4752 19722
rect 4816 18970 4844 20742
rect 4874 20700 5182 20709
rect 4874 20698 4880 20700
rect 4936 20698 4960 20700
rect 5016 20698 5040 20700
rect 5096 20698 5120 20700
rect 5176 20698 5182 20700
rect 4936 20646 4938 20698
rect 5118 20646 5120 20698
rect 4874 20644 4880 20646
rect 4936 20644 4960 20646
rect 5016 20644 5040 20646
rect 5096 20644 5120 20646
rect 5176 20644 5182 20646
rect 4874 20635 5182 20644
rect 6184 20528 6236 20534
rect 6184 20470 6236 20476
rect 5448 20460 5500 20466
rect 5448 20402 5500 20408
rect 5356 20324 5408 20330
rect 5356 20266 5408 20272
rect 5264 20256 5316 20262
rect 5264 20198 5316 20204
rect 5276 19786 5304 20198
rect 5368 19854 5396 20266
rect 5460 19922 5488 20402
rect 5448 19916 5500 19922
rect 5448 19858 5500 19864
rect 5356 19848 5408 19854
rect 5356 19790 5408 19796
rect 5264 19780 5316 19786
rect 5264 19722 5316 19728
rect 4874 19612 5182 19621
rect 4874 19610 4880 19612
rect 4936 19610 4960 19612
rect 5016 19610 5040 19612
rect 5096 19610 5120 19612
rect 5176 19610 5182 19612
rect 4936 19558 4938 19610
rect 5118 19558 5120 19610
rect 4874 19556 4880 19558
rect 4936 19556 4960 19558
rect 5016 19556 5040 19558
rect 5096 19556 5120 19558
rect 5176 19556 5182 19558
rect 4874 19547 5182 19556
rect 5460 19378 5488 19858
rect 5816 19780 5868 19786
rect 5816 19722 5868 19728
rect 5828 19378 5856 19722
rect 6000 19712 6052 19718
rect 6000 19654 6052 19660
rect 6012 19378 6040 19654
rect 6196 19378 6224 20470
rect 6380 19922 6408 20946
rect 6472 20874 6500 21422
rect 6564 21418 6592 21966
rect 6920 21888 6972 21894
rect 6920 21830 6972 21836
rect 6932 21554 6960 21830
rect 6920 21548 6972 21554
rect 6920 21490 6972 21496
rect 6552 21412 6604 21418
rect 6552 21354 6604 21360
rect 7288 21344 7340 21350
rect 7288 21286 7340 21292
rect 7300 21078 7328 21286
rect 7288 21072 7340 21078
rect 7288 21014 7340 21020
rect 6460 20868 6512 20874
rect 6460 20810 6512 20816
rect 7392 20534 7420 23054
rect 8128 22642 8156 24278
rect 8220 24274 8248 24647
rect 8496 24614 8524 24670
rect 8392 24608 8444 24614
rect 8392 24550 8444 24556
rect 8484 24608 8536 24614
rect 8484 24550 8536 24556
rect 8404 24410 8432 24550
rect 8588 24410 8616 25094
rect 9232 24954 9260 25162
rect 9220 24948 9272 24954
rect 9220 24890 9272 24896
rect 8760 24880 8812 24886
rect 8760 24822 8812 24828
rect 8668 24812 8720 24818
rect 8668 24754 8720 24760
rect 8300 24404 8352 24410
rect 8300 24346 8352 24352
rect 8392 24404 8444 24410
rect 8392 24346 8444 24352
rect 8576 24404 8628 24410
rect 8576 24346 8628 24352
rect 8208 24268 8260 24274
rect 8208 24210 8260 24216
rect 8116 22636 8168 22642
rect 8116 22578 8168 22584
rect 7656 21548 7708 21554
rect 7656 21490 7708 21496
rect 7380 20528 7432 20534
rect 7380 20470 7432 20476
rect 7104 20392 7156 20398
rect 7104 20334 7156 20340
rect 7116 19922 7144 20334
rect 7392 20330 7420 20470
rect 7668 20466 7696 21490
rect 8024 21480 8076 21486
rect 8024 21422 8076 21428
rect 7656 20460 7708 20466
rect 8036 20448 8064 21422
rect 8128 21010 8156 22578
rect 8312 21146 8340 24346
rect 8680 24274 8708 24754
rect 8772 24682 8800 24822
rect 9220 24812 9272 24818
rect 9220 24754 9272 24760
rect 9034 24712 9090 24721
rect 8760 24676 8812 24682
rect 9034 24647 9090 24656
rect 8760 24618 8812 24624
rect 9048 24614 9076 24647
rect 9036 24608 9088 24614
rect 9036 24550 9088 24556
rect 9232 24342 9260 24754
rect 9220 24336 9272 24342
rect 9220 24278 9272 24284
rect 8668 24268 8720 24274
rect 8668 24210 8720 24216
rect 8392 24200 8444 24206
rect 8392 24142 8444 24148
rect 8404 23730 8432 24142
rect 8392 23724 8444 23730
rect 8392 23666 8444 23672
rect 8404 23254 8432 23666
rect 8392 23248 8444 23254
rect 8392 23190 8444 23196
rect 8680 23118 8708 24210
rect 8760 23588 8812 23594
rect 8760 23530 8812 23536
rect 8668 23112 8720 23118
rect 8668 23054 8720 23060
rect 8392 22976 8444 22982
rect 8392 22918 8444 22924
rect 8404 22574 8432 22918
rect 8392 22568 8444 22574
rect 8392 22510 8444 22516
rect 8392 22160 8444 22166
rect 8392 22102 8444 22108
rect 8404 21554 8432 22102
rect 8680 22098 8708 23054
rect 8772 23050 8800 23530
rect 9036 23520 9088 23526
rect 9036 23462 9088 23468
rect 8760 23044 8812 23050
rect 8760 22986 8812 22992
rect 9048 22642 9076 23462
rect 9324 23050 9352 25638
rect 9956 25220 10008 25226
rect 9956 25162 10008 25168
rect 9404 24812 9456 24818
rect 9404 24754 9456 24760
rect 9416 24449 9444 24754
rect 9968 24682 9996 25162
rect 9956 24676 10008 24682
rect 9956 24618 10008 24624
rect 9402 24440 9458 24449
rect 9402 24375 9458 24384
rect 9588 23316 9640 23322
rect 9588 23258 9640 23264
rect 9312 23044 9364 23050
rect 9312 22986 9364 22992
rect 9496 23044 9548 23050
rect 9496 22986 9548 22992
rect 9128 22976 9180 22982
rect 9128 22918 9180 22924
rect 9140 22642 9168 22918
rect 8760 22636 8812 22642
rect 8760 22578 8812 22584
rect 8852 22636 8904 22642
rect 8852 22578 8904 22584
rect 9036 22636 9088 22642
rect 9036 22578 9088 22584
rect 9128 22636 9180 22642
rect 9128 22578 9180 22584
rect 8668 22092 8720 22098
rect 8668 22034 8720 22040
rect 8576 21888 8628 21894
rect 8576 21830 8628 21836
rect 8588 21554 8616 21830
rect 8392 21548 8444 21554
rect 8392 21490 8444 21496
rect 8576 21548 8628 21554
rect 8576 21490 8628 21496
rect 8300 21140 8352 21146
rect 8300 21082 8352 21088
rect 8116 21004 8168 21010
rect 8116 20946 8168 20952
rect 8576 20936 8628 20942
rect 8576 20878 8628 20884
rect 8300 20868 8352 20874
rect 8300 20810 8352 20816
rect 8208 20528 8260 20534
rect 8208 20470 8260 20476
rect 8036 20420 8156 20448
rect 7656 20402 7708 20408
rect 7380 20324 7432 20330
rect 7380 20266 7432 20272
rect 8128 20262 8156 20420
rect 7656 20256 7708 20262
rect 7656 20198 7708 20204
rect 8116 20256 8168 20262
rect 8116 20198 8168 20204
rect 6368 19916 6420 19922
rect 6368 19858 6420 19864
rect 7104 19916 7156 19922
rect 7288 19916 7340 19922
rect 7156 19876 7236 19904
rect 7104 19858 7156 19864
rect 6380 19378 6408 19858
rect 7104 19780 7156 19786
rect 7104 19722 7156 19728
rect 5448 19372 5500 19378
rect 5448 19314 5500 19320
rect 5816 19372 5868 19378
rect 5816 19314 5868 19320
rect 6000 19372 6052 19378
rect 6000 19314 6052 19320
rect 6184 19372 6236 19378
rect 6184 19314 6236 19320
rect 6368 19372 6420 19378
rect 6368 19314 6420 19320
rect 4804 18964 4856 18970
rect 4804 18906 4856 18912
rect 6092 18964 6144 18970
rect 6092 18906 6144 18912
rect 4804 18828 4856 18834
rect 4804 18770 4856 18776
rect 4816 18698 4844 18770
rect 5356 18760 5408 18766
rect 5356 18702 5408 18708
rect 4804 18692 4856 18698
rect 4804 18634 4856 18640
rect 4816 18340 4844 18634
rect 5264 18624 5316 18630
rect 5264 18566 5316 18572
rect 4874 18524 5182 18533
rect 4874 18522 4880 18524
rect 4936 18522 4960 18524
rect 5016 18522 5040 18524
rect 5096 18522 5120 18524
rect 5176 18522 5182 18524
rect 4936 18470 4938 18522
rect 5118 18470 5120 18522
rect 4874 18468 4880 18470
rect 4936 18468 4960 18470
rect 5016 18468 5040 18470
rect 5096 18468 5120 18470
rect 5176 18468 5182 18470
rect 4874 18459 5182 18468
rect 4988 18352 5040 18358
rect 4816 18312 4988 18340
rect 4988 18294 5040 18300
rect 5276 18086 5304 18566
rect 5368 18426 5396 18702
rect 5356 18420 5408 18426
rect 5356 18362 5408 18368
rect 6104 18290 6132 18906
rect 6380 18834 6408 19314
rect 6828 19236 6880 19242
rect 6828 19178 6880 19184
rect 6840 18834 6868 19178
rect 6368 18828 6420 18834
rect 6368 18770 6420 18776
rect 6828 18828 6880 18834
rect 6828 18770 6880 18776
rect 7116 18630 7144 19722
rect 7208 19514 7236 19876
rect 7288 19858 7340 19864
rect 7300 19718 7328 19858
rect 7288 19712 7340 19718
rect 7288 19654 7340 19660
rect 7472 19712 7524 19718
rect 7472 19654 7524 19660
rect 7196 19508 7248 19514
rect 7196 19450 7248 19456
rect 7380 19168 7432 19174
rect 7380 19110 7432 19116
rect 7104 18624 7156 18630
rect 7104 18566 7156 18572
rect 7116 18358 7144 18566
rect 7392 18426 7420 19110
rect 7380 18420 7432 18426
rect 7380 18362 7432 18368
rect 7484 18358 7512 19654
rect 7668 19242 7696 20198
rect 7932 19848 7984 19854
rect 7932 19790 7984 19796
rect 7656 19236 7708 19242
rect 7656 19178 7708 19184
rect 7564 18964 7616 18970
rect 7668 18952 7696 19178
rect 7616 18924 7696 18952
rect 7564 18906 7616 18912
rect 7944 18358 7972 19790
rect 8128 19718 8156 20198
rect 8220 19786 8248 20470
rect 8208 19780 8260 19786
rect 8208 19722 8260 19728
rect 8116 19712 8168 19718
rect 8116 19654 8168 19660
rect 8312 18902 8340 20810
rect 8392 20528 8444 20534
rect 8392 20470 8444 20476
rect 8404 19990 8432 20470
rect 8588 20398 8616 20878
rect 8680 20534 8708 22034
rect 8772 21350 8800 22578
rect 8864 22001 8892 22578
rect 9220 22568 9272 22574
rect 9220 22510 9272 22516
rect 8944 22432 8996 22438
rect 8944 22374 8996 22380
rect 8956 22234 8984 22374
rect 8944 22228 8996 22234
rect 8944 22170 8996 22176
rect 9232 22098 9260 22510
rect 9324 22438 9352 22986
rect 9508 22778 9536 22986
rect 9496 22772 9548 22778
rect 9496 22714 9548 22720
rect 9600 22642 9628 23258
rect 9772 23248 9824 23254
rect 9772 23190 9824 23196
rect 9680 23044 9732 23050
rect 9680 22986 9732 22992
rect 9692 22710 9720 22986
rect 9680 22704 9732 22710
rect 9680 22646 9732 22652
rect 9784 22642 9812 23190
rect 9864 22976 9916 22982
rect 9864 22918 9916 22924
rect 9404 22636 9456 22642
rect 9404 22578 9456 22584
rect 9588 22636 9640 22642
rect 9588 22578 9640 22584
rect 9772 22636 9824 22642
rect 9772 22578 9824 22584
rect 9312 22432 9364 22438
rect 9312 22374 9364 22380
rect 9220 22092 9272 22098
rect 9220 22034 9272 22040
rect 8850 21992 8906 22001
rect 8850 21927 8906 21936
rect 8760 21344 8812 21350
rect 8760 21286 8812 21292
rect 8668 20528 8720 20534
rect 8668 20470 8720 20476
rect 8576 20392 8628 20398
rect 8576 20334 8628 20340
rect 8392 19984 8444 19990
rect 8392 19926 8444 19932
rect 8300 18896 8352 18902
rect 8300 18838 8352 18844
rect 8116 18692 8168 18698
rect 8116 18634 8168 18640
rect 8128 18426 8156 18634
rect 8404 18630 8432 19926
rect 8668 19712 8720 19718
rect 8772 19700 8800 21286
rect 8720 19672 8800 19700
rect 8668 19654 8720 19660
rect 8668 19304 8720 19310
rect 8668 19246 8720 19252
rect 8392 18624 8444 18630
rect 8392 18566 8444 18572
rect 8116 18420 8168 18426
rect 8116 18362 8168 18368
rect 7104 18352 7156 18358
rect 7104 18294 7156 18300
rect 7472 18352 7524 18358
rect 7472 18294 7524 18300
rect 7932 18352 7984 18358
rect 7932 18294 7984 18300
rect 8680 18290 8708 19246
rect 8772 18766 8800 19672
rect 8864 18766 8892 21927
rect 9416 21690 9444 22578
rect 9404 21684 9456 21690
rect 9404 21626 9456 21632
rect 9600 20942 9628 22578
rect 9770 22536 9826 22545
rect 9770 22471 9826 22480
rect 9680 21888 9732 21894
rect 9680 21830 9732 21836
rect 9692 21146 9720 21830
rect 9784 21486 9812 22471
rect 9876 21962 9904 22918
rect 9968 22658 9996 24618
rect 10048 22976 10100 22982
rect 10048 22918 10100 22924
rect 10060 22778 10088 22918
rect 10048 22772 10100 22778
rect 10048 22714 10100 22720
rect 9968 22630 10088 22658
rect 9956 22228 10008 22234
rect 9956 22170 10008 22176
rect 9968 22098 9996 22170
rect 9956 22092 10008 22098
rect 10060 22094 10088 22630
rect 10152 22545 10180 25638
rect 10508 25152 10560 25158
rect 10508 25094 10560 25100
rect 10232 24608 10284 24614
rect 10232 24550 10284 24556
rect 10138 22536 10194 22545
rect 10138 22471 10194 22480
rect 10060 22066 10180 22094
rect 9956 22034 10008 22040
rect 9864 21956 9916 21962
rect 9864 21898 9916 21904
rect 9772 21480 9824 21486
rect 9772 21422 9824 21428
rect 9876 21418 10088 21434
rect 9864 21412 10100 21418
rect 9916 21406 10048 21412
rect 9864 21354 9916 21360
rect 10048 21354 10100 21360
rect 9680 21140 9732 21146
rect 9680 21082 9732 21088
rect 9864 21004 9916 21010
rect 9864 20946 9916 20952
rect 9588 20936 9640 20942
rect 9588 20878 9640 20884
rect 9312 20256 9364 20262
rect 9312 20198 9364 20204
rect 9324 19786 9352 20198
rect 9772 19848 9824 19854
rect 9772 19790 9824 19796
rect 9312 19780 9364 19786
rect 9312 19722 9364 19728
rect 9324 19514 9352 19722
rect 9680 19712 9732 19718
rect 9680 19654 9732 19660
rect 9312 19508 9364 19514
rect 9312 19450 9364 19456
rect 8944 19372 8996 19378
rect 8944 19314 8996 19320
rect 8760 18760 8812 18766
rect 8760 18702 8812 18708
rect 8852 18760 8904 18766
rect 8852 18702 8904 18708
rect 8772 18426 8800 18702
rect 8760 18420 8812 18426
rect 8760 18362 8812 18368
rect 6092 18284 6144 18290
rect 6092 18226 6144 18232
rect 8668 18284 8720 18290
rect 8668 18226 8720 18232
rect 5264 18080 5316 18086
rect 5264 18022 5316 18028
rect 4874 17436 5182 17445
rect 4874 17434 4880 17436
rect 4936 17434 4960 17436
rect 5016 17434 5040 17436
rect 5096 17434 5120 17436
rect 5176 17434 5182 17436
rect 4936 17382 4938 17434
rect 5118 17382 5120 17434
rect 4874 17380 4880 17382
rect 4936 17380 4960 17382
rect 5016 17380 5040 17382
rect 5096 17380 5120 17382
rect 5176 17380 5182 17382
rect 4874 17371 5182 17380
rect 4874 16348 5182 16357
rect 4874 16346 4880 16348
rect 4936 16346 4960 16348
rect 5016 16346 5040 16348
rect 5096 16346 5120 16348
rect 5176 16346 5182 16348
rect 4936 16294 4938 16346
rect 5118 16294 5120 16346
rect 4874 16292 4880 16294
rect 4936 16292 4960 16294
rect 5016 16292 5040 16294
rect 5096 16292 5120 16294
rect 5176 16292 5182 16294
rect 4874 16283 5182 16292
rect 4712 15632 4764 15638
rect 4712 15574 4764 15580
rect 4620 15564 4672 15570
rect 4620 15506 4672 15512
rect 3332 15428 3384 15434
rect 3332 15370 3384 15376
rect 3976 15428 4028 15434
rect 3976 15370 4028 15376
rect 3608 15360 3660 15366
rect 3608 15302 3660 15308
rect 3620 15026 3648 15302
rect 3988 15094 4016 15370
rect 4436 15360 4488 15366
rect 4436 15302 4488 15308
rect 3976 15088 4028 15094
rect 3976 15030 4028 15036
rect 3608 15020 3660 15026
rect 3608 14962 3660 14968
rect 3148 14952 3200 14958
rect 3148 14894 3200 14900
rect 3160 14482 3188 14894
rect 4448 14890 4476 15302
rect 4436 14884 4488 14890
rect 4436 14826 4488 14832
rect 4724 14822 4752 15574
rect 4874 15260 5182 15269
rect 4874 15258 4880 15260
rect 4936 15258 4960 15260
rect 5016 15258 5040 15260
rect 5096 15258 5120 15260
rect 5176 15258 5182 15260
rect 4936 15206 4938 15258
rect 5118 15206 5120 15258
rect 4874 15204 4880 15206
rect 4936 15204 4960 15206
rect 5016 15204 5040 15206
rect 5096 15204 5120 15206
rect 5176 15204 5182 15206
rect 4874 15195 5182 15204
rect 4712 14816 4764 14822
rect 4712 14758 4764 14764
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 3240 14612 3292 14618
rect 3240 14554 3292 14560
rect 3148 14476 3200 14482
rect 3148 14418 3200 14424
rect 3160 13462 3188 14418
rect 3148 13456 3200 13462
rect 3148 13398 3200 13404
rect 3252 13394 3280 14554
rect 3332 14408 3384 14414
rect 3332 14350 3384 14356
rect 3344 14006 3372 14350
rect 4436 14272 4488 14278
rect 4436 14214 4488 14220
rect 4528 14272 4580 14278
rect 4528 14214 4580 14220
rect 4712 14272 4764 14278
rect 4712 14214 4764 14220
rect 3332 14000 3384 14006
rect 3332 13942 3384 13948
rect 3240 13388 3292 13394
rect 3240 13330 3292 13336
rect 3252 12986 3280 13330
rect 3240 12980 3292 12986
rect 3240 12922 3292 12928
rect 3344 12434 3372 13942
rect 4448 13938 4476 14214
rect 4540 14074 4568 14214
rect 4528 14068 4580 14074
rect 4528 14010 4580 14016
rect 4436 13932 4488 13938
rect 4436 13874 4488 13880
rect 4724 13870 4752 14214
rect 4874 14172 5182 14181
rect 4874 14170 4880 14172
rect 4936 14170 4960 14172
rect 5016 14170 5040 14172
rect 5096 14170 5120 14172
rect 5176 14170 5182 14172
rect 4936 14118 4938 14170
rect 5118 14118 5120 14170
rect 4874 14116 4880 14118
rect 4936 14116 4960 14118
rect 5016 14116 5040 14118
rect 5096 14116 5120 14118
rect 5176 14116 5182 14118
rect 4874 14107 5182 14116
rect 4712 13864 4764 13870
rect 4712 13806 4764 13812
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4620 13388 4672 13394
rect 4620 13330 4672 13336
rect 4632 12918 4660 13330
rect 4724 13326 4752 13806
rect 4896 13728 4948 13734
rect 4896 13670 4948 13676
rect 4908 13394 4936 13670
rect 4896 13388 4948 13394
rect 4896 13330 4948 13336
rect 4712 13320 4764 13326
rect 4712 13262 4764 13268
rect 4620 12912 4672 12918
rect 4620 12854 4672 12860
rect 4068 12640 4120 12646
rect 4068 12582 4120 12588
rect 3252 12406 3372 12434
rect 4080 12434 4108 12582
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4080 12406 4200 12434
rect 3148 12096 3200 12102
rect 3148 12038 3200 12044
rect 3160 11694 3188 12038
rect 3148 11688 3200 11694
rect 3148 11630 3200 11636
rect 3160 10674 3188 11630
rect 3252 11150 3280 12406
rect 4172 12238 4200 12406
rect 4632 12306 4660 12854
rect 4724 12782 4752 13262
rect 4874 13084 5182 13093
rect 4874 13082 4880 13084
rect 4936 13082 4960 13084
rect 5016 13082 5040 13084
rect 5096 13082 5120 13084
rect 5176 13082 5182 13084
rect 4936 13030 4938 13082
rect 5118 13030 5120 13082
rect 4874 13028 4880 13030
rect 4936 13028 4960 13030
rect 5016 13028 5040 13030
rect 5096 13028 5120 13030
rect 5176 13028 5182 13030
rect 4874 13019 5182 13028
rect 4712 12776 4764 12782
rect 4712 12718 4764 12724
rect 4804 12640 4856 12646
rect 4804 12582 4856 12588
rect 4620 12300 4672 12306
rect 4620 12242 4672 12248
rect 3424 12232 3476 12238
rect 3424 12174 3476 12180
rect 4160 12232 4212 12238
rect 4160 12174 4212 12180
rect 3332 12096 3384 12102
rect 3332 12038 3384 12044
rect 3344 11762 3372 12038
rect 3332 11756 3384 11762
rect 3332 11698 3384 11704
rect 3436 11354 3464 12174
rect 4632 11694 4660 12242
rect 4816 11762 4844 12582
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 4804 11756 4856 11762
rect 4804 11698 4856 11704
rect 4068 11688 4120 11694
rect 4068 11630 4120 11636
rect 4620 11688 4672 11694
rect 4620 11630 4672 11636
rect 3424 11348 3476 11354
rect 3424 11290 3476 11296
rect 3240 11144 3292 11150
rect 3240 11086 3292 11092
rect 4080 11014 4108 11630
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4632 11218 4660 11630
rect 4712 11552 4764 11558
rect 4712 11494 4764 11500
rect 4620 11212 4672 11218
rect 4620 11154 4672 11160
rect 4160 11144 4212 11150
rect 4160 11086 4212 11092
rect 3240 11008 3292 11014
rect 3240 10950 3292 10956
rect 4068 11008 4120 11014
rect 4068 10950 4120 10956
rect 3148 10668 3200 10674
rect 3148 10610 3200 10616
rect 3148 10464 3200 10470
rect 3252 10452 3280 10950
rect 3424 10600 3476 10606
rect 3424 10542 3476 10548
rect 3976 10600 4028 10606
rect 3976 10542 4028 10548
rect 3200 10424 3280 10452
rect 3332 10464 3384 10470
rect 3148 10406 3200 10412
rect 3332 10406 3384 10412
rect 2964 10192 3016 10198
rect 2964 10134 3016 10140
rect 3160 10062 3188 10406
rect 3344 10062 3372 10406
rect 3436 10266 3464 10542
rect 3516 10532 3568 10538
rect 3516 10474 3568 10480
rect 3424 10260 3476 10266
rect 3424 10202 3476 10208
rect 2872 10056 2924 10062
rect 2872 9998 2924 10004
rect 3148 10056 3200 10062
rect 3148 9998 3200 10004
rect 3332 10056 3384 10062
rect 3332 9998 3384 10004
rect 2780 9648 2832 9654
rect 2780 9590 2832 9596
rect 2792 8974 2820 9590
rect 2780 8968 2832 8974
rect 2780 8910 2832 8916
rect 2504 8832 2556 8838
rect 2504 8774 2556 8780
rect 2516 8498 2544 8774
rect 2884 8498 2912 9998
rect 3160 9674 3188 9998
rect 3240 9920 3292 9926
rect 3240 9862 3292 9868
rect 3068 9646 3188 9674
rect 3068 9042 3096 9646
rect 3252 9382 3280 9862
rect 3330 9616 3386 9625
rect 3330 9551 3332 9560
rect 3384 9551 3386 9560
rect 3332 9522 3384 9528
rect 3240 9376 3292 9382
rect 3240 9318 3292 9324
rect 3332 9376 3384 9382
rect 3332 9318 3384 9324
rect 3056 9036 3108 9042
rect 3056 8978 3108 8984
rect 3252 8634 3280 9318
rect 3240 8628 3292 8634
rect 3240 8570 3292 8576
rect 2964 8560 3016 8566
rect 2964 8502 3016 8508
rect 3238 8528 3294 8537
rect 2504 8492 2556 8498
rect 2504 8434 2556 8440
rect 2872 8492 2924 8498
rect 2872 8434 2924 8440
rect 2228 8356 2280 8362
rect 2228 8298 2280 8304
rect 2136 6860 2188 6866
rect 2136 6802 2188 6808
rect 2240 6798 2268 8298
rect 2884 7993 2912 8434
rect 2976 8022 3004 8502
rect 3056 8492 3108 8498
rect 3056 8434 3108 8440
rect 3148 8492 3200 8498
rect 3238 8463 3240 8472
rect 3148 8434 3200 8440
rect 3292 8463 3294 8472
rect 3240 8434 3292 8440
rect 3068 8090 3096 8434
rect 3056 8084 3108 8090
rect 3056 8026 3108 8032
rect 2964 8016 3016 8022
rect 2870 7984 2926 7993
rect 2964 7958 3016 7964
rect 3160 7954 3188 8434
rect 3240 8356 3292 8362
rect 3240 8298 3292 8304
rect 3252 7954 3280 8298
rect 3344 8090 3372 9318
rect 3436 8838 3464 10202
rect 3528 10198 3556 10474
rect 3988 10198 4016 10542
rect 4172 10470 4200 11086
rect 4528 11076 4580 11082
rect 4528 11018 4580 11024
rect 4252 11008 4304 11014
rect 4252 10950 4304 10956
rect 4540 10962 4568 11018
rect 4724 10962 4752 11494
rect 4264 10606 4292 10950
rect 4540 10934 4752 10962
rect 4252 10600 4304 10606
rect 4252 10542 4304 10548
rect 4160 10464 4212 10470
rect 4160 10406 4212 10412
rect 4620 10464 4672 10470
rect 4620 10406 4672 10412
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4528 10260 4580 10266
rect 4528 10202 4580 10208
rect 3516 10192 3568 10198
rect 3516 10134 3568 10140
rect 3976 10192 4028 10198
rect 3976 10134 4028 10140
rect 4158 10160 4214 10169
rect 3988 9518 4016 10134
rect 4158 10095 4214 10104
rect 4344 10124 4396 10130
rect 4172 10062 4200 10095
rect 4344 10066 4396 10072
rect 4160 10056 4212 10062
rect 4160 9998 4212 10004
rect 4160 9920 4212 9926
rect 4160 9862 4212 9868
rect 4172 9586 4200 9862
rect 4356 9722 4384 10066
rect 4344 9716 4396 9722
rect 4344 9658 4396 9664
rect 4160 9580 4212 9586
rect 4160 9522 4212 9528
rect 3976 9512 4028 9518
rect 4172 9466 4200 9522
rect 3976 9454 4028 9460
rect 3608 8968 3660 8974
rect 3608 8910 3660 8916
rect 3988 8922 4016 9454
rect 4080 9438 4200 9466
rect 4080 9042 4108 9438
rect 4540 9382 4568 10202
rect 4528 9376 4580 9382
rect 4528 9318 4580 9324
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4436 9172 4488 9178
rect 4436 9114 4488 9120
rect 4068 9036 4120 9042
rect 4068 8978 4120 8984
rect 4344 9036 4396 9042
rect 4344 8978 4396 8984
rect 3516 8900 3568 8906
rect 3516 8842 3568 8848
rect 3424 8832 3476 8838
rect 3424 8774 3476 8780
rect 3332 8084 3384 8090
rect 3332 8026 3384 8032
rect 3422 7984 3478 7993
rect 2870 7919 2926 7928
rect 3148 7948 3200 7954
rect 3148 7890 3200 7896
rect 3240 7948 3292 7954
rect 3528 7970 3556 8842
rect 3620 8673 3648 8910
rect 3988 8894 4200 8922
rect 3792 8832 3844 8838
rect 3792 8774 3844 8780
rect 4068 8832 4120 8838
rect 4068 8774 4120 8780
rect 3606 8664 3662 8673
rect 3662 8622 3740 8650
rect 3606 8599 3662 8608
rect 3606 8528 3662 8537
rect 3606 8463 3662 8472
rect 3620 8090 3648 8463
rect 3608 8084 3660 8090
rect 3608 8026 3660 8032
rect 3528 7942 3648 7970
rect 3712 7954 3740 8622
rect 3422 7919 3478 7928
rect 3240 7890 3292 7896
rect 2872 7744 2924 7750
rect 2872 7686 2924 7692
rect 2884 7546 2912 7686
rect 3160 7562 3188 7890
rect 3436 7886 3464 7919
rect 3424 7880 3476 7886
rect 3424 7822 3476 7828
rect 2872 7540 2924 7546
rect 3160 7534 3280 7562
rect 2872 7482 2924 7488
rect 3148 7404 3200 7410
rect 3148 7346 3200 7352
rect 2504 6860 2556 6866
rect 2504 6802 2556 6808
rect 2228 6792 2280 6798
rect 2228 6734 2280 6740
rect 1676 6656 1728 6662
rect 1676 6598 1728 6604
rect 1688 6390 1716 6598
rect 2516 6458 2544 6802
rect 3160 6730 3188 7346
rect 3252 7206 3280 7534
rect 3620 7478 3648 7942
rect 3700 7948 3752 7954
rect 3700 7890 3752 7896
rect 3608 7472 3660 7478
rect 3608 7414 3660 7420
rect 3516 7404 3568 7410
rect 3516 7346 3568 7352
rect 3240 7200 3292 7206
rect 3240 7142 3292 7148
rect 3528 6798 3556 7346
rect 3620 7002 3648 7414
rect 3608 6996 3660 7002
rect 3608 6938 3660 6944
rect 3516 6792 3568 6798
rect 3568 6740 3648 6746
rect 3516 6734 3648 6740
rect 3148 6724 3200 6730
rect 3528 6718 3648 6734
rect 3148 6666 3200 6672
rect 3160 6458 3188 6666
rect 2504 6452 2556 6458
rect 2504 6394 2556 6400
rect 3148 6452 3200 6458
rect 3148 6394 3200 6400
rect 1676 6384 1728 6390
rect 1676 6326 1728 6332
rect 3620 6254 3648 6718
rect 3804 6458 3832 8774
rect 4080 8634 4108 8774
rect 4172 8634 4200 8894
rect 4252 8900 4304 8906
rect 4252 8842 4304 8848
rect 4068 8628 4120 8634
rect 4068 8570 4120 8576
rect 4160 8628 4212 8634
rect 4160 8570 4212 8576
rect 4158 8528 4214 8537
rect 3976 8492 4028 8498
rect 3896 8452 3976 8480
rect 3896 7993 3924 8452
rect 4158 8463 4160 8472
rect 3976 8434 4028 8440
rect 4212 8463 4214 8472
rect 4160 8434 4212 8440
rect 4264 8378 4292 8842
rect 4356 8498 4384 8978
rect 4448 8906 4476 9114
rect 4436 8900 4488 8906
rect 4436 8842 4488 8848
rect 4448 8537 4476 8842
rect 4434 8528 4490 8537
rect 4344 8492 4396 8498
rect 4434 8463 4490 8472
rect 4344 8434 4396 8440
rect 4080 8350 4292 8378
rect 3976 8288 4028 8294
rect 3976 8230 4028 8236
rect 3882 7984 3938 7993
rect 3882 7919 3938 7928
rect 3988 7886 4016 8230
rect 3976 7880 4028 7886
rect 3976 7822 4028 7828
rect 3884 7812 3936 7818
rect 3884 7754 3936 7760
rect 3896 7410 3924 7754
rect 4080 7546 4108 8350
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4344 7880 4396 7886
rect 4344 7822 4396 7828
rect 4252 7744 4304 7750
rect 4252 7686 4304 7692
rect 4068 7540 4120 7546
rect 4068 7482 4120 7488
rect 4160 7540 4212 7546
rect 4160 7482 4212 7488
rect 3884 7404 3936 7410
rect 3884 7346 3936 7352
rect 3896 6934 3924 7346
rect 4172 7290 4200 7482
rect 4264 7410 4292 7686
rect 4356 7546 4384 7822
rect 4344 7540 4396 7546
rect 4344 7482 4396 7488
rect 4252 7404 4304 7410
rect 4252 7346 4304 7352
rect 4264 7313 4292 7346
rect 4080 7262 4200 7290
rect 4250 7304 4306 7313
rect 4080 6984 4108 7262
rect 4250 7239 4306 7248
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4080 6956 4200 6984
rect 3884 6928 3936 6934
rect 3884 6870 3936 6876
rect 4172 6798 4200 6956
rect 4160 6792 4212 6798
rect 4160 6734 4212 6740
rect 4252 6724 4304 6730
rect 4252 6666 4304 6672
rect 3884 6656 3936 6662
rect 3884 6598 3936 6604
rect 3792 6452 3844 6458
rect 3792 6394 3844 6400
rect 1400 6248 1452 6254
rect 1400 6190 1452 6196
rect 2872 6248 2924 6254
rect 2872 6190 2924 6196
rect 3608 6248 3660 6254
rect 3608 6190 3660 6196
rect 1412 5778 1440 6190
rect 1400 5772 1452 5778
rect 1400 5714 1452 5720
rect 2884 5710 2912 6190
rect 3240 6112 3292 6118
rect 3240 6054 3292 6060
rect 3252 5914 3280 6054
rect 3240 5908 3292 5914
rect 3240 5850 3292 5856
rect 2872 5704 2924 5710
rect 2872 5646 2924 5652
rect 2884 5166 2912 5646
rect 3620 5574 3648 6190
rect 3700 5772 3752 5778
rect 3700 5714 3752 5720
rect 3608 5568 3660 5574
rect 3608 5510 3660 5516
rect 3712 5234 3740 5714
rect 3896 5302 3924 6598
rect 4264 6458 4292 6666
rect 4252 6452 4304 6458
rect 4252 6394 4304 6400
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4632 5778 4660 10406
rect 4724 10033 4752 10934
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 5276 10266 5304 18022
rect 5724 16584 5776 16590
rect 5724 16526 5776 16532
rect 5736 16250 5764 16526
rect 6104 16522 6132 18226
rect 8680 17202 8708 18226
rect 8668 17196 8720 17202
rect 8668 17138 8720 17144
rect 6920 16652 6972 16658
rect 6920 16594 6972 16600
rect 8208 16652 8260 16658
rect 8208 16594 8260 16600
rect 6092 16516 6144 16522
rect 6092 16458 6144 16464
rect 5724 16244 5776 16250
rect 5724 16186 5776 16192
rect 5908 16040 5960 16046
rect 5908 15982 5960 15988
rect 6000 16040 6052 16046
rect 6000 15982 6052 15988
rect 5356 15904 5408 15910
rect 5356 15846 5408 15852
rect 5368 15570 5396 15846
rect 5356 15564 5408 15570
rect 5356 15506 5408 15512
rect 5356 14816 5408 14822
rect 5356 14758 5408 14764
rect 5368 13802 5396 14758
rect 5920 14618 5948 15982
rect 6012 15094 6040 15982
rect 6104 15706 6132 16458
rect 6932 16250 6960 16594
rect 7840 16448 7892 16454
rect 7840 16390 7892 16396
rect 6920 16244 6972 16250
rect 6920 16186 6972 16192
rect 7852 16114 7880 16390
rect 6828 16108 6880 16114
rect 6828 16050 6880 16056
rect 7840 16108 7892 16114
rect 7840 16050 7892 16056
rect 6092 15700 6144 15706
rect 6092 15642 6144 15648
rect 6104 15434 6132 15642
rect 6840 15570 6868 16050
rect 8220 15706 8248 16594
rect 8680 16250 8708 17138
rect 8852 16788 8904 16794
rect 8852 16730 8904 16736
rect 8668 16244 8720 16250
rect 8668 16186 8720 16192
rect 7748 15700 7800 15706
rect 7748 15642 7800 15648
rect 8208 15700 8260 15706
rect 8208 15642 8260 15648
rect 6828 15564 6880 15570
rect 6828 15506 6880 15512
rect 6092 15428 6144 15434
rect 6092 15370 6144 15376
rect 6000 15088 6052 15094
rect 6000 15030 6052 15036
rect 5908 14612 5960 14618
rect 5908 14554 5960 14560
rect 6012 14482 6040 15030
rect 6000 14476 6052 14482
rect 6000 14418 6052 14424
rect 5632 14408 5684 14414
rect 5632 14350 5684 14356
rect 5540 14272 5592 14278
rect 5540 14214 5592 14220
rect 5356 13796 5408 13802
rect 5356 13738 5408 13744
rect 5368 12782 5396 13738
rect 5552 13394 5580 14214
rect 5644 13938 5672 14350
rect 6104 14346 6132 15370
rect 6828 15088 6880 15094
rect 6828 15030 6880 15036
rect 6644 15020 6696 15026
rect 6644 14962 6696 14968
rect 6552 14952 6604 14958
rect 6552 14894 6604 14900
rect 6460 14816 6512 14822
rect 6460 14758 6512 14764
rect 6472 14482 6500 14758
rect 6460 14476 6512 14482
rect 6460 14418 6512 14424
rect 6564 14414 6592 14894
rect 6656 14618 6684 14962
rect 6840 14634 6868 15030
rect 7656 14816 7708 14822
rect 7656 14758 7708 14764
rect 6644 14612 6696 14618
rect 6840 14606 6960 14634
rect 6644 14554 6696 14560
rect 6552 14408 6604 14414
rect 6552 14350 6604 14356
rect 6092 14340 6144 14346
rect 6092 14282 6144 14288
rect 5632 13932 5684 13938
rect 5632 13874 5684 13880
rect 5540 13388 5592 13394
rect 5540 13330 5592 13336
rect 6564 13190 6592 14350
rect 6656 14006 6684 14554
rect 6828 14544 6880 14550
rect 6748 14492 6828 14498
rect 6748 14486 6880 14492
rect 6748 14470 6868 14486
rect 6932 14482 6960 14606
rect 6920 14476 6972 14482
rect 6644 14000 6696 14006
rect 6644 13942 6696 13948
rect 6644 13864 6696 13870
rect 6748 13818 6776 14470
rect 6920 14418 6972 14424
rect 6828 14408 6880 14414
rect 6828 14350 6880 14356
rect 6696 13812 6776 13818
rect 6644 13806 6776 13812
rect 6656 13790 6776 13806
rect 6656 13326 6684 13790
rect 6736 13728 6788 13734
rect 6736 13670 6788 13676
rect 6644 13320 6696 13326
rect 6644 13262 6696 13268
rect 6552 13184 6604 13190
rect 6552 13126 6604 13132
rect 6276 12844 6328 12850
rect 6276 12786 6328 12792
rect 5356 12776 5408 12782
rect 5356 12718 5408 12724
rect 5724 12164 5776 12170
rect 5724 12106 5776 12112
rect 5736 11830 5764 12106
rect 6288 12102 6316 12786
rect 6276 12096 6328 12102
rect 6276 12038 6328 12044
rect 5724 11824 5776 11830
rect 5724 11766 5776 11772
rect 5736 11082 5764 11766
rect 6288 11150 6316 12038
rect 6564 11898 6592 13126
rect 6644 12980 6696 12986
rect 6644 12922 6696 12928
rect 6656 12442 6684 12922
rect 6748 12850 6776 13670
rect 6840 13394 6868 14350
rect 7380 14272 7432 14278
rect 7380 14214 7432 14220
rect 7392 14074 7420 14214
rect 7380 14068 7432 14074
rect 7380 14010 7432 14016
rect 7472 13932 7524 13938
rect 7472 13874 7524 13880
rect 6920 13796 6972 13802
rect 6920 13738 6972 13744
rect 6828 13388 6880 13394
rect 6828 13330 6880 13336
rect 6736 12844 6788 12850
rect 6736 12786 6788 12792
rect 6644 12436 6696 12442
rect 6644 12378 6696 12384
rect 6552 11892 6604 11898
rect 6552 11834 6604 11840
rect 6656 11830 6684 12378
rect 6840 12238 6868 13330
rect 6828 12232 6880 12238
rect 6828 12174 6880 12180
rect 6644 11824 6696 11830
rect 6644 11766 6696 11772
rect 6736 11756 6788 11762
rect 6736 11698 6788 11704
rect 6368 11552 6420 11558
rect 6368 11494 6420 11500
rect 6380 11218 6408 11494
rect 6748 11354 6776 11698
rect 6736 11348 6788 11354
rect 6736 11290 6788 11296
rect 6840 11218 6868 12174
rect 6932 11694 6960 13738
rect 7484 13734 7512 13874
rect 7196 13728 7248 13734
rect 7196 13670 7248 13676
rect 7472 13728 7524 13734
rect 7472 13670 7524 13676
rect 7208 13394 7236 13670
rect 7196 13388 7248 13394
rect 7196 13330 7248 13336
rect 7484 12986 7512 13670
rect 7472 12980 7524 12986
rect 7472 12922 7524 12928
rect 7104 12912 7156 12918
rect 7104 12854 7156 12860
rect 7116 12170 7144 12854
rect 7668 12434 7696 14758
rect 7760 13870 7788 15642
rect 7840 15360 7892 15366
rect 7840 15302 7892 15308
rect 7852 14958 7880 15302
rect 8680 14958 8708 16186
rect 8864 16182 8892 16730
rect 8852 16176 8904 16182
rect 8852 16118 8904 16124
rect 8864 15502 8892 16118
rect 8852 15496 8904 15502
rect 8852 15438 8904 15444
rect 8864 15094 8892 15438
rect 8852 15088 8904 15094
rect 8852 15030 8904 15036
rect 7840 14952 7892 14958
rect 7840 14894 7892 14900
rect 8668 14952 8720 14958
rect 8668 14894 8720 14900
rect 8956 14890 8984 19314
rect 9324 18902 9352 19450
rect 9312 18896 9364 18902
rect 9312 18838 9364 18844
rect 9220 18828 9272 18834
rect 9220 18770 9272 18776
rect 9232 18358 9260 18770
rect 9692 18766 9720 19654
rect 9784 19378 9812 19790
rect 9772 19372 9824 19378
rect 9772 19314 9824 19320
rect 9876 18970 9904 20946
rect 10048 20868 10100 20874
rect 10048 20810 10100 20816
rect 10060 20602 10088 20810
rect 10048 20596 10100 20602
rect 10048 20538 10100 20544
rect 9864 18964 9916 18970
rect 9864 18906 9916 18912
rect 9680 18760 9732 18766
rect 9680 18702 9732 18708
rect 9220 18352 9272 18358
rect 9220 18294 9272 18300
rect 9588 17672 9640 17678
rect 9588 17614 9640 17620
rect 9600 17202 9628 17614
rect 9876 17270 9904 18906
rect 10048 18284 10100 18290
rect 10152 18272 10180 22066
rect 10244 21010 10272 24550
rect 10520 24410 10548 25094
rect 10508 24404 10560 24410
rect 10508 24346 10560 24352
rect 10520 24206 10548 24346
rect 10416 24200 10468 24206
rect 10416 24142 10468 24148
rect 10508 24200 10560 24206
rect 10508 24142 10560 24148
rect 10324 23180 10376 23186
rect 10324 23122 10376 23128
rect 10336 22030 10364 23122
rect 10324 22024 10376 22030
rect 10324 21966 10376 21972
rect 10428 21146 10456 24142
rect 10508 22568 10560 22574
rect 10508 22510 10560 22516
rect 10520 22234 10548 22510
rect 10508 22228 10560 22234
rect 10508 22170 10560 22176
rect 10612 21962 10640 25774
rect 12808 25764 12860 25770
rect 12808 25706 12860 25712
rect 13912 25764 13964 25770
rect 13912 25706 13964 25712
rect 14648 25764 14700 25770
rect 14648 25706 14700 25712
rect 11060 25696 11112 25702
rect 11060 25638 11112 25644
rect 11888 25696 11940 25702
rect 11888 25638 11940 25644
rect 11072 25294 11100 25638
rect 11060 25288 11112 25294
rect 11060 25230 11112 25236
rect 11336 25220 11388 25226
rect 11336 25162 11388 25168
rect 10968 25152 11020 25158
rect 10968 25094 11020 25100
rect 11244 25152 11296 25158
rect 11244 25094 11296 25100
rect 10784 24812 10836 24818
rect 10784 24754 10836 24760
rect 10796 24342 10824 24754
rect 10784 24336 10836 24342
rect 10784 24278 10836 24284
rect 10796 24206 10824 24278
rect 10784 24200 10836 24206
rect 10784 24142 10836 24148
rect 10692 23520 10744 23526
rect 10692 23462 10744 23468
rect 10704 23118 10732 23462
rect 10692 23112 10744 23118
rect 10692 23054 10744 23060
rect 10692 22976 10744 22982
rect 10692 22918 10744 22924
rect 10704 22642 10732 22918
rect 10692 22636 10744 22642
rect 10744 22596 10916 22624
rect 10692 22578 10744 22584
rect 10600 21956 10652 21962
rect 10600 21898 10652 21904
rect 10612 21350 10640 21898
rect 10784 21548 10836 21554
rect 10784 21490 10836 21496
rect 10600 21344 10652 21350
rect 10600 21286 10652 21292
rect 10416 21140 10468 21146
rect 10416 21082 10468 21088
rect 10232 21004 10284 21010
rect 10232 20946 10284 20952
rect 10508 20936 10560 20942
rect 10508 20878 10560 20884
rect 10520 19310 10548 20878
rect 10612 20534 10640 21286
rect 10796 20874 10824 21490
rect 10784 20868 10836 20874
rect 10784 20810 10836 20816
rect 10600 20528 10652 20534
rect 10600 20470 10652 20476
rect 10600 20392 10652 20398
rect 10600 20334 10652 20340
rect 10508 19304 10560 19310
rect 10508 19246 10560 19252
rect 10612 18426 10640 20334
rect 10888 19514 10916 22596
rect 10980 22094 11008 25094
rect 11152 24404 11204 24410
rect 11152 24346 11204 24352
rect 11164 24206 11192 24346
rect 11152 24200 11204 24206
rect 11152 24142 11204 24148
rect 11060 24064 11112 24070
rect 11060 24006 11112 24012
rect 11072 23730 11100 24006
rect 11256 23866 11284 25094
rect 11244 23860 11296 23866
rect 11244 23802 11296 23808
rect 11060 23724 11112 23730
rect 11060 23666 11112 23672
rect 11060 23588 11112 23594
rect 11060 23530 11112 23536
rect 11152 23588 11204 23594
rect 11152 23530 11204 23536
rect 11072 23322 11100 23530
rect 11060 23316 11112 23322
rect 11060 23258 11112 23264
rect 11164 23202 11192 23530
rect 11244 23520 11296 23526
rect 11244 23462 11296 23468
rect 11256 23322 11284 23462
rect 11244 23316 11296 23322
rect 11244 23258 11296 23264
rect 11072 23186 11192 23202
rect 11060 23180 11192 23186
rect 11112 23174 11192 23180
rect 11060 23122 11112 23128
rect 10980 22066 11100 22094
rect 11072 22001 11100 22066
rect 11058 21992 11114 22001
rect 11058 21927 11114 21936
rect 10876 19508 10928 19514
rect 10876 19450 10928 19456
rect 10968 18692 11020 18698
rect 10968 18634 11020 18640
rect 10600 18420 10652 18426
rect 10600 18362 10652 18368
rect 10100 18244 10180 18272
rect 10048 18226 10100 18232
rect 9864 17264 9916 17270
rect 9864 17206 9916 17212
rect 9588 17196 9640 17202
rect 9588 17138 9640 17144
rect 9312 16516 9364 16522
rect 9312 16458 9364 16464
rect 9036 16448 9088 16454
rect 9036 16390 9088 16396
rect 9048 16182 9076 16390
rect 9036 16176 9088 16182
rect 9036 16118 9088 16124
rect 9324 15502 9352 16458
rect 9600 15570 9628 17138
rect 10060 16794 10088 18226
rect 10612 17746 10640 18362
rect 10980 18358 11008 18634
rect 10968 18352 11020 18358
rect 10968 18294 11020 18300
rect 11152 18352 11204 18358
rect 11152 18294 11204 18300
rect 10600 17740 10652 17746
rect 10600 17682 10652 17688
rect 11164 17338 11192 18294
rect 11348 17610 11376 25162
rect 11702 24168 11758 24177
rect 11702 24103 11758 24112
rect 11428 23112 11480 23118
rect 11428 23054 11480 23060
rect 11440 19446 11468 23054
rect 11520 22024 11572 22030
rect 11520 21966 11572 21972
rect 11532 21894 11560 21966
rect 11520 21888 11572 21894
rect 11520 21830 11572 21836
rect 11716 21554 11744 24103
rect 11796 24064 11848 24070
rect 11796 24006 11848 24012
rect 11808 23730 11836 24006
rect 11796 23724 11848 23730
rect 11796 23666 11848 23672
rect 11900 22817 11928 25638
rect 12072 25356 12124 25362
rect 12072 25298 12124 25304
rect 11886 22808 11942 22817
rect 11886 22743 11942 22752
rect 11900 22710 11928 22743
rect 11888 22704 11940 22710
rect 11888 22646 11940 22652
rect 11980 22432 12032 22438
rect 11980 22374 12032 22380
rect 11888 22024 11940 22030
rect 11888 21966 11940 21972
rect 11900 21622 11928 21966
rect 11888 21616 11940 21622
rect 11888 21558 11940 21564
rect 11520 21548 11572 21554
rect 11520 21490 11572 21496
rect 11704 21548 11756 21554
rect 11704 21490 11756 21496
rect 11532 19990 11560 21490
rect 11992 21418 12020 22374
rect 12084 22166 12112 25298
rect 12716 25220 12768 25226
rect 12716 25162 12768 25168
rect 12532 24812 12584 24818
rect 12532 24754 12584 24760
rect 12164 23860 12216 23866
rect 12164 23802 12216 23808
rect 12176 23594 12204 23802
rect 12440 23724 12492 23730
rect 12440 23666 12492 23672
rect 12164 23588 12216 23594
rect 12164 23530 12216 23536
rect 12348 23588 12400 23594
rect 12348 23530 12400 23536
rect 12176 23322 12204 23530
rect 12164 23316 12216 23322
rect 12164 23258 12216 23264
rect 12164 22636 12216 22642
rect 12164 22578 12216 22584
rect 12256 22636 12308 22642
rect 12256 22578 12308 22584
rect 12072 22160 12124 22166
rect 12072 22102 12124 22108
rect 12176 22098 12204 22578
rect 12164 22092 12216 22098
rect 12164 22034 12216 22040
rect 12072 22024 12124 22030
rect 12072 21966 12124 21972
rect 12162 21992 12218 22001
rect 12084 21690 12112 21966
rect 12162 21927 12218 21936
rect 12072 21684 12124 21690
rect 12072 21626 12124 21632
rect 12176 21593 12204 21927
rect 12268 21690 12296 22578
rect 12256 21684 12308 21690
rect 12256 21626 12308 21632
rect 12162 21584 12218 21593
rect 12162 21519 12164 21528
rect 12216 21519 12218 21528
rect 12164 21490 12216 21496
rect 11980 21412 12032 21418
rect 11980 21354 12032 21360
rect 11520 19984 11572 19990
rect 11520 19926 11572 19932
rect 12072 19984 12124 19990
rect 12360 19972 12388 23530
rect 12452 23118 12480 23666
rect 12544 23526 12572 24754
rect 12728 24750 12756 25162
rect 12716 24744 12768 24750
rect 12716 24686 12768 24692
rect 12728 24410 12756 24686
rect 12716 24404 12768 24410
rect 12716 24346 12768 24352
rect 12820 24274 12848 25706
rect 13820 25696 13872 25702
rect 13820 25638 13872 25644
rect 13360 25356 13412 25362
rect 13360 25298 13412 25304
rect 12992 25288 13044 25294
rect 12992 25230 13044 25236
rect 13004 24750 13032 25230
rect 13372 24750 13400 25298
rect 13544 25152 13596 25158
rect 13544 25094 13596 25100
rect 12992 24744 13044 24750
rect 12992 24686 13044 24692
rect 13360 24744 13412 24750
rect 13360 24686 13412 24692
rect 12900 24608 12952 24614
rect 12900 24550 12952 24556
rect 12912 24274 12940 24550
rect 13372 24410 13400 24686
rect 13360 24404 13412 24410
rect 13360 24346 13412 24352
rect 12808 24268 12860 24274
rect 12808 24210 12860 24216
rect 12900 24268 12952 24274
rect 12900 24210 12952 24216
rect 12624 24200 12676 24206
rect 12624 24142 12676 24148
rect 12636 23866 12664 24142
rect 12716 24064 12768 24070
rect 12716 24006 12768 24012
rect 12624 23860 12676 23866
rect 12624 23802 12676 23808
rect 12532 23520 12584 23526
rect 12532 23462 12584 23468
rect 12532 23316 12584 23322
rect 12532 23258 12584 23264
rect 12440 23112 12492 23118
rect 12440 23054 12492 23060
rect 12544 22778 12572 23258
rect 12532 22772 12584 22778
rect 12532 22714 12584 22720
rect 12532 22636 12584 22642
rect 12532 22578 12584 22584
rect 12440 22500 12492 22506
rect 12440 22442 12492 22448
rect 12452 21690 12480 22442
rect 12544 22098 12572 22578
rect 12728 22574 12756 24006
rect 12820 23848 12848 24210
rect 13556 24206 13584 25094
rect 13728 24744 13780 24750
rect 13728 24686 13780 24692
rect 13268 24200 13320 24206
rect 13360 24200 13412 24206
rect 13268 24142 13320 24148
rect 13358 24168 13360 24177
rect 13544 24200 13596 24206
rect 13412 24168 13414 24177
rect 12900 23860 12952 23866
rect 12820 23820 12900 23848
rect 12900 23802 12952 23808
rect 12992 23792 13044 23798
rect 12806 23760 12862 23769
rect 12992 23734 13044 23740
rect 12900 23724 12952 23730
rect 12862 23704 12900 23712
rect 12806 23695 12900 23704
rect 12820 23684 12900 23695
rect 12820 23254 12848 23684
rect 12900 23666 12952 23672
rect 13004 23254 13032 23734
rect 13084 23724 13136 23730
rect 13084 23666 13136 23672
rect 12808 23248 12860 23254
rect 12808 23190 12860 23196
rect 12992 23248 13044 23254
rect 12992 23190 13044 23196
rect 12716 22568 12768 22574
rect 12716 22510 12768 22516
rect 12728 22166 12756 22510
rect 12716 22160 12768 22166
rect 12716 22102 12768 22108
rect 12532 22092 12584 22098
rect 12532 22034 12584 22040
rect 12624 22024 12676 22030
rect 12624 21966 12676 21972
rect 12532 21956 12584 21962
rect 12532 21898 12584 21904
rect 12440 21684 12492 21690
rect 12440 21626 12492 21632
rect 12544 21554 12572 21898
rect 12636 21690 12664 21966
rect 12716 21888 12768 21894
rect 12716 21830 12768 21836
rect 12624 21684 12676 21690
rect 12624 21626 12676 21632
rect 12532 21548 12584 21554
rect 12532 21490 12584 21496
rect 12544 19990 12572 21490
rect 12124 19944 12388 19972
rect 12072 19926 12124 19932
rect 12164 19508 12216 19514
rect 12164 19450 12216 19456
rect 11428 19440 11480 19446
rect 11428 19382 11480 19388
rect 11888 19440 11940 19446
rect 11888 19382 11940 19388
rect 11900 18902 11928 19382
rect 12072 19168 12124 19174
rect 12072 19110 12124 19116
rect 11888 18896 11940 18902
rect 11888 18838 11940 18844
rect 12084 18766 12112 19110
rect 12176 18766 12204 19450
rect 12360 18850 12388 19944
rect 12532 19984 12584 19990
rect 12532 19926 12584 19932
rect 12544 19446 12572 19926
rect 12728 19718 12756 21830
rect 12820 20466 12848 23190
rect 12900 23112 12952 23118
rect 12900 23054 12952 23060
rect 12912 22710 12940 23054
rect 12992 22772 13044 22778
rect 12992 22714 13044 22720
rect 12900 22704 12952 22710
rect 12900 22646 12952 22652
rect 13004 22658 13032 22714
rect 13096 22658 13124 23666
rect 13280 23610 13308 24142
rect 13544 24142 13596 24148
rect 13358 24103 13414 24112
rect 13740 24070 13768 24686
rect 13728 24064 13780 24070
rect 13728 24006 13780 24012
rect 13360 23792 13412 23798
rect 13358 23760 13360 23769
rect 13412 23760 13414 23769
rect 13358 23695 13414 23704
rect 13280 23582 13492 23610
rect 13268 23520 13320 23526
rect 13268 23462 13320 23468
rect 13176 22772 13228 22778
rect 13176 22714 13228 22720
rect 12912 21486 12940 22646
rect 13004 22630 13124 22658
rect 13188 22642 13216 22714
rect 12992 22432 13044 22438
rect 12992 22374 13044 22380
rect 13004 22234 13032 22374
rect 13096 22250 13124 22630
rect 13176 22636 13228 22642
rect 13176 22578 13228 22584
rect 13096 22234 13140 22250
rect 13188 22234 13216 22578
rect 12992 22228 13044 22234
rect 12992 22170 13044 22176
rect 13084 22228 13140 22234
rect 13136 22188 13140 22228
rect 13176 22228 13228 22234
rect 13084 22170 13136 22176
rect 13176 22170 13228 22176
rect 13280 22098 13308 23462
rect 13464 22982 13492 23582
rect 13544 23112 13596 23118
rect 13544 23054 13596 23060
rect 13452 22976 13504 22982
rect 13452 22918 13504 22924
rect 13464 22420 13492 22918
rect 13556 22522 13584 23054
rect 13740 22778 13768 24006
rect 13728 22772 13780 22778
rect 13728 22714 13780 22720
rect 13832 22710 13860 25638
rect 13820 22704 13872 22710
rect 13820 22646 13872 22652
rect 13556 22494 13676 22522
rect 13372 22392 13492 22420
rect 13544 22432 13596 22438
rect 13372 22098 13400 22392
rect 13544 22374 13596 22380
rect 13452 22160 13504 22166
rect 13452 22102 13504 22108
rect 12992 22092 13044 22098
rect 12992 22034 13044 22040
rect 13084 22092 13136 22098
rect 13084 22034 13136 22040
rect 13268 22092 13320 22098
rect 13268 22034 13320 22040
rect 13360 22092 13412 22098
rect 13360 22034 13412 22040
rect 13004 21690 13032 22034
rect 12992 21684 13044 21690
rect 12992 21626 13044 21632
rect 12900 21480 12952 21486
rect 12900 21422 12952 21428
rect 12992 21344 13044 21350
rect 12992 21286 13044 21292
rect 13004 20942 13032 21286
rect 12992 20936 13044 20942
rect 12992 20878 13044 20884
rect 13096 20534 13124 22034
rect 13360 21956 13412 21962
rect 13360 21898 13412 21904
rect 13372 21554 13400 21898
rect 13464 21554 13492 22102
rect 13556 21962 13584 22374
rect 13648 22166 13676 22494
rect 13636 22160 13688 22166
rect 13636 22102 13688 22108
rect 13544 21956 13596 21962
rect 13544 21898 13596 21904
rect 13268 21548 13320 21554
rect 13268 21490 13320 21496
rect 13360 21548 13412 21554
rect 13360 21490 13412 21496
rect 13452 21548 13504 21554
rect 13452 21490 13504 21496
rect 13636 21548 13688 21554
rect 13636 21490 13688 21496
rect 13728 21548 13780 21554
rect 13728 21490 13780 21496
rect 13084 20528 13136 20534
rect 13084 20470 13136 20476
rect 12808 20460 12860 20466
rect 12808 20402 12860 20408
rect 12900 20392 12952 20398
rect 12900 20334 12952 20340
rect 12716 19712 12768 19718
rect 12716 19654 12768 19660
rect 12532 19440 12584 19446
rect 12532 19382 12584 19388
rect 12728 19310 12756 19654
rect 12440 19304 12492 19310
rect 12440 19246 12492 19252
rect 12716 19304 12768 19310
rect 12716 19246 12768 19252
rect 12452 18970 12480 19246
rect 12808 19168 12860 19174
rect 12808 19110 12860 19116
rect 12440 18964 12492 18970
rect 12440 18906 12492 18912
rect 12716 18964 12768 18970
rect 12716 18906 12768 18912
rect 12728 18873 12756 18906
rect 12438 18864 12494 18873
rect 12360 18822 12438 18850
rect 12438 18799 12494 18808
rect 12714 18864 12770 18873
rect 12714 18799 12770 18808
rect 12072 18760 12124 18766
rect 12072 18702 12124 18708
rect 12164 18760 12216 18766
rect 12164 18702 12216 18708
rect 12084 17882 12112 18702
rect 12176 18358 12204 18702
rect 12452 18358 12480 18799
rect 12820 18630 12848 19110
rect 12912 18714 12940 20334
rect 13096 19514 13124 20470
rect 13084 19508 13136 19514
rect 13084 19450 13136 19456
rect 13084 19304 13136 19310
rect 13084 19246 13136 19252
rect 13096 18766 13124 19246
rect 13084 18760 13136 18766
rect 12912 18686 13032 18714
rect 13084 18702 13136 18708
rect 12808 18624 12860 18630
rect 12808 18566 12860 18572
rect 12900 18624 12952 18630
rect 12900 18566 12952 18572
rect 12164 18352 12216 18358
rect 12164 18294 12216 18300
rect 12440 18352 12492 18358
rect 12440 18294 12492 18300
rect 12452 18086 12480 18294
rect 12440 18080 12492 18086
rect 12440 18022 12492 18028
rect 12716 18080 12768 18086
rect 12912 18068 12940 18566
rect 13004 18086 13032 18686
rect 13280 18426 13308 21490
rect 13360 21004 13412 21010
rect 13360 20946 13412 20952
rect 13372 20602 13400 20946
rect 13360 20596 13412 20602
rect 13360 20538 13412 20544
rect 13452 20460 13504 20466
rect 13452 20402 13504 20408
rect 13464 20058 13492 20402
rect 13648 20398 13676 21490
rect 13740 21146 13768 21490
rect 13728 21140 13780 21146
rect 13728 21082 13780 21088
rect 13832 20942 13860 22646
rect 13820 20936 13872 20942
rect 13820 20878 13872 20884
rect 13924 20874 13952 25706
rect 14464 24812 14516 24818
rect 14464 24754 14516 24760
rect 14476 24274 14504 24754
rect 14464 24268 14516 24274
rect 14464 24210 14516 24216
rect 14096 23656 14148 23662
rect 14096 23598 14148 23604
rect 14108 23322 14136 23598
rect 14278 23488 14334 23497
rect 14278 23423 14334 23432
rect 14096 23316 14148 23322
rect 14096 23258 14148 23264
rect 14108 22642 14136 23258
rect 14188 23180 14240 23186
rect 14188 23122 14240 23128
rect 14096 22636 14148 22642
rect 14096 22578 14148 22584
rect 14200 22420 14228 23122
rect 14292 23050 14320 23423
rect 14476 23118 14504 24210
rect 14464 23112 14516 23118
rect 14464 23054 14516 23060
rect 14280 23044 14332 23050
rect 14280 22986 14332 22992
rect 14464 22704 14516 22710
rect 14464 22646 14516 22652
rect 14280 22568 14332 22574
rect 14476 22556 14504 22646
rect 14332 22528 14504 22556
rect 14280 22510 14332 22516
rect 14280 22432 14332 22438
rect 14200 22392 14280 22420
rect 14280 22374 14332 22380
rect 13912 20868 13964 20874
rect 13912 20810 13964 20816
rect 14660 20534 14688 25706
rect 16948 25696 17000 25702
rect 16948 25638 17000 25644
rect 17408 25696 17460 25702
rect 17408 25638 17460 25644
rect 15292 25288 15344 25294
rect 15292 25230 15344 25236
rect 15476 25288 15528 25294
rect 15476 25230 15528 25236
rect 14740 24948 14792 24954
rect 14740 24890 14792 24896
rect 14752 22710 14780 24890
rect 14924 24744 14976 24750
rect 14924 24686 14976 24692
rect 14936 23322 14964 24686
rect 15016 24608 15068 24614
rect 15016 24550 15068 24556
rect 15028 24138 15056 24550
rect 15016 24132 15068 24138
rect 15016 24074 15068 24080
rect 15108 23792 15160 23798
rect 15108 23734 15160 23740
rect 15120 23526 15148 23734
rect 15304 23662 15332 25230
rect 15488 24682 15516 25230
rect 15844 25220 15896 25226
rect 15844 25162 15896 25168
rect 16856 25220 16908 25226
rect 16856 25162 16908 25168
rect 15856 24954 15884 25162
rect 15844 24948 15896 24954
rect 15844 24890 15896 24896
rect 16028 24812 16080 24818
rect 16028 24754 16080 24760
rect 15476 24676 15528 24682
rect 15476 24618 15528 24624
rect 15384 24200 15436 24206
rect 15488 24154 15516 24618
rect 15436 24148 15516 24154
rect 15384 24142 15516 24148
rect 15396 24126 15516 24142
rect 15292 23656 15344 23662
rect 15292 23598 15344 23604
rect 15108 23520 15160 23526
rect 15108 23462 15160 23468
rect 14924 23316 14976 23322
rect 14924 23258 14976 23264
rect 15488 23186 15516 24126
rect 15934 24168 15990 24177
rect 15934 24103 15990 24112
rect 15752 23860 15804 23866
rect 15752 23802 15804 23808
rect 14832 23180 14884 23186
rect 14832 23122 14884 23128
rect 15476 23180 15528 23186
rect 15476 23122 15528 23128
rect 14740 22704 14792 22710
rect 14740 22646 14792 22652
rect 14648 20528 14700 20534
rect 14648 20470 14700 20476
rect 13636 20392 13688 20398
rect 13636 20334 13688 20340
rect 13820 20256 13872 20262
rect 13820 20198 13872 20204
rect 13832 20058 13860 20198
rect 13452 20052 13504 20058
rect 13452 19994 13504 20000
rect 13820 20052 13872 20058
rect 13820 19994 13872 20000
rect 13912 19848 13964 19854
rect 13912 19790 13964 19796
rect 13636 18760 13688 18766
rect 13636 18702 13688 18708
rect 13452 18692 13504 18698
rect 13452 18634 13504 18640
rect 13268 18420 13320 18426
rect 13268 18362 13320 18368
rect 13176 18284 13228 18290
rect 13176 18226 13228 18232
rect 12768 18040 12940 18068
rect 12992 18080 13044 18086
rect 12716 18022 12768 18028
rect 12992 18022 13044 18028
rect 12072 17876 12124 17882
rect 12072 17818 12124 17824
rect 13004 17762 13032 18022
rect 13188 17882 13216 18226
rect 13280 18204 13308 18362
rect 13464 18290 13492 18634
rect 13648 18290 13676 18702
rect 13452 18284 13504 18290
rect 13452 18226 13504 18232
rect 13636 18284 13688 18290
rect 13636 18226 13688 18232
rect 13360 18216 13412 18222
rect 13280 18176 13360 18204
rect 13360 18158 13412 18164
rect 13648 17882 13676 18226
rect 13176 17876 13228 17882
rect 13176 17818 13228 17824
rect 13636 17876 13688 17882
rect 13636 17818 13688 17824
rect 12728 17734 13032 17762
rect 13924 17746 13952 19790
rect 14004 19780 14056 19786
rect 14004 19722 14056 19728
rect 13912 17740 13964 17746
rect 12728 17610 12756 17734
rect 13912 17682 13964 17688
rect 14016 17610 14044 19722
rect 14660 19378 14688 20470
rect 14844 19786 14872 23122
rect 15014 22808 15070 22817
rect 15014 22743 15070 22752
rect 14924 22432 14976 22438
rect 14924 22374 14976 22380
rect 14936 22166 14964 22374
rect 15028 22166 15056 22743
rect 14924 22160 14976 22166
rect 14924 22102 14976 22108
rect 15016 22160 15068 22166
rect 15016 22102 15068 22108
rect 15028 22030 15056 22102
rect 15016 22024 15068 22030
rect 15016 21966 15068 21972
rect 15016 21888 15068 21894
rect 15016 21830 15068 21836
rect 15028 21554 15056 21830
rect 15488 21554 15516 23122
rect 15568 22228 15620 22234
rect 15568 22170 15620 22176
rect 15016 21548 15068 21554
rect 15016 21490 15068 21496
rect 15476 21548 15528 21554
rect 15476 21490 15528 21496
rect 15108 21480 15160 21486
rect 15108 21422 15160 21428
rect 15120 20330 15148 21422
rect 15580 21418 15608 22170
rect 15764 21962 15792 23802
rect 15948 23322 15976 24103
rect 15936 23316 15988 23322
rect 15936 23258 15988 23264
rect 15936 23112 15988 23118
rect 15936 23054 15988 23060
rect 15948 22710 15976 23054
rect 16040 22778 16068 24754
rect 16120 24744 16172 24750
rect 16118 24712 16120 24721
rect 16172 24712 16174 24721
rect 16118 24647 16174 24656
rect 16132 24410 16160 24647
rect 16120 24404 16172 24410
rect 16120 24346 16172 24352
rect 16868 24274 16896 25162
rect 16856 24268 16908 24274
rect 16856 24210 16908 24216
rect 16580 24064 16632 24070
rect 16580 24006 16632 24012
rect 16592 23866 16620 24006
rect 16580 23860 16632 23866
rect 16580 23802 16632 23808
rect 16592 23474 16620 23802
rect 16960 23730 16988 25638
rect 17132 24812 17184 24818
rect 17052 24772 17132 24800
rect 17052 24342 17080 24772
rect 17132 24754 17184 24760
rect 17224 24812 17276 24818
rect 17224 24754 17276 24760
rect 17132 24676 17184 24682
rect 17132 24618 17184 24624
rect 17040 24336 17092 24342
rect 17040 24278 17092 24284
rect 17144 24206 17172 24618
rect 17236 24410 17264 24754
rect 17316 24744 17368 24750
rect 17316 24686 17368 24692
rect 17328 24410 17356 24686
rect 17224 24404 17276 24410
rect 17224 24346 17276 24352
rect 17316 24404 17368 24410
rect 17316 24346 17368 24352
rect 17132 24200 17184 24206
rect 17132 24142 17184 24148
rect 16948 23724 17000 23730
rect 16948 23666 17000 23672
rect 16500 23446 16620 23474
rect 16500 23050 16528 23446
rect 16960 23322 16988 23666
rect 17420 23497 17448 25638
rect 17512 24750 17540 25774
rect 17776 25764 17828 25770
rect 17776 25706 17828 25712
rect 18420 25764 18472 25770
rect 18420 25706 18472 25712
rect 17592 25152 17644 25158
rect 17592 25094 17644 25100
rect 17604 24886 17632 25094
rect 17592 24880 17644 24886
rect 17592 24822 17644 24828
rect 17500 24744 17552 24750
rect 17500 24686 17552 24692
rect 17406 23488 17462 23497
rect 17406 23423 17462 23432
rect 16672 23316 16724 23322
rect 16672 23258 16724 23264
rect 16948 23316 17000 23322
rect 16948 23258 17000 23264
rect 16488 23044 16540 23050
rect 16488 22986 16540 22992
rect 16028 22772 16080 22778
rect 16028 22714 16080 22720
rect 16304 22772 16356 22778
rect 16304 22714 16356 22720
rect 15936 22704 15988 22710
rect 15936 22646 15988 22652
rect 15948 22438 15976 22646
rect 15936 22432 15988 22438
rect 15936 22374 15988 22380
rect 16212 22160 16264 22166
rect 16212 22102 16264 22108
rect 16028 22024 16080 22030
rect 16028 21966 16080 21972
rect 15660 21956 15712 21962
rect 15660 21898 15712 21904
rect 15752 21956 15804 21962
rect 15752 21898 15804 21904
rect 15672 21622 15700 21898
rect 15660 21616 15712 21622
rect 15660 21558 15712 21564
rect 15568 21412 15620 21418
rect 15568 21354 15620 21360
rect 15580 20602 15608 21354
rect 15764 20942 15792 21898
rect 16040 21690 16068 21966
rect 16028 21684 16080 21690
rect 16028 21626 16080 21632
rect 15752 20936 15804 20942
rect 15752 20878 15804 20884
rect 16028 20936 16080 20942
rect 16028 20878 16080 20884
rect 15844 20868 15896 20874
rect 15844 20810 15896 20816
rect 15568 20596 15620 20602
rect 15568 20538 15620 20544
rect 15580 20466 15608 20538
rect 15856 20534 15884 20810
rect 15936 20596 15988 20602
rect 15936 20538 15988 20544
rect 15844 20528 15896 20534
rect 15844 20470 15896 20476
rect 15568 20460 15620 20466
rect 15568 20402 15620 20408
rect 15660 20392 15712 20398
rect 15660 20334 15712 20340
rect 15108 20324 15160 20330
rect 15108 20266 15160 20272
rect 14832 19780 14884 19786
rect 14832 19722 14884 19728
rect 15120 19378 15148 20266
rect 14648 19372 14700 19378
rect 14648 19314 14700 19320
rect 15108 19372 15160 19378
rect 15108 19314 15160 19320
rect 15120 18698 15148 19314
rect 15200 19304 15252 19310
rect 15200 19246 15252 19252
rect 15212 18970 15240 19246
rect 15200 18964 15252 18970
rect 15200 18906 15252 18912
rect 15108 18692 15160 18698
rect 15108 18634 15160 18640
rect 15120 18426 15148 18634
rect 15108 18420 15160 18426
rect 15108 18362 15160 18368
rect 14740 17876 14792 17882
rect 14740 17818 14792 17824
rect 14752 17610 14780 17818
rect 11336 17604 11388 17610
rect 11336 17546 11388 17552
rect 12716 17604 12768 17610
rect 12716 17546 12768 17552
rect 14004 17604 14056 17610
rect 14004 17546 14056 17552
rect 14740 17604 14792 17610
rect 14740 17546 14792 17552
rect 11152 17332 11204 17338
rect 11152 17274 11204 17280
rect 11348 17202 11376 17546
rect 15212 17542 15240 18906
rect 15672 18902 15700 20334
rect 15856 19922 15884 20470
rect 15948 20466 15976 20538
rect 15936 20460 15988 20466
rect 15936 20402 15988 20408
rect 15936 20256 15988 20262
rect 15936 20198 15988 20204
rect 15948 19990 15976 20198
rect 15936 19984 15988 19990
rect 15936 19926 15988 19932
rect 15844 19916 15896 19922
rect 15844 19858 15896 19864
rect 15844 19168 15896 19174
rect 15844 19110 15896 19116
rect 15752 18964 15804 18970
rect 15752 18906 15804 18912
rect 15660 18896 15712 18902
rect 15660 18838 15712 18844
rect 15672 18358 15700 18838
rect 15764 18766 15792 18906
rect 15752 18760 15804 18766
rect 15752 18702 15804 18708
rect 15856 18698 15884 19110
rect 15936 18964 15988 18970
rect 15936 18906 15988 18912
rect 15844 18692 15896 18698
rect 15844 18634 15896 18640
rect 15476 18352 15528 18358
rect 15660 18352 15712 18358
rect 15528 18312 15608 18340
rect 15476 18294 15528 18300
rect 15580 17882 15608 18312
rect 15660 18294 15712 18300
rect 15568 17876 15620 17882
rect 15568 17818 15620 17824
rect 15580 17610 15608 17818
rect 15568 17604 15620 17610
rect 15568 17546 15620 17552
rect 15200 17536 15252 17542
rect 15200 17478 15252 17484
rect 15948 17270 15976 18906
rect 16040 18766 16068 20878
rect 16224 20602 16252 22102
rect 16316 22030 16344 22714
rect 16500 22030 16528 22986
rect 16304 22024 16356 22030
rect 16304 21966 16356 21972
rect 16488 22024 16540 22030
rect 16488 21966 16540 21972
rect 16396 21956 16448 21962
rect 16396 21898 16448 21904
rect 16304 21548 16356 21554
rect 16304 21490 16356 21496
rect 16316 20806 16344 21490
rect 16408 21010 16436 21898
rect 16684 21554 16712 23258
rect 16764 23248 16816 23254
rect 16764 23190 16816 23196
rect 16776 22642 16804 23190
rect 17408 23112 17460 23118
rect 17408 23054 17460 23060
rect 17132 22976 17184 22982
rect 17132 22918 17184 22924
rect 16764 22636 16816 22642
rect 16764 22578 16816 22584
rect 16764 22500 16816 22506
rect 16764 22442 16816 22448
rect 16776 21554 16804 22442
rect 17144 22234 17172 22918
rect 17420 22778 17448 23054
rect 17408 22772 17460 22778
rect 17408 22714 17460 22720
rect 17512 22710 17540 24686
rect 17604 24206 17632 24822
rect 17788 24818 17816 25706
rect 17868 24880 17920 24886
rect 18432 24857 18460 25706
rect 19524 25356 19576 25362
rect 19524 25298 19576 25304
rect 19432 25220 19484 25226
rect 19432 25162 19484 25168
rect 18418 24848 18474 24857
rect 17920 24828 18184 24834
rect 17868 24822 18184 24828
rect 17880 24818 18184 24822
rect 17776 24812 17828 24818
rect 17880 24812 18196 24818
rect 17880 24806 18144 24812
rect 17776 24754 17828 24760
rect 19444 24818 19472 25162
rect 18418 24783 18474 24792
rect 19432 24812 19484 24818
rect 18144 24754 18196 24760
rect 17684 24744 17736 24750
rect 17684 24686 17736 24692
rect 17592 24200 17644 24206
rect 17592 24142 17644 24148
rect 17500 22704 17552 22710
rect 17500 22646 17552 22652
rect 17604 22506 17632 24142
rect 17696 24138 17724 24686
rect 17684 24132 17736 24138
rect 17684 24074 17736 24080
rect 17788 24070 17816 24754
rect 17960 24132 18012 24138
rect 17960 24074 18012 24080
rect 17776 24064 17828 24070
rect 17972 24018 18000 24074
rect 17776 24006 17828 24012
rect 17788 23798 17816 24006
rect 17880 23990 18000 24018
rect 17880 23798 17908 23990
rect 17776 23792 17828 23798
rect 17776 23734 17828 23740
rect 17868 23792 17920 23798
rect 17868 23734 17920 23740
rect 17788 23594 17816 23734
rect 17684 23588 17736 23594
rect 17684 23530 17736 23536
rect 17776 23588 17828 23594
rect 17776 23530 17828 23536
rect 17696 23118 17724 23530
rect 17880 23118 17908 23734
rect 18432 23594 18460 24783
rect 19432 24754 19484 24760
rect 19536 24750 19564 25298
rect 24860 25288 24912 25294
rect 24858 25256 24860 25265
rect 24912 25256 24914 25265
rect 21088 25220 21140 25226
rect 24858 25191 24914 25200
rect 21088 25162 21140 25168
rect 20996 25152 21048 25158
rect 20996 25094 21048 25100
rect 19892 24948 19944 24954
rect 19892 24890 19944 24896
rect 19340 24744 19392 24750
rect 19340 24686 19392 24692
rect 19524 24744 19576 24750
rect 19524 24686 19576 24692
rect 19800 24744 19852 24750
rect 19800 24686 19852 24692
rect 18880 24404 18932 24410
rect 18880 24346 18932 24352
rect 19076 24398 19288 24426
rect 18604 24064 18656 24070
rect 18604 24006 18656 24012
rect 18512 23656 18564 23662
rect 18512 23598 18564 23604
rect 18420 23588 18472 23594
rect 18420 23530 18472 23536
rect 18328 23520 18380 23526
rect 18328 23462 18380 23468
rect 17684 23112 17736 23118
rect 17684 23054 17736 23060
rect 17868 23112 17920 23118
rect 17868 23054 17920 23060
rect 17960 22976 18012 22982
rect 17960 22918 18012 22924
rect 17592 22500 17644 22506
rect 17592 22442 17644 22448
rect 17972 22234 18000 22918
rect 17132 22228 17184 22234
rect 17132 22170 17184 22176
rect 17960 22228 18012 22234
rect 17960 22170 18012 22176
rect 18236 22160 18288 22166
rect 18236 22102 18288 22108
rect 17960 22024 18012 22030
rect 17960 21966 18012 21972
rect 17776 21956 17828 21962
rect 17776 21898 17828 21904
rect 17500 21888 17552 21894
rect 17500 21830 17552 21836
rect 16672 21548 16724 21554
rect 16672 21490 16724 21496
rect 16764 21548 16816 21554
rect 16764 21490 16816 21496
rect 16948 21548 17000 21554
rect 16948 21490 17000 21496
rect 17040 21548 17092 21554
rect 17040 21490 17092 21496
rect 17132 21548 17184 21554
rect 17132 21490 17184 21496
rect 16960 21078 16988 21490
rect 16948 21072 17000 21078
rect 16948 21014 17000 21020
rect 16396 21004 16448 21010
rect 16396 20946 16448 20952
rect 16304 20800 16356 20806
rect 16304 20742 16356 20748
rect 16212 20596 16264 20602
rect 16212 20538 16264 20544
rect 16212 19508 16264 19514
rect 16212 19450 16264 19456
rect 16120 18828 16172 18834
rect 16120 18770 16172 18776
rect 16028 18760 16080 18766
rect 16028 18702 16080 18708
rect 16132 17610 16160 18770
rect 16120 17604 16172 17610
rect 16120 17546 16172 17552
rect 15936 17264 15988 17270
rect 15936 17206 15988 17212
rect 11336 17196 11388 17202
rect 11336 17138 11388 17144
rect 10048 16788 10100 16794
rect 10048 16730 10100 16736
rect 10600 16040 10652 16046
rect 10600 15982 10652 15988
rect 10140 15904 10192 15910
rect 10140 15846 10192 15852
rect 10152 15570 10180 15846
rect 10612 15706 10640 15982
rect 10600 15700 10652 15706
rect 10600 15642 10652 15648
rect 9588 15564 9640 15570
rect 9588 15506 9640 15512
rect 10140 15564 10192 15570
rect 10140 15506 10192 15512
rect 9312 15496 9364 15502
rect 9312 15438 9364 15444
rect 9220 15360 9272 15366
rect 9220 15302 9272 15308
rect 8944 14884 8996 14890
rect 8944 14826 8996 14832
rect 8116 14408 8168 14414
rect 8116 14350 8168 14356
rect 8128 13938 8156 14350
rect 8208 14068 8260 14074
rect 8208 14010 8260 14016
rect 8116 13932 8168 13938
rect 8116 13874 8168 13880
rect 7748 13864 7800 13870
rect 7748 13806 7800 13812
rect 8220 13258 8248 14010
rect 8392 13864 8444 13870
rect 8392 13806 8444 13812
rect 8484 13864 8536 13870
rect 8484 13806 8536 13812
rect 8404 13462 8432 13806
rect 8496 13530 8524 13806
rect 8484 13524 8536 13530
rect 8484 13466 8536 13472
rect 8392 13456 8444 13462
rect 8392 13398 8444 13404
rect 8208 13252 8260 13258
rect 8208 13194 8260 13200
rect 7668 12406 7880 12434
rect 7104 12164 7156 12170
rect 7104 12106 7156 12112
rect 6920 11688 6972 11694
rect 6920 11630 6972 11636
rect 6368 11212 6420 11218
rect 6368 11154 6420 11160
rect 6828 11212 6880 11218
rect 6828 11154 6880 11160
rect 6276 11144 6328 11150
rect 6276 11086 6328 11092
rect 6840 11098 6868 11154
rect 5724 11076 5776 11082
rect 6840 11070 6960 11098
rect 5724 11018 5776 11024
rect 6932 10674 6960 11070
rect 6920 10668 6972 10674
rect 6920 10610 6972 10616
rect 5356 10464 5408 10470
rect 5356 10406 5408 10412
rect 5264 10260 5316 10266
rect 5264 10202 5316 10208
rect 4804 10192 4856 10198
rect 4804 10134 4856 10140
rect 4894 10160 4950 10169
rect 4710 10024 4766 10033
rect 4710 9959 4766 9968
rect 4712 9920 4764 9926
rect 4712 9862 4764 9868
rect 4724 8974 4752 9862
rect 4816 9586 4844 10134
rect 4894 10095 4950 10104
rect 4908 9926 4936 10095
rect 4896 9920 4948 9926
rect 4896 9862 4948 9868
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 5368 9722 5396 10406
rect 6092 10192 6144 10198
rect 6092 10134 6144 10140
rect 5448 10056 5500 10062
rect 5448 9998 5500 10004
rect 4896 9716 4948 9722
rect 4896 9658 4948 9664
rect 5356 9716 5408 9722
rect 5356 9658 5408 9664
rect 4804 9580 4856 9586
rect 4804 9522 4856 9528
rect 4804 9444 4856 9450
rect 4804 9386 4856 9392
rect 4816 9178 4844 9386
rect 4804 9172 4856 9178
rect 4804 9114 4856 9120
rect 4908 9058 4936 9658
rect 5170 9616 5226 9625
rect 5170 9551 5172 9560
rect 5224 9551 5226 9560
rect 5264 9580 5316 9586
rect 5172 9522 5224 9528
rect 5264 9522 5316 9528
rect 4816 9042 4936 9058
rect 4804 9036 4936 9042
rect 4856 9030 4936 9036
rect 4804 8978 4856 8984
rect 5276 8974 5304 9522
rect 5460 9450 5488 9998
rect 5540 9648 5592 9654
rect 5540 9590 5592 9596
rect 5448 9444 5500 9450
rect 5448 9386 5500 9392
rect 4712 8968 4764 8974
rect 4712 8910 4764 8916
rect 5264 8968 5316 8974
rect 5264 8910 5316 8916
rect 5356 8968 5408 8974
rect 5356 8910 5408 8916
rect 4804 8900 4856 8906
rect 4804 8842 4856 8848
rect 4710 8664 4766 8673
rect 4816 8634 4844 8842
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 5276 8634 5304 8910
rect 4710 8599 4766 8608
rect 4804 8628 4856 8634
rect 4724 8430 4752 8599
rect 4804 8570 4856 8576
rect 5264 8628 5316 8634
rect 5264 8570 5316 8576
rect 5078 8528 5134 8537
rect 4804 8492 4856 8498
rect 5078 8463 5134 8472
rect 5172 8492 5224 8498
rect 4804 8434 4856 8440
rect 4712 8424 4764 8430
rect 4710 8392 4712 8401
rect 4764 8392 4766 8401
rect 4710 8327 4766 8336
rect 4712 7812 4764 7818
rect 4712 7754 4764 7760
rect 4724 7002 4752 7754
rect 4816 7324 4844 8434
rect 4896 8356 4948 8362
rect 4896 8298 4948 8304
rect 4908 7954 4936 8298
rect 4896 7948 4948 7954
rect 4896 7890 4948 7896
rect 5092 7868 5120 8463
rect 5172 8434 5224 8440
rect 5264 8492 5316 8498
rect 5264 8434 5316 8440
rect 5184 8294 5212 8434
rect 5172 8288 5224 8294
rect 5172 8230 5224 8236
rect 5184 7993 5212 8230
rect 5276 8022 5304 8434
rect 5264 8016 5316 8022
rect 5170 7984 5226 7993
rect 5264 7958 5316 7964
rect 5170 7919 5226 7928
rect 5092 7840 5304 7868
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 5276 7546 5304 7840
rect 5368 7546 5396 8910
rect 5460 7886 5488 9386
rect 5552 9110 5580 9590
rect 5908 9376 5960 9382
rect 5908 9318 5960 9324
rect 5540 9104 5592 9110
rect 5540 9046 5592 9052
rect 5632 9036 5684 9042
rect 5632 8978 5684 8984
rect 5724 9036 5776 9042
rect 5724 8978 5776 8984
rect 5540 8968 5592 8974
rect 5540 8910 5592 8916
rect 5552 8498 5580 8910
rect 5540 8492 5592 8498
rect 5540 8434 5592 8440
rect 5644 8294 5672 8978
rect 5736 8498 5764 8978
rect 5920 8906 5948 9318
rect 6104 9178 6132 10134
rect 6932 10130 6960 10610
rect 6920 10124 6972 10130
rect 6920 10066 6972 10072
rect 6552 10056 6604 10062
rect 6552 9998 6604 10004
rect 6564 9722 6592 9998
rect 6644 9988 6696 9994
rect 6644 9930 6696 9936
rect 6552 9716 6604 9722
rect 6552 9658 6604 9664
rect 6460 9648 6512 9654
rect 6460 9590 6512 9596
rect 6368 9580 6420 9586
rect 6368 9522 6420 9528
rect 6276 9512 6328 9518
rect 6276 9454 6328 9460
rect 6288 9178 6316 9454
rect 6092 9172 6144 9178
rect 6092 9114 6144 9120
rect 6276 9172 6328 9178
rect 6276 9114 6328 9120
rect 5908 8900 5960 8906
rect 5908 8842 5960 8848
rect 5724 8492 5776 8498
rect 5724 8434 5776 8440
rect 5736 8401 5764 8434
rect 5722 8392 5778 8401
rect 6380 8362 6408 9522
rect 5722 8327 5778 8336
rect 6368 8356 6420 8362
rect 5632 8288 5684 8294
rect 5632 8230 5684 8236
rect 5736 7954 5764 8327
rect 6368 8298 6420 8304
rect 6380 8022 6408 8298
rect 6368 8016 6420 8022
rect 6368 7958 6420 7964
rect 5724 7948 5776 7954
rect 5724 7890 5776 7896
rect 5448 7880 5500 7886
rect 5448 7822 5500 7828
rect 5448 7744 5500 7750
rect 5448 7686 5500 7692
rect 5908 7744 5960 7750
rect 5908 7686 5960 7692
rect 5264 7540 5316 7546
rect 5264 7482 5316 7488
rect 5356 7540 5408 7546
rect 5356 7482 5408 7488
rect 5172 7472 5224 7478
rect 5224 7420 5304 7426
rect 5172 7414 5304 7420
rect 5184 7398 5304 7414
rect 4896 7336 4948 7342
rect 4816 7296 4896 7324
rect 4896 7278 4948 7284
rect 5078 7304 5134 7313
rect 4908 7002 4936 7278
rect 4988 7268 5040 7274
rect 5078 7239 5134 7248
rect 4988 7210 5040 7216
rect 4712 6996 4764 7002
rect 4712 6938 4764 6944
rect 4896 6996 4948 7002
rect 4896 6938 4948 6944
rect 4896 6860 4948 6866
rect 5000 6848 5028 7210
rect 5092 7002 5120 7239
rect 5080 6996 5132 7002
rect 5080 6938 5132 6944
rect 5276 6866 5304 7398
rect 5356 7404 5408 7410
rect 5356 7346 5408 7352
rect 4948 6820 5028 6848
rect 5264 6860 5316 6866
rect 4896 6802 4948 6808
rect 5264 6802 5316 6808
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 4620 5772 4672 5778
rect 4620 5714 4672 5720
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 5276 5370 5304 6802
rect 5368 6798 5396 7346
rect 5356 6792 5408 6798
rect 5356 6734 5408 6740
rect 5368 5914 5396 6734
rect 5460 6458 5488 7686
rect 5920 7410 5948 7686
rect 5908 7404 5960 7410
rect 5908 7346 5960 7352
rect 6000 7200 6052 7206
rect 6000 7142 6052 7148
rect 6012 6458 6040 7142
rect 5448 6452 5500 6458
rect 5448 6394 5500 6400
rect 6000 6452 6052 6458
rect 6000 6394 6052 6400
rect 6472 6254 6500 9590
rect 6564 7410 6592 9658
rect 6656 9518 6684 9930
rect 6932 9654 6960 10066
rect 7012 9920 7064 9926
rect 7012 9862 7064 9868
rect 6920 9648 6972 9654
rect 6920 9590 6972 9596
rect 6644 9512 6696 9518
rect 6644 9454 6696 9460
rect 6656 9110 6684 9454
rect 6644 9104 6696 9110
rect 6644 9046 6696 9052
rect 6736 8900 6788 8906
rect 6736 8842 6788 8848
rect 6748 7886 6776 8842
rect 6932 8498 6960 9590
rect 6920 8492 6972 8498
rect 6920 8434 6972 8440
rect 6920 8016 6972 8022
rect 6920 7958 6972 7964
rect 6932 7886 6960 7958
rect 6736 7880 6788 7886
rect 6736 7822 6788 7828
rect 6920 7880 6972 7886
rect 6920 7822 6972 7828
rect 6736 7744 6788 7750
rect 6736 7686 6788 7692
rect 6748 7478 6776 7686
rect 6736 7472 6788 7478
rect 6736 7414 6788 7420
rect 6552 7404 6604 7410
rect 6552 7346 6604 7352
rect 6564 6662 6592 7346
rect 7024 6866 7052 9862
rect 7116 9674 7144 12106
rect 7852 11694 7880 12406
rect 7840 11688 7892 11694
rect 7840 11630 7892 11636
rect 7288 11552 7340 11558
rect 7288 11494 7340 11500
rect 7300 11218 7328 11494
rect 7288 11212 7340 11218
rect 7288 11154 7340 11160
rect 7748 10600 7800 10606
rect 7748 10542 7800 10548
rect 7116 9646 7328 9674
rect 7300 8906 7328 9646
rect 7760 9450 7788 10542
rect 7748 9444 7800 9450
rect 7748 9386 7800 9392
rect 7288 8900 7340 8906
rect 7116 8860 7288 8888
rect 7012 6860 7064 6866
rect 7012 6802 7064 6808
rect 6828 6724 6880 6730
rect 6828 6666 6880 6672
rect 6552 6656 6604 6662
rect 6552 6598 6604 6604
rect 6840 6458 6868 6666
rect 6828 6452 6880 6458
rect 6828 6394 6880 6400
rect 6460 6248 6512 6254
rect 6460 6190 6512 6196
rect 6552 6112 6604 6118
rect 6552 6054 6604 6060
rect 5356 5908 5408 5914
rect 5356 5850 5408 5856
rect 6564 5778 6592 6054
rect 6552 5772 6604 5778
rect 6552 5714 6604 5720
rect 6092 5636 6144 5642
rect 6092 5578 6144 5584
rect 7012 5636 7064 5642
rect 7116 5624 7144 8860
rect 7288 8842 7340 8848
rect 7380 8832 7432 8838
rect 7380 8774 7432 8780
rect 7392 8498 7420 8774
rect 7288 8492 7340 8498
rect 7288 8434 7340 8440
rect 7380 8492 7432 8498
rect 7380 8434 7432 8440
rect 7196 8288 7248 8294
rect 7196 8230 7248 8236
rect 7208 7886 7236 8230
rect 7300 7886 7328 8434
rect 7196 7880 7248 7886
rect 7196 7822 7248 7828
rect 7288 7880 7340 7886
rect 7288 7822 7340 7828
rect 7380 7744 7432 7750
rect 7380 7686 7432 7692
rect 7392 7546 7420 7686
rect 7380 7540 7432 7546
rect 7380 7482 7432 7488
rect 7852 6798 7880 11630
rect 8024 9648 8076 9654
rect 8024 9590 8076 9596
rect 7932 9376 7984 9382
rect 7932 9318 7984 9324
rect 7944 8906 7972 9318
rect 8036 9042 8064 9590
rect 8024 9036 8076 9042
rect 8024 8978 8076 8984
rect 7932 8900 7984 8906
rect 7932 8842 7984 8848
rect 8036 8634 8064 8978
rect 8024 8628 8076 8634
rect 8024 8570 8076 8576
rect 8036 6798 8064 8570
rect 8220 8566 8248 13194
rect 8668 12096 8720 12102
rect 8668 12038 8720 12044
rect 8300 11892 8352 11898
rect 8300 11834 8352 11840
rect 8312 11082 8340 11834
rect 8680 11762 8708 12038
rect 8668 11756 8720 11762
rect 8668 11698 8720 11704
rect 8680 11354 8708 11698
rect 8484 11348 8536 11354
rect 8484 11290 8536 11296
rect 8668 11348 8720 11354
rect 8668 11290 8720 11296
rect 8300 11076 8352 11082
rect 8300 11018 8352 11024
rect 8312 10742 8340 11018
rect 8300 10736 8352 10742
rect 8300 10678 8352 10684
rect 8496 9518 8524 11290
rect 8956 10810 8984 14826
rect 9232 14822 9260 15302
rect 9220 14816 9272 14822
rect 9220 14758 9272 14764
rect 9128 12640 9180 12646
rect 9128 12582 9180 12588
rect 9140 12306 9168 12582
rect 9232 12434 9260 14758
rect 9324 14346 9352 15438
rect 9680 15360 9732 15366
rect 9680 15302 9732 15308
rect 9692 15026 9720 15302
rect 9680 15020 9732 15026
rect 9680 14962 9732 14968
rect 9680 14408 9732 14414
rect 9680 14350 9732 14356
rect 9312 14340 9364 14346
rect 9312 14282 9364 14288
rect 9692 14074 9720 14350
rect 10140 14340 10192 14346
rect 10140 14282 10192 14288
rect 9680 14068 9732 14074
rect 9680 14010 9732 14016
rect 9864 13728 9916 13734
rect 9864 13670 9916 13676
rect 9404 13388 9456 13394
rect 9404 13330 9456 13336
rect 9772 13388 9824 13394
rect 9772 13330 9824 13336
rect 9232 12406 9352 12434
rect 9128 12300 9180 12306
rect 9128 12242 9180 12248
rect 9220 12232 9272 12238
rect 9220 12174 9272 12180
rect 9232 11762 9260 12174
rect 9220 11756 9272 11762
rect 9220 11698 9272 11704
rect 8944 10804 8996 10810
rect 8944 10746 8996 10752
rect 9036 10804 9088 10810
rect 9036 10746 9088 10752
rect 8956 10062 8984 10746
rect 8944 10056 8996 10062
rect 8944 9998 8996 10004
rect 9048 9722 9076 10746
rect 9324 10130 9352 12406
rect 9312 10124 9364 10130
rect 9312 10066 9364 10072
rect 9312 9920 9364 9926
rect 9312 9862 9364 9868
rect 9036 9716 9088 9722
rect 9036 9658 9088 9664
rect 8484 9512 8536 9518
rect 8484 9454 8536 9460
rect 8208 8560 8260 8566
rect 8208 8502 8260 8508
rect 8300 7200 8352 7206
rect 8300 7142 8352 7148
rect 7840 6792 7892 6798
rect 7840 6734 7892 6740
rect 8024 6792 8076 6798
rect 8024 6734 8076 6740
rect 7288 6656 7340 6662
rect 7288 6598 7340 6604
rect 7564 6656 7616 6662
rect 7564 6598 7616 6604
rect 7300 5710 7328 6598
rect 7576 5914 7604 6598
rect 8036 6322 8064 6734
rect 8116 6656 8168 6662
rect 8116 6598 8168 6604
rect 8128 6322 8156 6598
rect 8024 6316 8076 6322
rect 8024 6258 8076 6264
rect 8116 6316 8168 6322
rect 8116 6258 8168 6264
rect 7564 5908 7616 5914
rect 7564 5850 7616 5856
rect 8036 5778 8064 6258
rect 8024 5772 8076 5778
rect 8024 5714 8076 5720
rect 7288 5704 7340 5710
rect 7288 5646 7340 5652
rect 7064 5596 7144 5624
rect 7012 5578 7064 5584
rect 5264 5364 5316 5370
rect 5264 5306 5316 5312
rect 6104 5302 6132 5578
rect 3884 5296 3936 5302
rect 3884 5238 3936 5244
rect 6092 5296 6144 5302
rect 6092 5238 6144 5244
rect 3700 5228 3752 5234
rect 3700 5170 3752 5176
rect 2872 5160 2924 5166
rect 2872 5102 2924 5108
rect 7116 5030 7144 5596
rect 8036 5234 8064 5714
rect 8312 5234 8340 7142
rect 8496 6866 8524 9454
rect 8852 8900 8904 8906
rect 8852 8842 8904 8848
rect 8864 8566 8892 8842
rect 8852 8560 8904 8566
rect 8852 8502 8904 8508
rect 9324 8498 9352 9862
rect 9312 8492 9364 8498
rect 9312 8434 9364 8440
rect 9416 7546 9444 13330
rect 9784 12782 9812 13330
rect 9876 13190 9904 13670
rect 9864 13184 9916 13190
rect 9864 13126 9916 13132
rect 9588 12776 9640 12782
rect 9588 12718 9640 12724
rect 9772 12776 9824 12782
rect 9772 12718 9824 12724
rect 9600 12442 9628 12718
rect 9588 12436 9640 12442
rect 9784 12434 9812 12718
rect 9784 12406 9904 12434
rect 9588 12378 9640 12384
rect 9600 9110 9628 12378
rect 9680 12164 9732 12170
rect 9680 12106 9732 12112
rect 9692 11898 9720 12106
rect 9680 11892 9732 11898
rect 9680 11834 9732 11840
rect 9772 11688 9824 11694
rect 9772 11630 9824 11636
rect 9784 11354 9812 11630
rect 9876 11558 9904 12406
rect 10152 11898 10180 14282
rect 10416 14272 10468 14278
rect 10416 14214 10468 14220
rect 10428 14074 10456 14214
rect 10416 14068 10468 14074
rect 10416 14010 10468 14016
rect 10508 13864 10560 13870
rect 10508 13806 10560 13812
rect 10140 11892 10192 11898
rect 10140 11834 10192 11840
rect 9864 11552 9916 11558
rect 9864 11494 9916 11500
rect 9772 11348 9824 11354
rect 9772 11290 9824 11296
rect 10152 11286 10180 11834
rect 10324 11552 10376 11558
rect 10324 11494 10376 11500
rect 10140 11280 10192 11286
rect 10140 11222 10192 11228
rect 10336 11218 10364 11494
rect 10324 11212 10376 11218
rect 10324 11154 10376 11160
rect 10324 11076 10376 11082
rect 10324 11018 10376 11024
rect 9680 10056 9732 10062
rect 9680 9998 9732 10004
rect 9588 9104 9640 9110
rect 9588 9046 9640 9052
rect 9692 9042 9720 9998
rect 10140 9920 10192 9926
rect 10140 9862 10192 9868
rect 9680 9036 9732 9042
rect 9680 8978 9732 8984
rect 9692 7886 9720 8978
rect 10152 8498 10180 9862
rect 10232 9648 10284 9654
rect 10232 9590 10284 9596
rect 10244 9178 10272 9590
rect 10232 9172 10284 9178
rect 10232 9114 10284 9120
rect 10140 8492 10192 8498
rect 10140 8434 10192 8440
rect 10244 8430 10272 9114
rect 10232 8424 10284 8430
rect 10232 8366 10284 8372
rect 9680 7880 9732 7886
rect 9680 7822 9732 7828
rect 9404 7540 9456 7546
rect 9404 7482 9456 7488
rect 9692 7342 9720 7822
rect 9864 7404 9916 7410
rect 9864 7346 9916 7352
rect 10140 7404 10192 7410
rect 10140 7346 10192 7352
rect 9680 7336 9732 7342
rect 9680 7278 9732 7284
rect 9588 6996 9640 7002
rect 9692 6984 9720 7278
rect 9772 7200 9824 7206
rect 9772 7142 9824 7148
rect 9640 6956 9720 6984
rect 9588 6938 9640 6944
rect 9784 6866 9812 7142
rect 8484 6860 8536 6866
rect 8484 6802 8536 6808
rect 9772 6860 9824 6866
rect 9772 6802 9824 6808
rect 9588 6656 9640 6662
rect 9588 6598 9640 6604
rect 9600 6390 9628 6598
rect 9588 6384 9640 6390
rect 9876 6361 9904 7346
rect 10152 7002 10180 7346
rect 10140 6996 10192 7002
rect 10140 6938 10192 6944
rect 10140 6724 10192 6730
rect 10244 6712 10272 8366
rect 10336 7546 10364 11018
rect 10520 10130 10548 13806
rect 10612 13802 10640 15642
rect 10968 15496 11020 15502
rect 10968 15438 11020 15444
rect 10692 15360 10744 15366
rect 10692 15302 10744 15308
rect 10784 15360 10836 15366
rect 10784 15302 10836 15308
rect 10704 15026 10732 15302
rect 10796 15094 10824 15302
rect 10980 15178 11008 15438
rect 11348 15434 11376 17138
rect 16132 17066 16160 17546
rect 16120 17060 16172 17066
rect 16120 17002 16172 17008
rect 16224 16998 16252 19450
rect 16316 18222 16344 20742
rect 16408 19378 16436 20946
rect 16764 20936 16816 20942
rect 16764 20878 16816 20884
rect 16672 20324 16724 20330
rect 16672 20266 16724 20272
rect 16684 19786 16712 20266
rect 16672 19780 16724 19786
rect 16672 19722 16724 19728
rect 16684 19446 16712 19722
rect 16672 19440 16724 19446
rect 16672 19382 16724 19388
rect 16396 19372 16448 19378
rect 16396 19314 16448 19320
rect 16408 18290 16436 19314
rect 16684 18630 16712 19382
rect 16672 18624 16724 18630
rect 16672 18566 16724 18572
rect 16684 18358 16712 18566
rect 16672 18352 16724 18358
rect 16672 18294 16724 18300
rect 16396 18284 16448 18290
rect 16396 18226 16448 18232
rect 16304 18216 16356 18222
rect 16304 18158 16356 18164
rect 16316 17746 16344 18158
rect 16304 17740 16356 17746
rect 16304 17682 16356 17688
rect 16316 17202 16344 17682
rect 16580 17604 16632 17610
rect 16580 17546 16632 17552
rect 16396 17536 16448 17542
rect 16396 17478 16448 17484
rect 16408 17270 16436 17478
rect 16396 17264 16448 17270
rect 16396 17206 16448 17212
rect 16304 17196 16356 17202
rect 16304 17138 16356 17144
rect 16592 17134 16620 17546
rect 16580 17128 16632 17134
rect 16580 17070 16632 17076
rect 16212 16992 16264 16998
rect 16212 16934 16264 16940
rect 11980 16176 12032 16182
rect 11980 16118 12032 16124
rect 11336 15428 11388 15434
rect 11336 15370 11388 15376
rect 10888 15150 11008 15178
rect 10784 15088 10836 15094
rect 10784 15030 10836 15036
rect 10692 15020 10744 15026
rect 10692 14962 10744 14968
rect 10600 13796 10652 13802
rect 10600 13738 10652 13744
rect 10612 13394 10640 13738
rect 10600 13388 10652 13394
rect 10600 13330 10652 13336
rect 10692 12844 10744 12850
rect 10692 12786 10744 12792
rect 10704 12442 10732 12786
rect 10692 12436 10744 12442
rect 10692 12378 10744 12384
rect 10888 11098 10916 15150
rect 11520 15020 11572 15026
rect 11520 14962 11572 14968
rect 11532 14414 11560 14962
rect 11704 14952 11756 14958
rect 11704 14894 11756 14900
rect 11520 14408 11572 14414
rect 11520 14350 11572 14356
rect 11612 14408 11664 14414
rect 11612 14350 11664 14356
rect 11428 14340 11480 14346
rect 11428 14282 11480 14288
rect 11336 13796 11388 13802
rect 11336 13738 11388 13744
rect 11348 12238 11376 13738
rect 11440 13326 11468 14282
rect 11428 13320 11480 13326
rect 11428 13262 11480 13268
rect 11440 12238 11468 13262
rect 11532 13258 11560 14350
rect 11520 13252 11572 13258
rect 11520 13194 11572 13200
rect 11532 12238 11560 13194
rect 11624 13190 11652 14350
rect 11716 13938 11744 14894
rect 11796 14340 11848 14346
rect 11796 14282 11848 14288
rect 11704 13932 11756 13938
rect 11704 13874 11756 13880
rect 11716 13530 11744 13874
rect 11704 13524 11756 13530
rect 11704 13466 11756 13472
rect 11808 13462 11836 14282
rect 11796 13456 11848 13462
rect 11796 13398 11848 13404
rect 11612 13184 11664 13190
rect 11612 13126 11664 13132
rect 11624 12306 11652 13126
rect 11612 12300 11664 12306
rect 11612 12242 11664 12248
rect 11336 12232 11388 12238
rect 11336 12174 11388 12180
rect 11428 12232 11480 12238
rect 11428 12174 11480 12180
rect 11520 12232 11572 12238
rect 11520 12174 11572 12180
rect 11440 11830 11468 12174
rect 11532 11898 11560 12174
rect 11520 11892 11572 11898
rect 11520 11834 11572 11840
rect 11428 11824 11480 11830
rect 11428 11766 11480 11772
rect 10704 11082 10916 11098
rect 11440 11082 11468 11766
rect 11624 11762 11652 12242
rect 11612 11756 11664 11762
rect 11612 11698 11664 11704
rect 11624 11286 11652 11698
rect 11612 11280 11664 11286
rect 11612 11222 11664 11228
rect 10692 11076 10916 11082
rect 10744 11070 10916 11076
rect 11428 11076 11480 11082
rect 10692 11018 10744 11024
rect 11428 11018 11480 11024
rect 10508 10124 10560 10130
rect 10508 10066 10560 10072
rect 10416 9920 10468 9926
rect 10416 9862 10468 9868
rect 10428 9042 10456 9862
rect 10416 9036 10468 9042
rect 10416 8978 10468 8984
rect 10324 7540 10376 7546
rect 10324 7482 10376 7488
rect 10704 7206 10732 11018
rect 10876 11008 10928 11014
rect 10876 10950 10928 10956
rect 10888 10810 10916 10950
rect 10876 10804 10928 10810
rect 10876 10746 10928 10752
rect 10784 10056 10836 10062
rect 10784 9998 10836 10004
rect 10796 9722 10824 9998
rect 11888 9920 11940 9926
rect 11888 9862 11940 9868
rect 10784 9716 10836 9722
rect 10784 9658 10836 9664
rect 11900 9178 11928 9862
rect 11992 9654 12020 16118
rect 12256 16108 12308 16114
rect 12256 16050 12308 16056
rect 13728 16108 13780 16114
rect 13728 16050 13780 16056
rect 15476 16108 15528 16114
rect 15476 16050 15528 16056
rect 15660 16108 15712 16114
rect 15660 16050 15712 16056
rect 12268 15570 12296 16050
rect 13740 15910 13768 16050
rect 14096 16040 14148 16046
rect 14280 16040 14332 16046
rect 14148 16000 14280 16028
rect 14096 15982 14148 15988
rect 14280 15982 14332 15988
rect 14740 16040 14792 16046
rect 14740 15982 14792 15988
rect 14832 16040 14884 16046
rect 14832 15982 14884 15988
rect 15384 16040 15436 16046
rect 15384 15982 15436 15988
rect 12808 15904 12860 15910
rect 12808 15846 12860 15852
rect 13728 15904 13780 15910
rect 13728 15846 13780 15852
rect 14096 15904 14148 15910
rect 14096 15846 14148 15852
rect 12440 15632 12492 15638
rect 12440 15574 12492 15580
rect 12256 15564 12308 15570
rect 12256 15506 12308 15512
rect 12268 15366 12296 15506
rect 12256 15360 12308 15366
rect 12256 15302 12308 15308
rect 12268 15026 12296 15302
rect 12452 15026 12480 15574
rect 12532 15360 12584 15366
rect 12532 15302 12584 15308
rect 12544 15094 12572 15302
rect 12820 15094 12848 15846
rect 13740 15722 13768 15846
rect 13740 15694 13860 15722
rect 13728 15632 13780 15638
rect 13728 15574 13780 15580
rect 13740 15502 13768 15574
rect 12900 15496 12952 15502
rect 12900 15438 12952 15444
rect 13728 15496 13780 15502
rect 13728 15438 13780 15444
rect 12532 15088 12584 15094
rect 12532 15030 12584 15036
rect 12808 15088 12860 15094
rect 12808 15030 12860 15036
rect 12256 15020 12308 15026
rect 12440 15020 12492 15026
rect 12256 14962 12308 14968
rect 12360 14980 12440 15008
rect 12072 14884 12124 14890
rect 12072 14826 12124 14832
rect 12084 14550 12112 14826
rect 12072 14544 12124 14550
rect 12072 14486 12124 14492
rect 12084 14006 12112 14486
rect 12268 14385 12296 14962
rect 12360 14618 12388 14980
rect 12912 15008 12940 15438
rect 13832 15434 13860 15694
rect 14108 15638 14136 15846
rect 14096 15632 14148 15638
rect 14096 15574 14148 15580
rect 14096 15496 14148 15502
rect 14292 15450 14320 15982
rect 14148 15444 14320 15450
rect 14096 15438 14320 15444
rect 13360 15428 13412 15434
rect 13360 15370 13412 15376
rect 13820 15428 13872 15434
rect 13820 15370 13872 15376
rect 14108 15422 14320 15438
rect 13176 15360 13228 15366
rect 13176 15302 13228 15308
rect 12992 15020 13044 15026
rect 12912 14980 12992 15008
rect 12440 14962 12492 14968
rect 12992 14962 13044 14968
rect 12440 14816 12492 14822
rect 12440 14758 12492 14764
rect 12624 14816 12676 14822
rect 12624 14758 12676 14764
rect 12348 14612 12400 14618
rect 12348 14554 12400 14560
rect 12452 14482 12480 14758
rect 12440 14476 12492 14482
rect 12440 14418 12492 14424
rect 12254 14376 12310 14385
rect 12254 14311 12256 14320
rect 12308 14311 12310 14320
rect 12256 14282 12308 14288
rect 12636 14278 12664 14758
rect 13004 14414 13032 14962
rect 13188 14822 13216 15302
rect 13372 15026 13400 15370
rect 13452 15360 13504 15366
rect 13452 15302 13504 15308
rect 13360 15020 13412 15026
rect 13360 14962 13412 14968
rect 13176 14816 13228 14822
rect 13176 14758 13228 14764
rect 13268 14816 13320 14822
rect 13268 14758 13320 14764
rect 13188 14414 13216 14758
rect 12992 14408 13044 14414
rect 13084 14408 13136 14414
rect 12992 14350 13044 14356
rect 13082 14376 13084 14385
rect 13176 14408 13228 14414
rect 13136 14376 13138 14385
rect 12624 14272 12676 14278
rect 12624 14214 12676 14220
rect 12716 14272 12768 14278
rect 12716 14214 12768 14220
rect 12808 14272 12860 14278
rect 12808 14214 12860 14220
rect 12728 14006 12756 14214
rect 12072 14000 12124 14006
rect 12072 13942 12124 13948
rect 12716 14000 12768 14006
rect 12716 13942 12768 13948
rect 12072 13864 12124 13870
rect 12072 13806 12124 13812
rect 12084 12850 12112 13806
rect 12820 13802 12848 14214
rect 13004 14074 13032 14350
rect 13176 14350 13228 14356
rect 13082 14311 13138 14320
rect 12992 14068 13044 14074
rect 12992 14010 13044 14016
rect 12808 13796 12860 13802
rect 12808 13738 12860 13744
rect 13096 13258 13124 14311
rect 13280 13870 13308 14758
rect 13464 14414 13492 15302
rect 13820 14612 13872 14618
rect 13820 14554 13872 14560
rect 13360 14408 13412 14414
rect 13360 14350 13412 14356
rect 13452 14408 13504 14414
rect 13452 14350 13504 14356
rect 13372 13920 13400 14350
rect 13728 14340 13780 14346
rect 13648 14300 13728 14328
rect 13648 13938 13676 14300
rect 13728 14282 13780 14288
rect 13636 13932 13688 13938
rect 13372 13892 13636 13920
rect 13636 13874 13688 13880
rect 13268 13864 13320 13870
rect 13268 13806 13320 13812
rect 13832 13802 13860 14554
rect 14108 14550 14136 15422
rect 14752 15366 14780 15982
rect 14844 15706 14872 15982
rect 14832 15700 14884 15706
rect 14832 15642 14884 15648
rect 15396 15638 15424 15982
rect 15384 15632 15436 15638
rect 15384 15574 15436 15580
rect 14740 15360 14792 15366
rect 14740 15302 14792 15308
rect 14924 15020 14976 15026
rect 14924 14962 14976 14968
rect 15292 15020 15344 15026
rect 15396 15008 15424 15574
rect 15488 15502 15516 16050
rect 15568 15904 15620 15910
rect 15568 15846 15620 15852
rect 15580 15502 15608 15846
rect 15476 15496 15528 15502
rect 15476 15438 15528 15444
rect 15568 15496 15620 15502
rect 15568 15438 15620 15444
rect 15672 15162 15700 16050
rect 16028 15972 16080 15978
rect 16028 15914 16080 15920
rect 15752 15632 15804 15638
rect 15752 15574 15804 15580
rect 15660 15156 15712 15162
rect 15660 15098 15712 15104
rect 15764 15026 15792 15574
rect 15844 15496 15896 15502
rect 15844 15438 15896 15444
rect 15344 14980 15424 15008
rect 15476 15020 15528 15026
rect 15292 14962 15344 14968
rect 15476 14962 15528 14968
rect 15752 15020 15804 15026
rect 15752 14962 15804 14968
rect 14936 14618 14964 14962
rect 14924 14612 14976 14618
rect 14924 14554 14976 14560
rect 14096 14544 14148 14550
rect 14096 14486 14148 14492
rect 14188 14476 14240 14482
rect 14188 14418 14240 14424
rect 14096 14340 14148 14346
rect 14200 14328 14228 14418
rect 14148 14300 14228 14328
rect 15292 14340 15344 14346
rect 14096 14282 14148 14288
rect 15292 14282 15344 14288
rect 13360 13796 13412 13802
rect 13360 13738 13412 13744
rect 13820 13796 13872 13802
rect 13820 13738 13872 13744
rect 13084 13252 13136 13258
rect 13084 13194 13136 13200
rect 12072 12844 12124 12850
rect 12072 12786 12124 12792
rect 12164 12640 12216 12646
rect 12164 12582 12216 12588
rect 12176 12238 12204 12582
rect 12348 12368 12400 12374
rect 12348 12310 12400 12316
rect 12256 12300 12308 12306
rect 12256 12242 12308 12248
rect 12164 12232 12216 12238
rect 12164 12174 12216 12180
rect 12072 12164 12124 12170
rect 12072 12106 12124 12112
rect 12084 11830 12112 12106
rect 12268 11898 12296 12242
rect 12256 11892 12308 11898
rect 12256 11834 12308 11840
rect 12072 11824 12124 11830
rect 12072 11766 12124 11772
rect 12084 11218 12112 11766
rect 12360 11762 12388 12310
rect 13372 12238 13400 13738
rect 13832 12850 13860 13738
rect 14108 13530 14136 14282
rect 14280 14272 14332 14278
rect 14280 14214 14332 14220
rect 14292 14006 14320 14214
rect 14280 14000 14332 14006
rect 14280 13942 14332 13948
rect 14096 13524 14148 13530
rect 14096 13466 14148 13472
rect 15304 13326 15332 14282
rect 15488 14074 15516 14962
rect 15856 14618 15884 15438
rect 16040 15026 16068 15914
rect 16580 15564 16632 15570
rect 16580 15506 16632 15512
rect 16304 15496 16356 15502
rect 16304 15438 16356 15444
rect 16212 15360 16264 15366
rect 16212 15302 16264 15308
rect 16224 15026 16252 15302
rect 16316 15162 16344 15438
rect 16304 15156 16356 15162
rect 16304 15098 16356 15104
rect 16028 15020 16080 15026
rect 16028 14962 16080 14968
rect 16212 15020 16264 15026
rect 16212 14962 16264 14968
rect 15844 14612 15896 14618
rect 15844 14554 15896 14560
rect 15752 14272 15804 14278
rect 15752 14214 15804 14220
rect 15476 14068 15528 14074
rect 15476 14010 15528 14016
rect 15764 13326 15792 14214
rect 16224 13326 16252 14962
rect 16592 14958 16620 15506
rect 16776 15094 16804 20878
rect 17052 20602 17080 21490
rect 17040 20596 17092 20602
rect 17040 20538 17092 20544
rect 17144 19922 17172 21490
rect 17512 21486 17540 21830
rect 17788 21554 17816 21898
rect 17972 21690 18000 21966
rect 17960 21684 18012 21690
rect 17960 21626 18012 21632
rect 18052 21616 18104 21622
rect 18052 21558 18104 21564
rect 17776 21548 17828 21554
rect 17776 21490 17828 21496
rect 17500 21480 17552 21486
rect 17500 21422 17552 21428
rect 17500 20868 17552 20874
rect 17500 20810 17552 20816
rect 17512 20466 17540 20810
rect 17500 20460 17552 20466
rect 17500 20402 17552 20408
rect 17132 19916 17184 19922
rect 17132 19858 17184 19864
rect 17408 18828 17460 18834
rect 17408 18770 17460 18776
rect 17040 18692 17092 18698
rect 17040 18634 17092 18640
rect 16856 18624 16908 18630
rect 16856 18566 16908 18572
rect 16868 17882 16896 18566
rect 17052 18426 17080 18634
rect 17040 18420 17092 18426
rect 17040 18362 17092 18368
rect 17224 18080 17276 18086
rect 17224 18022 17276 18028
rect 16856 17876 16908 17882
rect 16856 17818 16908 17824
rect 17040 17808 17092 17814
rect 17040 17750 17092 17756
rect 17052 17270 17080 17750
rect 17236 17678 17264 18022
rect 17420 17814 17448 18770
rect 17788 18766 17816 21490
rect 17960 21072 18012 21078
rect 17960 21014 18012 21020
rect 17868 20868 17920 20874
rect 17868 20810 17920 20816
rect 17880 19514 17908 20810
rect 17972 20466 18000 21014
rect 17960 20460 18012 20466
rect 17960 20402 18012 20408
rect 17972 19514 18000 20402
rect 17868 19508 17920 19514
rect 17868 19450 17920 19456
rect 17960 19508 18012 19514
rect 17960 19450 18012 19456
rect 17880 19394 17908 19450
rect 17880 19366 17954 19394
rect 17926 19360 17954 19366
rect 17926 19332 18000 19360
rect 17776 18760 17828 18766
rect 17776 18702 17828 18708
rect 17684 18080 17736 18086
rect 17684 18022 17736 18028
rect 17408 17808 17460 17814
rect 17408 17750 17460 17756
rect 17224 17672 17276 17678
rect 17224 17614 17276 17620
rect 17696 17338 17724 18022
rect 17972 17678 18000 19332
rect 18064 18698 18092 21558
rect 18248 21146 18276 22102
rect 18340 21554 18368 23462
rect 18420 22024 18472 22030
rect 18420 21966 18472 21972
rect 18432 21690 18460 21966
rect 18524 21690 18552 23598
rect 18420 21684 18472 21690
rect 18420 21626 18472 21632
rect 18512 21684 18564 21690
rect 18512 21626 18564 21632
rect 18328 21548 18380 21554
rect 18328 21490 18380 21496
rect 18236 21140 18288 21146
rect 18236 21082 18288 21088
rect 18144 20392 18196 20398
rect 18144 20334 18196 20340
rect 18616 20346 18644 24006
rect 18892 23662 18920 24346
rect 18972 24200 19024 24206
rect 18972 24142 19024 24148
rect 18880 23656 18932 23662
rect 18880 23598 18932 23604
rect 18892 23186 18920 23598
rect 18984 23594 19012 24142
rect 19076 23730 19104 24398
rect 19156 24336 19208 24342
rect 19156 24278 19208 24284
rect 19168 23798 19196 24278
rect 19260 24274 19288 24398
rect 19248 24268 19300 24274
rect 19248 24210 19300 24216
rect 19246 24168 19302 24177
rect 19246 24103 19302 24112
rect 19260 23866 19288 24103
rect 19248 23860 19300 23866
rect 19248 23802 19300 23808
rect 19156 23792 19208 23798
rect 19156 23734 19208 23740
rect 19064 23724 19116 23730
rect 19064 23666 19116 23672
rect 18972 23588 19024 23594
rect 18972 23530 19024 23536
rect 19352 23526 19380 24686
rect 19432 24608 19484 24614
rect 19432 24550 19484 24556
rect 19444 24290 19472 24550
rect 19812 24410 19840 24686
rect 19800 24404 19852 24410
rect 19800 24346 19852 24352
rect 19444 24262 19748 24290
rect 19904 24274 19932 24890
rect 20812 24676 20864 24682
rect 20812 24618 20864 24624
rect 20536 24608 20588 24614
rect 20536 24550 20588 24556
rect 19720 24206 19748 24262
rect 19892 24268 19944 24274
rect 19892 24210 19944 24216
rect 19708 24200 19760 24206
rect 19708 24142 19760 24148
rect 20076 24200 20128 24206
rect 20076 24142 20128 24148
rect 19616 24064 19668 24070
rect 19616 24006 19668 24012
rect 19892 24064 19944 24070
rect 19892 24006 19944 24012
rect 19628 23798 19656 24006
rect 19904 23798 19932 24006
rect 19616 23792 19668 23798
rect 19616 23734 19668 23740
rect 19892 23792 19944 23798
rect 19892 23734 19944 23740
rect 19708 23724 19760 23730
rect 19708 23666 19760 23672
rect 19340 23520 19392 23526
rect 19340 23462 19392 23468
rect 18880 23180 18932 23186
rect 18880 23122 18932 23128
rect 18892 21554 18920 23122
rect 19720 22094 19748 23666
rect 19800 23656 19852 23662
rect 19800 23598 19852 23604
rect 19892 23656 19944 23662
rect 19892 23598 19944 23604
rect 19812 23526 19840 23598
rect 19800 23520 19852 23526
rect 19800 23462 19852 23468
rect 19798 22264 19854 22273
rect 19798 22199 19854 22208
rect 19812 22166 19840 22199
rect 19800 22160 19852 22166
rect 19800 22102 19852 22108
rect 19536 22066 19748 22094
rect 19064 21888 19116 21894
rect 19064 21830 19116 21836
rect 19248 21888 19300 21894
rect 19248 21830 19300 21836
rect 19432 21888 19484 21894
rect 19432 21830 19484 21836
rect 18880 21548 18932 21554
rect 18880 21490 18932 21496
rect 19076 21010 19104 21830
rect 19260 21622 19288 21830
rect 19248 21616 19300 21622
rect 19248 21558 19300 21564
rect 19248 21344 19300 21350
rect 19248 21286 19300 21292
rect 19064 21004 19116 21010
rect 19064 20946 19116 20952
rect 19076 20874 19104 20946
rect 19260 20942 19288 21286
rect 19248 20936 19300 20942
rect 19248 20878 19300 20884
rect 19064 20868 19116 20874
rect 19064 20810 19116 20816
rect 19260 20806 19288 20878
rect 19444 20806 19472 21830
rect 18696 20800 18748 20806
rect 18696 20742 18748 20748
rect 19248 20800 19300 20806
rect 19248 20742 19300 20748
rect 19432 20800 19484 20806
rect 19432 20742 19484 20748
rect 18708 20534 18736 20742
rect 18696 20528 18748 20534
rect 18696 20470 18748 20476
rect 18788 20460 18840 20466
rect 18788 20402 18840 20408
rect 18052 18692 18104 18698
rect 18052 18634 18104 18640
rect 17960 17672 18012 17678
rect 17960 17614 18012 17620
rect 18064 17338 18092 18634
rect 18156 18358 18184 20334
rect 18616 20318 18736 20346
rect 18420 20256 18472 20262
rect 18420 20198 18472 20204
rect 18432 19922 18460 20198
rect 18420 19916 18472 19922
rect 18420 19858 18472 19864
rect 18236 19508 18288 19514
rect 18236 19450 18288 19456
rect 18248 18766 18276 19450
rect 18708 18766 18736 20318
rect 18800 20058 18828 20402
rect 18788 20052 18840 20058
rect 18788 19994 18840 20000
rect 19444 19786 19472 20742
rect 19432 19780 19484 19786
rect 19432 19722 19484 19728
rect 18800 19094 19104 19122
rect 18800 18970 18828 19094
rect 19076 18970 19104 19094
rect 18788 18964 18840 18970
rect 18788 18906 18840 18912
rect 18880 18964 18932 18970
rect 19064 18964 19116 18970
rect 18932 18924 19012 18952
rect 18880 18906 18932 18912
rect 18236 18760 18288 18766
rect 18236 18702 18288 18708
rect 18696 18760 18748 18766
rect 18696 18702 18748 18708
rect 18880 18624 18932 18630
rect 18880 18566 18932 18572
rect 18144 18352 18196 18358
rect 18144 18294 18196 18300
rect 18892 17882 18920 18566
rect 18984 17882 19012 18924
rect 19064 18906 19116 18912
rect 19156 18692 19208 18698
rect 19156 18634 19208 18640
rect 19064 18148 19116 18154
rect 19064 18090 19116 18096
rect 18880 17876 18932 17882
rect 18880 17818 18932 17824
rect 18972 17876 19024 17882
rect 18972 17818 19024 17824
rect 18420 17740 18472 17746
rect 18420 17682 18472 17688
rect 18328 17536 18380 17542
rect 18328 17478 18380 17484
rect 17684 17332 17736 17338
rect 17684 17274 17736 17280
rect 18052 17332 18104 17338
rect 18052 17274 18104 17280
rect 18340 17270 18368 17478
rect 17040 17264 17092 17270
rect 17040 17206 17092 17212
rect 17500 17264 17552 17270
rect 17500 17206 17552 17212
rect 18328 17264 18380 17270
rect 18328 17206 18380 17212
rect 17512 17134 17540 17206
rect 17500 17128 17552 17134
rect 17500 17070 17552 17076
rect 17512 15434 17540 17070
rect 18432 16114 18460 17682
rect 19076 17678 19104 18090
rect 19168 18086 19196 18634
rect 19156 18080 19208 18086
rect 19156 18022 19208 18028
rect 19064 17672 19116 17678
rect 19064 17614 19116 17620
rect 19168 17338 19196 18022
rect 19156 17332 19208 17338
rect 19156 17274 19208 17280
rect 19444 17202 19472 19722
rect 19536 19514 19564 22066
rect 19812 20942 19840 22102
rect 19904 21894 19932 23598
rect 19984 22160 20036 22166
rect 19984 22102 20036 22108
rect 19996 21894 20024 22102
rect 19892 21888 19944 21894
rect 19892 21830 19944 21836
rect 19984 21888 20036 21894
rect 19984 21830 20036 21836
rect 19996 21706 20024 21830
rect 19904 21678 20024 21706
rect 19904 21486 19932 21678
rect 20088 21570 20116 24142
rect 20168 24064 20220 24070
rect 20168 24006 20220 24012
rect 20180 23798 20208 24006
rect 20168 23792 20220 23798
rect 20168 23734 20220 23740
rect 20548 23474 20576 24550
rect 20628 24268 20680 24274
rect 20628 24210 20680 24216
rect 20640 23662 20668 24210
rect 20824 23866 20852 24618
rect 21008 24342 21036 25094
rect 21100 24886 21128 25162
rect 21088 24880 21140 24886
rect 21088 24822 21140 24828
rect 21548 24880 21600 24886
rect 21548 24822 21600 24828
rect 21730 24848 21786 24857
rect 21364 24812 21416 24818
rect 21364 24754 21416 24760
rect 21086 24712 21142 24721
rect 21086 24647 21142 24656
rect 21100 24410 21128 24647
rect 21180 24608 21232 24614
rect 21180 24550 21232 24556
rect 21088 24404 21140 24410
rect 21088 24346 21140 24352
rect 20996 24336 21048 24342
rect 20996 24278 21048 24284
rect 20904 24200 20956 24206
rect 20904 24142 20956 24148
rect 20812 23860 20864 23866
rect 20812 23802 20864 23808
rect 20916 23662 20944 24142
rect 21088 24064 21140 24070
rect 21088 24006 21140 24012
rect 21100 23866 21128 24006
rect 21088 23860 21140 23866
rect 21088 23802 21140 23808
rect 20996 23792 21048 23798
rect 20996 23734 21048 23740
rect 20628 23656 20680 23662
rect 20628 23598 20680 23604
rect 20904 23656 20956 23662
rect 20904 23598 20956 23604
rect 20812 23520 20864 23526
rect 20548 23446 20760 23474
rect 21008 23497 21036 23734
rect 21100 23594 21128 23802
rect 21192 23730 21220 24550
rect 21272 24200 21324 24206
rect 21270 24168 21272 24177
rect 21324 24168 21326 24177
rect 21270 24103 21326 24112
rect 21180 23724 21232 23730
rect 21180 23666 21232 23672
rect 21088 23588 21140 23594
rect 21088 23530 21140 23536
rect 20812 23462 20864 23468
rect 20994 23488 21050 23497
rect 20444 22092 20496 22098
rect 20444 22034 20496 22040
rect 20168 21956 20220 21962
rect 20168 21898 20220 21904
rect 19996 21542 20116 21570
rect 19892 21480 19944 21486
rect 19892 21422 19944 21428
rect 19708 20936 19760 20942
rect 19708 20878 19760 20884
rect 19800 20936 19852 20942
rect 19800 20878 19852 20884
rect 19720 20602 19748 20878
rect 19708 20596 19760 20602
rect 19708 20538 19760 20544
rect 19616 19848 19668 19854
rect 19616 19790 19668 19796
rect 19524 19508 19576 19514
rect 19524 19450 19576 19456
rect 19524 18624 19576 18630
rect 19524 18566 19576 18572
rect 19536 17610 19564 18566
rect 19628 18426 19656 19790
rect 19720 19360 19748 20538
rect 19812 20466 19840 20878
rect 19996 20482 20024 21542
rect 20076 21480 20128 21486
rect 20076 21422 20128 21428
rect 20088 20602 20116 21422
rect 20180 20942 20208 21898
rect 20168 20936 20220 20942
rect 20168 20878 20220 20884
rect 20076 20596 20128 20602
rect 20076 20538 20128 20544
rect 19800 20460 19852 20466
rect 19996 20454 20116 20482
rect 19800 20402 19852 20408
rect 19984 20256 20036 20262
rect 19984 20198 20036 20204
rect 19996 20058 20024 20198
rect 19984 20052 20036 20058
rect 19984 19994 20036 20000
rect 19892 19712 19944 19718
rect 19892 19654 19944 19660
rect 19904 19378 19932 19654
rect 19892 19372 19944 19378
rect 19720 19332 19840 19360
rect 19708 19168 19760 19174
rect 19708 19110 19760 19116
rect 19720 18970 19748 19110
rect 19708 18964 19760 18970
rect 19708 18906 19760 18912
rect 19616 18420 19668 18426
rect 19616 18362 19668 18368
rect 19524 17604 19576 17610
rect 19524 17546 19576 17552
rect 19432 17196 19484 17202
rect 19432 17138 19484 17144
rect 18420 16108 18472 16114
rect 18420 16050 18472 16056
rect 17776 15904 17828 15910
rect 17776 15846 17828 15852
rect 17500 15428 17552 15434
rect 17500 15370 17552 15376
rect 17224 15360 17276 15366
rect 17224 15302 17276 15308
rect 16764 15088 16816 15094
rect 16764 15030 16816 15036
rect 17236 15026 17264 15302
rect 17224 15020 17276 15026
rect 17224 14962 17276 14968
rect 16580 14952 16632 14958
rect 16580 14894 16632 14900
rect 16304 13524 16356 13530
rect 16304 13466 16356 13472
rect 15292 13320 15344 13326
rect 15292 13262 15344 13268
rect 15752 13320 15804 13326
rect 15752 13262 15804 13268
rect 16028 13320 16080 13326
rect 16028 13262 16080 13268
rect 16212 13320 16264 13326
rect 16212 13262 16264 13268
rect 15016 13184 15068 13190
rect 15016 13126 15068 13132
rect 15028 12850 15056 13126
rect 13820 12844 13872 12850
rect 13820 12786 13872 12792
rect 15016 12844 15068 12850
rect 15016 12786 15068 12792
rect 12808 12232 12860 12238
rect 12808 12174 12860 12180
rect 13360 12232 13412 12238
rect 13360 12174 13412 12180
rect 12716 12096 12768 12102
rect 12716 12038 12768 12044
rect 12348 11756 12400 11762
rect 12348 11698 12400 11704
rect 12728 11694 12756 12038
rect 12820 11830 12848 12174
rect 13176 12164 13228 12170
rect 13176 12106 13228 12112
rect 12808 11824 12860 11830
rect 12808 11766 12860 11772
rect 13188 11762 13216 12106
rect 13372 11762 13400 12174
rect 13176 11756 13228 11762
rect 13176 11698 13228 11704
rect 13360 11756 13412 11762
rect 13360 11698 13412 11704
rect 12716 11688 12768 11694
rect 12716 11630 12768 11636
rect 13452 11620 13504 11626
rect 13452 11562 13504 11568
rect 12072 11212 12124 11218
rect 12072 11154 12124 11160
rect 13360 11144 13412 11150
rect 13360 11086 13412 11092
rect 12900 11008 12952 11014
rect 12900 10950 12952 10956
rect 13268 11008 13320 11014
rect 13268 10950 13320 10956
rect 12912 10810 12940 10950
rect 12900 10804 12952 10810
rect 12900 10746 12952 10752
rect 13280 10674 13308 10950
rect 13372 10674 13400 11086
rect 13464 10674 13492 11562
rect 13832 11150 13860 12786
rect 14648 12776 14700 12782
rect 14648 12718 14700 12724
rect 14660 12434 14688 12718
rect 15304 12434 15332 13262
rect 16040 12434 16068 13262
rect 16316 12918 16344 13466
rect 16304 12912 16356 12918
rect 16304 12854 16356 12860
rect 14660 12406 14872 12434
rect 15304 12406 15424 12434
rect 14844 12238 14872 12406
rect 14832 12232 14884 12238
rect 14832 12174 14884 12180
rect 13912 12096 13964 12102
rect 13912 12038 13964 12044
rect 13924 11762 13952 12038
rect 13912 11756 13964 11762
rect 13912 11698 13964 11704
rect 14844 11218 14872 12174
rect 14832 11212 14884 11218
rect 14832 11154 14884 11160
rect 13636 11144 13688 11150
rect 13820 11144 13872 11150
rect 13688 11104 13768 11132
rect 13636 11086 13688 11092
rect 13740 10674 13768 11104
rect 13820 11086 13872 11092
rect 13832 10810 13860 11086
rect 13912 11008 13964 11014
rect 13912 10950 13964 10956
rect 13820 10804 13872 10810
rect 13820 10746 13872 10752
rect 13832 10674 13860 10746
rect 13268 10668 13320 10674
rect 13268 10610 13320 10616
rect 13360 10668 13412 10674
rect 13360 10610 13412 10616
rect 13452 10668 13504 10674
rect 13452 10610 13504 10616
rect 13728 10668 13780 10674
rect 13728 10610 13780 10616
rect 13820 10668 13872 10674
rect 13820 10610 13872 10616
rect 13372 10062 13400 10610
rect 13464 10130 13492 10610
rect 13740 10538 13768 10610
rect 13728 10532 13780 10538
rect 13728 10474 13780 10480
rect 13924 10470 13952 10950
rect 13544 10464 13596 10470
rect 13544 10406 13596 10412
rect 13912 10464 13964 10470
rect 13912 10406 13964 10412
rect 14004 10464 14056 10470
rect 14004 10406 14056 10412
rect 14372 10464 14424 10470
rect 14372 10406 14424 10412
rect 15200 10464 15252 10470
rect 15200 10406 15252 10412
rect 13452 10124 13504 10130
rect 13452 10066 13504 10072
rect 13556 10062 13584 10406
rect 14016 10130 14044 10406
rect 14004 10124 14056 10130
rect 14004 10066 14056 10072
rect 14384 10062 14412 10406
rect 13360 10056 13412 10062
rect 13360 9998 13412 10004
rect 13544 10056 13596 10062
rect 13544 9998 13596 10004
rect 13912 10056 13964 10062
rect 13912 9998 13964 10004
rect 14188 10056 14240 10062
rect 14188 9998 14240 10004
rect 14372 10056 14424 10062
rect 14372 9998 14424 10004
rect 11980 9648 12032 9654
rect 11980 9590 12032 9596
rect 13636 9648 13688 9654
rect 13636 9590 13688 9596
rect 12164 9580 12216 9586
rect 12164 9522 12216 9528
rect 12176 9450 12204 9522
rect 12164 9444 12216 9450
rect 12164 9386 12216 9392
rect 10968 9172 11020 9178
rect 10968 9114 11020 9120
rect 11888 9172 11940 9178
rect 11888 9114 11940 9120
rect 10784 9036 10836 9042
rect 10784 8978 10836 8984
rect 10796 8498 10824 8978
rect 10980 8906 11008 9114
rect 11796 9036 11848 9042
rect 11796 8978 11848 8984
rect 10968 8900 11020 8906
rect 10968 8842 11020 8848
rect 10784 8492 10836 8498
rect 10784 8434 10836 8440
rect 11704 7404 11756 7410
rect 11704 7346 11756 7352
rect 10324 7200 10376 7206
rect 10324 7142 10376 7148
rect 10692 7200 10744 7206
rect 10692 7142 10744 7148
rect 10192 6684 10272 6712
rect 10140 6666 10192 6672
rect 10152 6458 10180 6666
rect 10140 6452 10192 6458
rect 10140 6394 10192 6400
rect 9588 6326 9640 6332
rect 9862 6352 9918 6361
rect 9036 6316 9088 6322
rect 10152 6322 10180 6394
rect 10336 6322 10364 7142
rect 11716 7002 11744 7346
rect 11060 6996 11112 7002
rect 11060 6938 11112 6944
rect 11612 6996 11664 7002
rect 11612 6938 11664 6944
rect 11704 6996 11756 7002
rect 11704 6938 11756 6944
rect 10876 6452 10928 6458
rect 10876 6394 10928 6400
rect 9862 6287 9918 6296
rect 10140 6316 10192 6322
rect 9036 6258 9088 6264
rect 9048 5642 9076 6258
rect 9036 5636 9088 5642
rect 9036 5578 9088 5584
rect 9048 5302 9076 5578
rect 9876 5302 9904 6287
rect 10140 6258 10192 6264
rect 10324 6316 10376 6322
rect 10324 6258 10376 6264
rect 10336 5370 10364 6258
rect 10888 5914 10916 6394
rect 10416 5908 10468 5914
rect 10416 5850 10468 5856
rect 10876 5908 10928 5914
rect 10876 5850 10928 5856
rect 10428 5642 10456 5850
rect 10508 5840 10560 5846
rect 10508 5782 10560 5788
rect 10520 5642 10548 5782
rect 10888 5710 10916 5850
rect 11072 5846 11100 6938
rect 11624 6866 11652 6938
rect 11612 6860 11664 6866
rect 11612 6802 11664 6808
rect 11624 6730 11652 6802
rect 11808 6730 11836 8978
rect 12176 8974 12204 9386
rect 12900 9376 12952 9382
rect 12900 9318 12952 9324
rect 12348 9172 12400 9178
rect 12348 9114 12400 9120
rect 12360 8974 12388 9114
rect 12164 8968 12216 8974
rect 12164 8910 12216 8916
rect 12348 8968 12400 8974
rect 12348 8910 12400 8916
rect 12532 8968 12584 8974
rect 12532 8910 12584 8916
rect 11888 8832 11940 8838
rect 11888 8774 11940 8780
rect 11900 6769 11928 8774
rect 12176 8430 12204 8910
rect 12544 8498 12572 8910
rect 12912 8906 12940 9318
rect 13648 9178 13676 9590
rect 13924 9518 13952 9998
rect 14200 9722 14228 9998
rect 14188 9716 14240 9722
rect 14188 9658 14240 9664
rect 15212 9586 15240 10406
rect 15292 9920 15344 9926
rect 15292 9862 15344 9868
rect 15108 9580 15160 9586
rect 15108 9522 15160 9528
rect 15200 9580 15252 9586
rect 15200 9522 15252 9528
rect 13912 9512 13964 9518
rect 13912 9454 13964 9460
rect 14280 9512 14332 9518
rect 14280 9454 14332 9460
rect 15120 9466 15148 9522
rect 15304 9466 15332 9862
rect 13636 9172 13688 9178
rect 13636 9114 13688 9120
rect 14292 9042 14320 9454
rect 15120 9438 15332 9466
rect 15396 9178 15424 12406
rect 15856 12406 16068 12434
rect 15568 11348 15620 11354
rect 15568 11290 15620 11296
rect 15580 11150 15608 11290
rect 15568 11144 15620 11150
rect 15568 11086 15620 11092
rect 15752 10056 15804 10062
rect 15752 9998 15804 10004
rect 15764 9518 15792 9998
rect 15856 9994 15884 12406
rect 16396 12164 16448 12170
rect 16396 12106 16448 12112
rect 15936 11212 15988 11218
rect 15936 11154 15988 11160
rect 15948 10674 15976 11154
rect 16408 11082 16436 12106
rect 16592 11218 16620 14894
rect 17040 13932 17092 13938
rect 17040 13874 17092 13880
rect 16764 13320 16816 13326
rect 16764 13262 16816 13268
rect 16776 12986 16804 13262
rect 17052 13190 17080 13874
rect 17236 13258 17264 14962
rect 17316 14952 17368 14958
rect 17316 14894 17368 14900
rect 17328 14618 17356 14894
rect 17316 14612 17368 14618
rect 17316 14554 17368 14560
rect 17788 14482 17816 15846
rect 19812 15706 19840 19332
rect 19892 19314 19944 19320
rect 20088 19122 20116 20454
rect 20180 19446 20208 20878
rect 20456 19854 20484 22034
rect 20732 21554 20760 23446
rect 20824 23322 20852 23462
rect 20994 23423 21050 23432
rect 20812 23316 20864 23322
rect 20812 23258 20864 23264
rect 21008 22710 21036 23423
rect 20996 22704 21048 22710
rect 20996 22646 21048 22652
rect 21100 22642 21128 23530
rect 21284 23526 21312 24103
rect 21376 23798 21404 24754
rect 21560 24206 21588 24822
rect 21730 24783 21786 24792
rect 22376 24812 22428 24818
rect 21548 24200 21600 24206
rect 21548 24142 21600 24148
rect 21364 23792 21416 23798
rect 21364 23734 21416 23740
rect 21272 23520 21324 23526
rect 21272 23462 21324 23468
rect 21088 22636 21140 22642
rect 21088 22578 21140 22584
rect 21560 22094 21588 24142
rect 21744 22642 21772 24783
rect 22376 24754 22428 24760
rect 22652 24812 22704 24818
rect 22652 24754 22704 24760
rect 22388 24410 22416 24754
rect 22376 24404 22428 24410
rect 22376 24346 22428 24352
rect 22388 23866 22416 24346
rect 22664 23866 22692 24754
rect 23020 24608 23072 24614
rect 23020 24550 23072 24556
rect 22928 24268 22980 24274
rect 22928 24210 22980 24216
rect 22744 24064 22796 24070
rect 22744 24006 22796 24012
rect 22376 23860 22428 23866
rect 22376 23802 22428 23808
rect 22652 23860 22704 23866
rect 22652 23802 22704 23808
rect 22756 23746 22784 24006
rect 22284 23724 22336 23730
rect 22284 23666 22336 23672
rect 22664 23718 22784 23746
rect 21732 22636 21784 22642
rect 21732 22578 21784 22584
rect 21468 22066 21588 22094
rect 20996 21888 21048 21894
rect 20996 21830 21048 21836
rect 20720 21548 20772 21554
rect 20720 21490 20772 21496
rect 21008 20466 21036 21830
rect 21180 21344 21232 21350
rect 21180 21286 21232 21292
rect 20996 20460 21048 20466
rect 20996 20402 21048 20408
rect 21192 20398 21220 21286
rect 20720 20392 20772 20398
rect 20720 20334 20772 20340
rect 21180 20392 21232 20398
rect 21180 20334 21232 20340
rect 20444 19848 20496 19854
rect 20444 19790 20496 19796
rect 20168 19440 20220 19446
rect 20168 19382 20220 19388
rect 19904 19094 20116 19122
rect 19904 16046 19932 19094
rect 20180 18970 20208 19382
rect 20628 19372 20680 19378
rect 20628 19314 20680 19320
rect 20168 18964 20220 18970
rect 20168 18906 20220 18912
rect 20180 18766 20208 18906
rect 20640 18834 20668 19314
rect 20628 18828 20680 18834
rect 20628 18770 20680 18776
rect 20168 18760 20220 18766
rect 20168 18702 20220 18708
rect 19984 18692 20036 18698
rect 19984 18634 20036 18640
rect 19996 18426 20024 18634
rect 19984 18420 20036 18426
rect 19984 18362 20036 18368
rect 20076 18352 20128 18358
rect 20076 18294 20128 18300
rect 20088 17610 20116 18294
rect 20180 18222 20208 18702
rect 20640 18698 20668 18770
rect 20732 18698 20760 20334
rect 20996 20256 21048 20262
rect 20996 20198 21048 20204
rect 20812 19508 20864 19514
rect 20812 19450 20864 19456
rect 20824 18714 20852 19450
rect 21008 19310 21036 20198
rect 21272 19372 21324 19378
rect 21272 19314 21324 19320
rect 20996 19304 21048 19310
rect 20996 19246 21048 19252
rect 20904 19168 20956 19174
rect 20904 19110 20956 19116
rect 20916 18970 20944 19110
rect 20904 18964 20956 18970
rect 20904 18906 20956 18912
rect 21284 18902 21312 19314
rect 21272 18896 21324 18902
rect 21272 18838 21324 18844
rect 20824 18698 21220 18714
rect 20260 18692 20312 18698
rect 20260 18634 20312 18640
rect 20628 18692 20680 18698
rect 20628 18634 20680 18640
rect 20720 18692 20772 18698
rect 20720 18634 20772 18640
rect 20824 18692 21232 18698
rect 20824 18686 21180 18692
rect 20168 18216 20220 18222
rect 20168 18158 20220 18164
rect 20272 18154 20300 18634
rect 20824 18630 20852 18686
rect 21180 18634 21232 18640
rect 20812 18624 20864 18630
rect 20812 18566 20864 18572
rect 20904 18624 20956 18630
rect 20904 18566 20956 18572
rect 21088 18624 21140 18630
rect 21088 18566 21140 18572
rect 20260 18148 20312 18154
rect 20260 18090 20312 18096
rect 20824 17882 20852 18566
rect 20916 18086 20944 18566
rect 21100 18358 21128 18566
rect 21088 18352 21140 18358
rect 21088 18294 21140 18300
rect 20904 18080 20956 18086
rect 20904 18022 20956 18028
rect 20812 17876 20864 17882
rect 20812 17818 20864 17824
rect 20076 17604 20128 17610
rect 20076 17546 20128 17552
rect 20088 16522 20116 17546
rect 21088 16720 21140 16726
rect 21088 16662 21140 16668
rect 20076 16516 20128 16522
rect 20076 16458 20128 16464
rect 20088 16182 20116 16458
rect 20076 16176 20128 16182
rect 20076 16118 20128 16124
rect 19892 16040 19944 16046
rect 19892 15982 19944 15988
rect 20812 16040 20864 16046
rect 20812 15982 20864 15988
rect 20352 15972 20404 15978
rect 20352 15914 20404 15920
rect 19800 15700 19852 15706
rect 19800 15642 19852 15648
rect 20364 15638 20392 15914
rect 20628 15904 20680 15910
rect 20628 15846 20680 15852
rect 20352 15632 20404 15638
rect 20352 15574 20404 15580
rect 20364 15502 20392 15574
rect 20640 15502 20668 15846
rect 20720 15564 20772 15570
rect 20720 15506 20772 15512
rect 20352 15496 20404 15502
rect 20352 15438 20404 15444
rect 20628 15496 20680 15502
rect 20732 15473 20760 15506
rect 20628 15438 20680 15444
rect 20718 15464 20774 15473
rect 19340 15428 19392 15434
rect 20718 15399 20774 15408
rect 19340 15370 19392 15376
rect 18880 15156 18932 15162
rect 18880 15098 18932 15104
rect 18512 15088 18564 15094
rect 18512 15030 18564 15036
rect 18052 14816 18104 14822
rect 18052 14758 18104 14764
rect 17776 14476 17828 14482
rect 17776 14418 17828 14424
rect 18064 14414 18092 14758
rect 18052 14408 18104 14414
rect 17972 14368 18052 14396
rect 17500 13932 17552 13938
rect 17500 13874 17552 13880
rect 17408 13456 17460 13462
rect 17408 13398 17460 13404
rect 17224 13252 17276 13258
rect 17224 13194 17276 13200
rect 16948 13184 17000 13190
rect 16948 13126 17000 13132
rect 17040 13184 17092 13190
rect 17040 13126 17092 13132
rect 16764 12980 16816 12986
rect 16764 12922 16816 12928
rect 16776 12850 16804 12922
rect 16764 12844 16816 12850
rect 16764 12786 16816 12792
rect 16960 12306 16988 13126
rect 17052 12850 17080 13126
rect 17132 12912 17184 12918
rect 17132 12854 17184 12860
rect 17040 12844 17092 12850
rect 17040 12786 17092 12792
rect 17052 12442 17080 12786
rect 17040 12436 17092 12442
rect 17040 12378 17092 12384
rect 16948 12300 17000 12306
rect 16948 12242 17000 12248
rect 17144 12102 17172 12854
rect 17224 12844 17276 12850
rect 17224 12786 17276 12792
rect 17132 12096 17184 12102
rect 17132 12038 17184 12044
rect 17132 11348 17184 11354
rect 17132 11290 17184 11296
rect 16580 11212 16632 11218
rect 16580 11154 16632 11160
rect 16396 11076 16448 11082
rect 16396 11018 16448 11024
rect 15936 10668 15988 10674
rect 15936 10610 15988 10616
rect 15948 10130 15976 10610
rect 16028 10192 16080 10198
rect 16028 10134 16080 10140
rect 15936 10124 15988 10130
rect 15936 10066 15988 10072
rect 15844 9988 15896 9994
rect 15844 9930 15896 9936
rect 15752 9512 15804 9518
rect 15752 9454 15804 9460
rect 15476 9376 15528 9382
rect 15476 9318 15528 9324
rect 15936 9376 15988 9382
rect 15936 9318 15988 9324
rect 15384 9172 15436 9178
rect 15384 9114 15436 9120
rect 14280 9036 14332 9042
rect 14280 8978 14332 8984
rect 12900 8900 12952 8906
rect 12900 8842 12952 8848
rect 12912 8634 12940 8842
rect 13176 8832 13228 8838
rect 13176 8774 13228 8780
rect 12900 8628 12952 8634
rect 12900 8570 12952 8576
rect 12532 8492 12584 8498
rect 12532 8434 12584 8440
rect 12808 8492 12860 8498
rect 12808 8434 12860 8440
rect 12164 8424 12216 8430
rect 12164 8366 12216 8372
rect 12176 6934 12204 8366
rect 12256 8084 12308 8090
rect 12256 8026 12308 8032
rect 12268 7410 12296 8026
rect 12348 7880 12400 7886
rect 12348 7822 12400 7828
rect 12440 7880 12492 7886
rect 12440 7822 12492 7828
rect 12360 7410 12388 7822
rect 12256 7404 12308 7410
rect 12256 7346 12308 7352
rect 12348 7404 12400 7410
rect 12348 7346 12400 7352
rect 12268 7002 12296 7346
rect 12452 7342 12480 7822
rect 12440 7336 12492 7342
rect 12440 7278 12492 7284
rect 12256 6996 12308 7002
rect 12452 6984 12480 7278
rect 12532 6996 12584 7002
rect 12452 6956 12532 6984
rect 12256 6938 12308 6944
rect 12532 6938 12584 6944
rect 12164 6928 12216 6934
rect 12164 6870 12216 6876
rect 12440 6792 12492 6798
rect 11886 6760 11942 6769
rect 11152 6724 11204 6730
rect 11152 6666 11204 6672
rect 11612 6724 11664 6730
rect 11612 6666 11664 6672
rect 11796 6724 11848 6730
rect 11886 6695 11888 6704
rect 11796 6666 11848 6672
rect 11940 6695 11942 6704
rect 12268 6752 12440 6780
rect 11888 6666 11940 6672
rect 11060 5840 11112 5846
rect 11060 5782 11112 5788
rect 10876 5704 10928 5710
rect 10876 5646 10928 5652
rect 11072 5642 11100 5782
rect 11164 5710 11192 6666
rect 11808 6458 11836 6666
rect 11796 6452 11848 6458
rect 11796 6394 11848 6400
rect 11702 6352 11758 6361
rect 11758 6296 11836 6304
rect 11702 6287 11704 6296
rect 11756 6276 11836 6296
rect 11704 6258 11756 6264
rect 11704 6112 11756 6118
rect 11704 6054 11756 6060
rect 11336 5908 11388 5914
rect 11336 5850 11388 5856
rect 11152 5704 11204 5710
rect 11152 5646 11204 5652
rect 11348 5642 11376 5850
rect 11716 5710 11744 6054
rect 11704 5704 11756 5710
rect 11704 5646 11756 5652
rect 10416 5636 10468 5642
rect 10416 5578 10468 5584
rect 10508 5636 10560 5642
rect 10508 5578 10560 5584
rect 11060 5636 11112 5642
rect 11060 5578 11112 5584
rect 11336 5636 11388 5642
rect 11336 5578 11388 5584
rect 11072 5370 11100 5578
rect 11244 5568 11296 5574
rect 11244 5510 11296 5516
rect 10324 5364 10376 5370
rect 10324 5306 10376 5312
rect 11060 5364 11112 5370
rect 11060 5306 11112 5312
rect 9036 5296 9088 5302
rect 9036 5238 9088 5244
rect 9864 5296 9916 5302
rect 9864 5238 9916 5244
rect 8024 5228 8076 5234
rect 8024 5170 8076 5176
rect 8300 5228 8352 5234
rect 8300 5170 8352 5176
rect 11256 5098 11284 5510
rect 11348 5234 11376 5578
rect 11336 5228 11388 5234
rect 11336 5170 11388 5176
rect 11704 5228 11756 5234
rect 11808 5216 11836 6276
rect 11900 6254 11928 6666
rect 12268 6662 12296 6752
rect 12624 6792 12676 6798
rect 12440 6734 12492 6740
rect 12622 6760 12624 6769
rect 12676 6760 12678 6769
rect 12820 6730 12848 8434
rect 12992 8288 13044 8294
rect 12992 8230 13044 8236
rect 13004 7954 13032 8230
rect 12992 7948 13044 7954
rect 12992 7890 13044 7896
rect 13188 7818 13216 8774
rect 13360 8492 13412 8498
rect 13360 8434 13412 8440
rect 13268 7880 13320 7886
rect 13268 7822 13320 7828
rect 13176 7812 13228 7818
rect 13176 7754 13228 7760
rect 13280 7546 13308 7822
rect 13372 7750 13400 8434
rect 13636 8288 13688 8294
rect 13636 8230 13688 8236
rect 13360 7744 13412 7750
rect 13360 7686 13412 7692
rect 13452 7744 13504 7750
rect 13452 7686 13504 7692
rect 13268 7540 13320 7546
rect 13268 7482 13320 7488
rect 13464 7410 13492 7686
rect 13648 7478 13676 8230
rect 13820 8016 13872 8022
rect 13820 7958 13872 7964
rect 13636 7472 13688 7478
rect 13636 7414 13688 7420
rect 12900 7404 12952 7410
rect 12900 7346 12952 7352
rect 13452 7404 13504 7410
rect 13452 7346 13504 7352
rect 12912 6934 12940 7346
rect 13832 7342 13860 7958
rect 14292 7954 14320 8978
rect 15488 8974 15516 9318
rect 15948 9178 15976 9318
rect 15936 9172 15988 9178
rect 15936 9114 15988 9120
rect 15476 8968 15528 8974
rect 15476 8910 15528 8916
rect 15948 8430 15976 9114
rect 16040 8566 16068 10134
rect 16408 9926 16436 11018
rect 17144 10810 17172 11290
rect 17236 11082 17264 12786
rect 17420 12646 17448 13398
rect 17512 12918 17540 13874
rect 17868 13864 17920 13870
rect 17868 13806 17920 13812
rect 17776 13456 17828 13462
rect 17776 13398 17828 13404
rect 17788 13326 17816 13398
rect 17684 13320 17736 13326
rect 17684 13262 17736 13268
rect 17776 13320 17828 13326
rect 17776 13262 17828 13268
rect 17592 13252 17644 13258
rect 17592 13194 17644 13200
rect 17500 12912 17552 12918
rect 17500 12854 17552 12860
rect 17408 12640 17460 12646
rect 17408 12582 17460 12588
rect 17420 12170 17448 12582
rect 17500 12436 17552 12442
rect 17500 12378 17552 12384
rect 17512 12306 17540 12378
rect 17500 12300 17552 12306
rect 17500 12242 17552 12248
rect 17604 12238 17632 13194
rect 17696 12918 17724 13262
rect 17684 12912 17736 12918
rect 17684 12854 17736 12860
rect 17696 12434 17724 12854
rect 17880 12442 17908 13806
rect 17868 12436 17920 12442
rect 17696 12406 17816 12434
rect 17592 12232 17644 12238
rect 17592 12174 17644 12180
rect 17408 12164 17460 12170
rect 17408 12106 17460 12112
rect 17684 12096 17736 12102
rect 17684 12038 17736 12044
rect 17224 11076 17276 11082
rect 17224 11018 17276 11024
rect 17592 11076 17644 11082
rect 17592 11018 17644 11024
rect 17604 10810 17632 11018
rect 17132 10804 17184 10810
rect 17132 10746 17184 10752
rect 17592 10804 17644 10810
rect 17592 10746 17644 10752
rect 16764 10668 16816 10674
rect 16764 10610 16816 10616
rect 16672 10124 16724 10130
rect 16672 10066 16724 10072
rect 16580 10056 16632 10062
rect 16580 9998 16632 10004
rect 16396 9920 16448 9926
rect 16396 9862 16448 9868
rect 16120 9512 16172 9518
rect 16120 9454 16172 9460
rect 16132 9178 16160 9454
rect 16120 9172 16172 9178
rect 16120 9114 16172 9120
rect 16408 8906 16436 9862
rect 16592 9722 16620 9998
rect 16580 9716 16632 9722
rect 16580 9658 16632 9664
rect 16684 8974 16712 10066
rect 16672 8968 16724 8974
rect 16672 8910 16724 8916
rect 16396 8900 16448 8906
rect 16396 8842 16448 8848
rect 16028 8560 16080 8566
rect 16028 8502 16080 8508
rect 15936 8424 15988 8430
rect 15936 8366 15988 8372
rect 14280 7948 14332 7954
rect 14280 7890 14332 7896
rect 14648 7880 14700 7886
rect 14648 7822 14700 7828
rect 14660 7546 14688 7822
rect 16408 7818 16436 8842
rect 16580 8084 16632 8090
rect 16580 8026 16632 8032
rect 16396 7812 16448 7818
rect 16396 7754 16448 7760
rect 14648 7540 14700 7546
rect 14648 7482 14700 7488
rect 16592 7478 16620 8026
rect 16580 7472 16632 7478
rect 16580 7414 16632 7420
rect 13820 7336 13872 7342
rect 13820 7278 13872 7284
rect 13728 7268 13780 7274
rect 13728 7210 13780 7216
rect 12900 6928 12952 6934
rect 12900 6870 12952 6876
rect 12900 6792 12952 6798
rect 12900 6734 12952 6740
rect 12622 6695 12678 6704
rect 12808 6724 12860 6730
rect 12256 6656 12308 6662
rect 12256 6598 12308 6604
rect 11888 6248 11940 6254
rect 11888 6190 11940 6196
rect 11888 5840 11940 5846
rect 11888 5782 11940 5788
rect 11900 5574 11928 5782
rect 11888 5568 11940 5574
rect 11888 5510 11940 5516
rect 11756 5188 11836 5216
rect 11704 5170 11756 5176
rect 11900 5166 11928 5510
rect 12268 5302 12296 6598
rect 12256 5296 12308 5302
rect 12256 5238 12308 5244
rect 12636 5234 12664 6695
rect 12808 6666 12860 6672
rect 12820 6390 12848 6666
rect 12808 6384 12860 6390
rect 12912 6361 12940 6734
rect 13740 6662 13768 7210
rect 15660 6724 15712 6730
rect 15660 6666 15712 6672
rect 16580 6724 16632 6730
rect 16580 6666 16632 6672
rect 13728 6656 13780 6662
rect 13728 6598 13780 6604
rect 12808 6326 12860 6332
rect 12898 6352 12954 6361
rect 12716 6316 12768 6322
rect 12716 6258 12768 6264
rect 12728 5574 12756 6258
rect 12820 5710 12848 6326
rect 13740 6322 13768 6598
rect 15672 6458 15700 6666
rect 16592 6474 16620 6666
rect 16500 6458 16620 6474
rect 15660 6452 15712 6458
rect 15660 6394 15712 6400
rect 16488 6452 16620 6458
rect 16540 6446 16620 6452
rect 16488 6394 16540 6400
rect 14740 6384 14792 6390
rect 14740 6326 14792 6332
rect 12898 6287 12954 6296
rect 13636 6316 13688 6322
rect 12808 5704 12860 5710
rect 12808 5646 12860 5652
rect 12716 5568 12768 5574
rect 12716 5510 12768 5516
rect 12624 5228 12676 5234
rect 12624 5170 12676 5176
rect 11888 5160 11940 5166
rect 12912 5148 12940 6287
rect 13636 6258 13688 6264
rect 13728 6316 13780 6322
rect 13728 6258 13780 6264
rect 14556 6316 14608 6322
rect 14556 6258 14608 6264
rect 13084 6112 13136 6118
rect 13084 6054 13136 6060
rect 13268 6112 13320 6118
rect 13268 6054 13320 6060
rect 13096 5642 13124 6054
rect 13084 5636 13136 5642
rect 13084 5578 13136 5584
rect 13096 5234 13124 5578
rect 13084 5228 13136 5234
rect 13084 5170 13136 5176
rect 12992 5160 13044 5166
rect 12912 5120 12992 5148
rect 11888 5102 11940 5108
rect 12992 5102 13044 5108
rect 11244 5092 11296 5098
rect 11244 5034 11296 5040
rect 7104 5024 7156 5030
rect 7104 4966 7156 4972
rect 12900 5024 12952 5030
rect 12900 4966 12952 4972
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 12912 4622 12940 4966
rect 13280 4690 13308 6054
rect 13648 5914 13676 6258
rect 13636 5908 13688 5914
rect 13636 5850 13688 5856
rect 14568 5710 14596 6258
rect 14648 6180 14700 6186
rect 14648 6122 14700 6128
rect 14556 5704 14608 5710
rect 14556 5646 14608 5652
rect 14660 5574 14688 6122
rect 14752 5710 14780 6326
rect 16684 6322 16712 8910
rect 16776 8838 16804 10610
rect 17316 10600 17368 10606
rect 17316 10542 17368 10548
rect 17224 9512 17276 9518
rect 17224 9454 17276 9460
rect 17040 8968 17092 8974
rect 17040 8910 17092 8916
rect 16764 8832 16816 8838
rect 16764 8774 16816 8780
rect 17052 8634 17080 8910
rect 17040 8628 17092 8634
rect 17040 8570 17092 8576
rect 17236 8498 17264 9454
rect 17224 8492 17276 8498
rect 17224 8434 17276 8440
rect 17328 8378 17356 10542
rect 17696 10266 17724 12038
rect 17684 10260 17736 10266
rect 17684 10202 17736 10208
rect 17696 9738 17724 10202
rect 17604 9722 17724 9738
rect 17592 9716 17724 9722
rect 17644 9710 17724 9716
rect 17592 9658 17644 9664
rect 17500 9580 17552 9586
rect 17500 9522 17552 9528
rect 17512 9042 17540 9522
rect 17500 9036 17552 9042
rect 17500 8978 17552 8984
rect 17408 8832 17460 8838
rect 17408 8774 17460 8780
rect 17420 8634 17448 8774
rect 17408 8628 17460 8634
rect 17408 8570 17460 8576
rect 17236 8350 17356 8378
rect 16948 7404 17000 7410
rect 16948 7346 17000 7352
rect 17132 7404 17184 7410
rect 17132 7346 17184 7352
rect 16960 7002 16988 7346
rect 16948 6996 17000 7002
rect 16948 6938 17000 6944
rect 17144 6866 17172 7346
rect 17236 7342 17264 8350
rect 17788 8090 17816 12406
rect 17868 12378 17920 12384
rect 17972 11830 18000 14368
rect 18052 14350 18104 14356
rect 18052 13796 18104 13802
rect 18052 13738 18104 13744
rect 18064 13394 18092 13738
rect 18328 13728 18380 13734
rect 18328 13670 18380 13676
rect 18052 13388 18104 13394
rect 18052 13330 18104 13336
rect 18064 11898 18092 13330
rect 18144 13184 18196 13190
rect 18144 13126 18196 13132
rect 18052 11892 18104 11898
rect 18052 11834 18104 11840
rect 17960 11824 18012 11830
rect 17960 11766 18012 11772
rect 18064 11558 18092 11834
rect 18156 11762 18184 13126
rect 18340 12782 18368 13670
rect 18524 13530 18552 15030
rect 18696 14068 18748 14074
rect 18696 14010 18748 14016
rect 18512 13524 18564 13530
rect 18512 13466 18564 13472
rect 18420 13184 18472 13190
rect 18420 13126 18472 13132
rect 18328 12776 18380 12782
rect 18328 12718 18380 12724
rect 18236 12708 18288 12714
rect 18236 12650 18288 12656
rect 18248 12238 18276 12650
rect 18432 12646 18460 13126
rect 18420 12640 18472 12646
rect 18420 12582 18472 12588
rect 18432 12238 18460 12582
rect 18524 12345 18552 13466
rect 18708 12986 18736 14010
rect 18696 12980 18748 12986
rect 18696 12922 18748 12928
rect 18708 12850 18736 12922
rect 18696 12844 18748 12850
rect 18696 12786 18748 12792
rect 18788 12776 18840 12782
rect 18788 12718 18840 12724
rect 18800 12442 18828 12718
rect 18788 12436 18840 12442
rect 18788 12378 18840 12384
rect 18510 12336 18566 12345
rect 18566 12294 18644 12322
rect 18510 12271 18566 12280
rect 18236 12232 18288 12238
rect 18236 12174 18288 12180
rect 18420 12232 18472 12238
rect 18420 12174 18472 12180
rect 18512 12232 18564 12238
rect 18512 12174 18564 12180
rect 18524 11898 18552 12174
rect 18512 11892 18564 11898
rect 18512 11834 18564 11840
rect 18144 11756 18196 11762
rect 18144 11698 18196 11704
rect 17960 11552 18012 11558
rect 17960 11494 18012 11500
rect 18052 11552 18104 11558
rect 18052 11494 18104 11500
rect 17972 10130 18000 11494
rect 18616 10282 18644 12294
rect 18788 12232 18840 12238
rect 18788 12174 18840 12180
rect 18800 11898 18828 12174
rect 18788 11892 18840 11898
rect 18788 11834 18840 11840
rect 18892 11082 18920 15098
rect 19064 12232 19116 12238
rect 19064 12174 19116 12180
rect 19076 11898 19104 12174
rect 19064 11892 19116 11898
rect 19064 11834 19116 11840
rect 18880 11076 18932 11082
rect 18880 11018 18932 11024
rect 19352 11014 19380 15370
rect 20720 15360 20772 15366
rect 20720 15302 20772 15308
rect 20732 15076 20760 15302
rect 20824 15094 20852 15982
rect 20904 15564 20956 15570
rect 20904 15506 20956 15512
rect 20812 15088 20864 15094
rect 20732 15048 20812 15076
rect 20812 15030 20864 15036
rect 19524 14952 19576 14958
rect 19524 14894 19576 14900
rect 19536 14618 19564 14894
rect 20916 14822 20944 15506
rect 21100 15434 21128 16662
rect 21364 16108 21416 16114
rect 21364 16050 21416 16056
rect 21180 15904 21232 15910
rect 21180 15846 21232 15852
rect 21192 15434 21220 15846
rect 21376 15706 21404 16050
rect 21364 15700 21416 15706
rect 21364 15642 21416 15648
rect 21088 15428 21140 15434
rect 21088 15370 21140 15376
rect 21180 15428 21232 15434
rect 21180 15370 21232 15376
rect 21376 15366 21404 15642
rect 20996 15360 21048 15366
rect 20996 15302 21048 15308
rect 21364 15360 21416 15366
rect 21468 15337 21496 22066
rect 21548 21548 21600 21554
rect 21600 21508 21680 21536
rect 21548 21490 21600 21496
rect 21652 21146 21680 21508
rect 21744 21350 21772 22578
rect 22100 22500 22152 22506
rect 22100 22442 22152 22448
rect 22192 22500 22244 22506
rect 22192 22442 22244 22448
rect 22006 21584 22062 21593
rect 22112 21554 22140 22442
rect 22204 21690 22232 22442
rect 22296 22438 22324 23666
rect 22284 22432 22336 22438
rect 22284 22374 22336 22380
rect 22296 22030 22324 22374
rect 22376 22228 22428 22234
rect 22428 22188 22508 22216
rect 22376 22170 22428 22176
rect 22284 22024 22336 22030
rect 22284 21966 22336 21972
rect 22480 21962 22508 22188
rect 22468 21956 22520 21962
rect 22468 21898 22520 21904
rect 22192 21684 22244 21690
rect 22192 21626 22244 21632
rect 22374 21584 22430 21593
rect 22006 21519 22062 21528
rect 22100 21548 22152 21554
rect 21916 21480 21968 21486
rect 21916 21422 21968 21428
rect 21732 21344 21784 21350
rect 21732 21286 21784 21292
rect 21640 21140 21692 21146
rect 21640 21082 21692 21088
rect 21652 20806 21680 21082
rect 21928 21078 21956 21422
rect 21916 21072 21968 21078
rect 21916 21014 21968 21020
rect 21640 20800 21692 20806
rect 21640 20742 21692 20748
rect 21652 18766 21680 20742
rect 22020 20602 22048 21519
rect 22374 21519 22376 21528
rect 22100 21490 22152 21496
rect 22428 21519 22430 21528
rect 22376 21490 22428 21496
rect 22664 21486 22692 23718
rect 22940 23662 22968 24210
rect 23032 24138 23060 24550
rect 23020 24132 23072 24138
rect 23020 24074 23072 24080
rect 22928 23656 22980 23662
rect 22928 23598 22980 23604
rect 23204 23656 23256 23662
rect 23204 23598 23256 23604
rect 23112 22772 23164 22778
rect 23112 22714 23164 22720
rect 23020 22704 23072 22710
rect 23020 22646 23072 22652
rect 22836 22432 22888 22438
rect 22836 22374 22888 22380
rect 22848 22234 22876 22374
rect 22836 22228 22888 22234
rect 22836 22170 22888 22176
rect 22848 22030 22876 22170
rect 22928 22092 22980 22098
rect 22928 22034 22980 22040
rect 22836 22024 22888 22030
rect 22836 21966 22888 21972
rect 22848 21690 22876 21966
rect 22836 21684 22888 21690
rect 22836 21626 22888 21632
rect 22940 21622 22968 22034
rect 23032 21894 23060 22646
rect 23124 22030 23152 22714
rect 23216 22094 23244 23598
rect 23216 22066 23428 22094
rect 23112 22024 23164 22030
rect 23112 21966 23164 21972
rect 23020 21888 23072 21894
rect 23020 21830 23072 21836
rect 22928 21616 22980 21622
rect 22928 21558 22980 21564
rect 22652 21480 22704 21486
rect 22652 21422 22704 21428
rect 22468 21412 22520 21418
rect 22468 21354 22520 21360
rect 22100 21344 22152 21350
rect 22100 21286 22152 21292
rect 22008 20596 22060 20602
rect 22008 20538 22060 20544
rect 22112 20466 22140 21286
rect 22376 21004 22428 21010
rect 22376 20946 22428 20952
rect 22192 20528 22244 20534
rect 22192 20470 22244 20476
rect 22100 20460 22152 20466
rect 22100 20402 22152 20408
rect 22008 19780 22060 19786
rect 22008 19722 22060 19728
rect 22020 19446 22048 19722
rect 22008 19440 22060 19446
rect 22008 19382 22060 19388
rect 22112 19378 22140 20402
rect 22100 19372 22152 19378
rect 22100 19314 22152 19320
rect 21640 18760 21692 18766
rect 21640 18702 21692 18708
rect 21652 18222 21680 18702
rect 22112 18630 22140 19314
rect 22100 18624 22152 18630
rect 22100 18566 22152 18572
rect 22204 18290 22232 20470
rect 22284 19508 22336 19514
rect 22284 19450 22336 19456
rect 22296 18834 22324 19450
rect 22388 19242 22416 20946
rect 22480 20466 22508 21354
rect 22664 21146 22692 21422
rect 23032 21350 23060 21830
rect 23020 21344 23072 21350
rect 23020 21286 23072 21292
rect 22652 21140 22704 21146
rect 22652 21082 22704 21088
rect 22664 20466 22692 21082
rect 23032 20942 23060 21286
rect 23124 21078 23152 21966
rect 23216 21962 23244 22066
rect 23204 21956 23256 21962
rect 23204 21898 23256 21904
rect 23204 21616 23256 21622
rect 23204 21558 23256 21564
rect 23112 21072 23164 21078
rect 23112 21014 23164 21020
rect 23020 20936 23072 20942
rect 23020 20878 23072 20884
rect 22744 20800 22796 20806
rect 22744 20742 22796 20748
rect 22468 20460 22520 20466
rect 22468 20402 22520 20408
rect 22652 20460 22704 20466
rect 22652 20402 22704 20408
rect 22756 20398 22784 20742
rect 23216 20534 23244 21558
rect 23400 20942 23428 22066
rect 23480 21072 23532 21078
rect 23480 21014 23532 21020
rect 23492 20942 23520 21014
rect 23388 20936 23440 20942
rect 23388 20878 23440 20884
rect 23480 20936 23532 20942
rect 23480 20878 23532 20884
rect 23664 20936 23716 20942
rect 23664 20878 23716 20884
rect 23204 20528 23256 20534
rect 23204 20470 23256 20476
rect 22744 20392 22796 20398
rect 22744 20334 22796 20340
rect 22376 19236 22428 19242
rect 22376 19178 22428 19184
rect 22388 18970 22416 19178
rect 22376 18964 22428 18970
rect 22376 18906 22428 18912
rect 22284 18828 22336 18834
rect 22284 18770 22336 18776
rect 22192 18284 22244 18290
rect 22192 18226 22244 18232
rect 22296 18222 22324 18770
rect 23216 18714 23244 20470
rect 23216 18698 23336 18714
rect 23216 18692 23348 18698
rect 23216 18686 23296 18692
rect 21640 18216 21692 18222
rect 21640 18158 21692 18164
rect 22284 18216 22336 18222
rect 22284 18158 22336 18164
rect 21652 17746 21680 18158
rect 21640 17740 21692 17746
rect 21640 17682 21692 17688
rect 22008 17740 22060 17746
rect 22008 17682 22060 17688
rect 22020 16574 22048 17682
rect 22928 16652 22980 16658
rect 22928 16594 22980 16600
rect 22284 16584 22336 16590
rect 22020 16546 22140 16574
rect 21640 16516 21692 16522
rect 21640 16458 21692 16464
rect 21652 15434 21680 16458
rect 22112 16114 22140 16546
rect 22284 16526 22336 16532
rect 22192 16516 22244 16522
rect 22192 16458 22244 16464
rect 22100 16108 22152 16114
rect 22100 16050 22152 16056
rect 22008 15904 22060 15910
rect 22008 15846 22060 15852
rect 21824 15564 21876 15570
rect 21824 15506 21876 15512
rect 21640 15428 21692 15434
rect 21640 15370 21692 15376
rect 21364 15302 21416 15308
rect 21454 15328 21510 15337
rect 20904 14816 20956 14822
rect 20904 14758 20956 14764
rect 19524 14612 19576 14618
rect 19524 14554 19576 14560
rect 21008 14482 21036 15302
rect 21454 15263 21510 15272
rect 21272 14952 21324 14958
rect 21272 14894 21324 14900
rect 21284 14550 21312 14894
rect 21732 14816 21784 14822
rect 21732 14758 21784 14764
rect 21364 14612 21416 14618
rect 21364 14554 21416 14560
rect 21088 14544 21140 14550
rect 21088 14486 21140 14492
rect 21272 14544 21324 14550
rect 21272 14486 21324 14492
rect 20996 14476 21048 14482
rect 20996 14418 21048 14424
rect 20996 14340 21048 14346
rect 20996 14282 21048 14288
rect 21008 14006 21036 14282
rect 20996 14000 21048 14006
rect 20996 13942 21048 13948
rect 21008 13326 21036 13942
rect 21100 13326 21128 14486
rect 21272 13456 21324 13462
rect 21272 13398 21324 13404
rect 20996 13320 21048 13326
rect 20996 13262 21048 13268
rect 21088 13320 21140 13326
rect 21088 13262 21140 13268
rect 20628 13184 20680 13190
rect 20628 13126 20680 13132
rect 19708 12844 19760 12850
rect 19708 12786 19760 12792
rect 19720 12374 19748 12786
rect 19984 12640 20036 12646
rect 19984 12582 20036 12588
rect 19708 12368 19760 12374
rect 19708 12310 19760 12316
rect 19616 12232 19668 12238
rect 19616 12174 19668 12180
rect 19892 12232 19944 12238
rect 19892 12174 19944 12180
rect 19628 11694 19656 12174
rect 19904 11898 19932 12174
rect 19892 11892 19944 11898
rect 19892 11834 19944 11840
rect 19996 11762 20024 12582
rect 20640 12238 20668 13126
rect 21100 12782 21128 13262
rect 21180 13184 21232 13190
rect 21180 13126 21232 13132
rect 20904 12776 20956 12782
rect 20904 12718 20956 12724
rect 21088 12776 21140 12782
rect 21088 12718 21140 12724
rect 20916 12322 20944 12718
rect 20996 12640 21048 12646
rect 20996 12582 21048 12588
rect 20732 12306 20944 12322
rect 20720 12300 20944 12306
rect 20772 12294 20944 12300
rect 20720 12242 20772 12248
rect 20628 12232 20680 12238
rect 20904 12232 20956 12238
rect 20628 12174 20680 12180
rect 20902 12200 20904 12209
rect 20956 12200 20958 12209
rect 20076 12164 20128 12170
rect 20902 12135 20958 12144
rect 20076 12106 20128 12112
rect 19984 11756 20036 11762
rect 19984 11698 20036 11704
rect 19616 11688 19668 11694
rect 19616 11630 19668 11636
rect 19340 11008 19392 11014
rect 19340 10950 19392 10956
rect 18524 10254 18644 10282
rect 17960 10124 18012 10130
rect 17960 10066 18012 10072
rect 17960 9920 18012 9926
rect 17960 9862 18012 9868
rect 17868 9376 17920 9382
rect 17972 9330 18000 9862
rect 17920 9324 18000 9330
rect 17868 9318 18000 9324
rect 18052 9376 18104 9382
rect 18052 9318 18104 9324
rect 17880 9302 18000 9318
rect 17776 8084 17828 8090
rect 17776 8026 17828 8032
rect 17224 7336 17276 7342
rect 17224 7278 17276 7284
rect 17132 6860 17184 6866
rect 17132 6802 17184 6808
rect 17236 6730 17264 7278
rect 18064 6866 18092 9318
rect 18524 7886 18552 10254
rect 19524 10192 19576 10198
rect 19524 10134 19576 10140
rect 18604 10124 18656 10130
rect 18604 10066 18656 10072
rect 18616 8430 18644 10066
rect 19536 10062 19564 10134
rect 19524 10056 19576 10062
rect 19524 9998 19576 10004
rect 18788 9920 18840 9926
rect 18788 9862 18840 9868
rect 18800 9654 18828 9862
rect 18788 9648 18840 9654
rect 18788 9590 18840 9596
rect 18800 8974 18828 9590
rect 19536 9586 19564 9998
rect 19524 9580 19576 9586
rect 19524 9522 19576 9528
rect 18788 8968 18840 8974
rect 18788 8910 18840 8916
rect 19064 8968 19116 8974
rect 19064 8910 19116 8916
rect 18604 8424 18656 8430
rect 18604 8366 18656 8372
rect 18512 7880 18564 7886
rect 18564 7840 18644 7868
rect 18512 7822 18564 7828
rect 18616 7478 18644 7840
rect 18800 7750 18828 8910
rect 18788 7744 18840 7750
rect 18788 7686 18840 7692
rect 18604 7472 18656 7478
rect 18604 7414 18656 7420
rect 18144 7336 18196 7342
rect 18144 7278 18196 7284
rect 18156 6866 18184 7278
rect 18616 7002 18644 7414
rect 18604 6996 18656 7002
rect 18604 6938 18656 6944
rect 18052 6860 18104 6866
rect 18052 6802 18104 6808
rect 18144 6860 18196 6866
rect 18144 6802 18196 6808
rect 17224 6724 17276 6730
rect 17224 6666 17276 6672
rect 14924 6316 14976 6322
rect 14924 6258 14976 6264
rect 15660 6316 15712 6322
rect 15660 6258 15712 6264
rect 16120 6316 16172 6322
rect 16120 6258 16172 6264
rect 16212 6316 16264 6322
rect 16212 6258 16264 6264
rect 16672 6316 16724 6322
rect 16672 6258 16724 6264
rect 14936 5710 14964 6258
rect 15476 6248 15528 6254
rect 15476 6190 15528 6196
rect 15488 5846 15516 6190
rect 15476 5840 15528 5846
rect 15476 5782 15528 5788
rect 14740 5704 14792 5710
rect 14740 5646 14792 5652
rect 14924 5704 14976 5710
rect 14924 5646 14976 5652
rect 13636 5568 13688 5574
rect 13636 5510 13688 5516
rect 14648 5568 14700 5574
rect 14648 5510 14700 5516
rect 13648 5234 13676 5510
rect 14752 5370 14780 5646
rect 14740 5364 14792 5370
rect 14740 5306 14792 5312
rect 13636 5228 13688 5234
rect 13636 5170 13688 5176
rect 13648 5098 13676 5170
rect 14936 5166 14964 5646
rect 15488 5574 15516 5782
rect 15568 5636 15620 5642
rect 15568 5578 15620 5584
rect 15292 5568 15344 5574
rect 15292 5510 15344 5516
rect 15476 5568 15528 5574
rect 15476 5510 15528 5516
rect 15304 5370 15332 5510
rect 15292 5364 15344 5370
rect 15292 5306 15344 5312
rect 14924 5160 14976 5166
rect 14924 5102 14976 5108
rect 13636 5092 13688 5098
rect 13636 5034 13688 5040
rect 13912 5092 13964 5098
rect 13912 5034 13964 5040
rect 13360 5024 13412 5030
rect 13360 4966 13412 4972
rect 13820 5024 13872 5030
rect 13820 4966 13872 4972
rect 13268 4684 13320 4690
rect 13268 4626 13320 4632
rect 12900 4616 12952 4622
rect 12900 4558 12952 4564
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 13372 4146 13400 4966
rect 13832 4162 13860 4966
rect 13740 4146 13860 4162
rect 13924 4146 13952 5034
rect 15108 4480 15160 4486
rect 15108 4422 15160 4428
rect 15120 4214 15148 4422
rect 15304 4282 15332 5306
rect 15580 5302 15608 5578
rect 15568 5296 15620 5302
rect 15568 5238 15620 5244
rect 15672 5234 15700 6258
rect 15936 5704 15988 5710
rect 15936 5646 15988 5652
rect 15948 5370 15976 5646
rect 16132 5574 16160 6258
rect 16224 5914 16252 6258
rect 16396 6248 16448 6254
rect 16396 6190 16448 6196
rect 16212 5908 16264 5914
rect 16212 5850 16264 5856
rect 16408 5846 16436 6190
rect 17236 5846 17264 6666
rect 17316 6656 17368 6662
rect 17316 6598 17368 6604
rect 17500 6656 17552 6662
rect 17500 6598 17552 6604
rect 16396 5840 16448 5846
rect 16396 5782 16448 5788
rect 17224 5840 17276 5846
rect 17224 5782 17276 5788
rect 17328 5778 17356 6598
rect 17512 6458 17540 6598
rect 17500 6452 17552 6458
rect 17500 6394 17552 6400
rect 17500 6248 17552 6254
rect 17500 6190 17552 6196
rect 17512 5914 17540 6190
rect 18064 6186 18092 6802
rect 18800 6390 18828 7686
rect 19076 6798 19104 8910
rect 19064 6792 19116 6798
rect 19064 6734 19116 6740
rect 19076 6474 19104 6734
rect 18984 6446 19104 6474
rect 18788 6384 18840 6390
rect 18788 6326 18840 6332
rect 18984 6186 19012 6446
rect 18052 6180 18104 6186
rect 18052 6122 18104 6128
rect 18972 6180 19024 6186
rect 18972 6122 19024 6128
rect 18788 6112 18840 6118
rect 18788 6054 18840 6060
rect 17500 5908 17552 5914
rect 17500 5850 17552 5856
rect 16672 5772 16724 5778
rect 16672 5714 16724 5720
rect 17316 5772 17368 5778
rect 17316 5714 17368 5720
rect 16580 5704 16632 5710
rect 16580 5646 16632 5652
rect 16120 5568 16172 5574
rect 16120 5510 16172 5516
rect 15936 5364 15988 5370
rect 15936 5306 15988 5312
rect 16592 5302 16620 5646
rect 16684 5370 16712 5714
rect 18800 5642 18828 6054
rect 19536 5710 19564 9522
rect 19628 7546 19656 11630
rect 20088 11218 20116 12106
rect 20444 12096 20496 12102
rect 20444 12038 20496 12044
rect 20260 11756 20312 11762
rect 20260 11698 20312 11704
rect 20168 11688 20220 11694
rect 20168 11630 20220 11636
rect 20180 11354 20208 11630
rect 20272 11354 20300 11698
rect 20168 11348 20220 11354
rect 20168 11290 20220 11296
rect 20260 11348 20312 11354
rect 20260 11290 20312 11296
rect 20352 11280 20404 11286
rect 20272 11228 20352 11234
rect 20272 11222 20404 11228
rect 20076 11212 20128 11218
rect 20076 11154 20128 11160
rect 20272 11206 20392 11222
rect 19892 11144 19944 11150
rect 19892 11086 19944 11092
rect 19904 10810 19932 11086
rect 19892 10804 19944 10810
rect 19892 10746 19944 10752
rect 19904 10266 19932 10746
rect 19892 10260 19944 10266
rect 19892 10202 19944 10208
rect 20088 10062 20116 11154
rect 20272 11150 20300 11206
rect 20456 11150 20484 12038
rect 21008 11898 21036 12582
rect 21100 12481 21128 12718
rect 21192 12646 21220 13126
rect 21180 12640 21232 12646
rect 21180 12582 21232 12588
rect 21086 12472 21142 12481
rect 21086 12407 21142 12416
rect 21088 12300 21140 12306
rect 21088 12242 21140 12248
rect 21100 12102 21128 12242
rect 21284 12102 21312 13398
rect 21376 12986 21404 14554
rect 21744 14414 21772 14758
rect 21640 14408 21692 14414
rect 21640 14350 21692 14356
rect 21732 14408 21784 14414
rect 21732 14350 21784 14356
rect 21456 14068 21508 14074
rect 21456 14010 21508 14016
rect 21468 13326 21496 14010
rect 21456 13320 21508 13326
rect 21456 13262 21508 13268
rect 21548 13320 21600 13326
rect 21548 13262 21600 13268
rect 21454 13152 21510 13161
rect 21454 13087 21510 13096
rect 21468 12986 21496 13087
rect 21364 12980 21416 12986
rect 21364 12922 21416 12928
rect 21456 12980 21508 12986
rect 21456 12922 21508 12928
rect 21088 12096 21140 12102
rect 21088 12038 21140 12044
rect 21272 12096 21324 12102
rect 21272 12038 21324 12044
rect 20996 11892 21048 11898
rect 20996 11834 21048 11840
rect 21376 11694 21404 12922
rect 21560 12434 21588 13262
rect 21652 12986 21680 14350
rect 21640 12980 21692 12986
rect 21640 12922 21692 12928
rect 21744 12434 21772 14350
rect 21468 12406 21588 12434
rect 21652 12406 21772 12434
rect 21468 12374 21496 12406
rect 21456 12368 21508 12374
rect 21456 12310 21508 12316
rect 21468 12238 21496 12310
rect 21652 12306 21680 12406
rect 21640 12300 21692 12306
rect 21640 12242 21692 12248
rect 21456 12232 21508 12238
rect 21456 12174 21508 12180
rect 21364 11688 21416 11694
rect 21364 11630 21416 11636
rect 21836 11626 21864 15506
rect 21916 14816 21968 14822
rect 21916 14758 21968 14764
rect 21928 14414 21956 14758
rect 22020 14618 22048 15846
rect 22204 15094 22232 16458
rect 22296 15978 22324 16526
rect 22652 16040 22704 16046
rect 22652 15982 22704 15988
rect 22284 15972 22336 15978
rect 22284 15914 22336 15920
rect 22296 15178 22324 15914
rect 22664 15638 22692 15982
rect 22652 15632 22704 15638
rect 22652 15574 22704 15580
rect 22468 15428 22520 15434
rect 22388 15388 22468 15416
rect 22388 15178 22416 15388
rect 22468 15370 22520 15376
rect 22296 15150 22416 15178
rect 22192 15088 22244 15094
rect 22244 15036 22324 15042
rect 22192 15030 22324 15036
rect 22204 15014 22324 15030
rect 22192 14952 22244 14958
rect 22192 14894 22244 14900
rect 22008 14612 22060 14618
rect 22008 14554 22060 14560
rect 22204 14414 22232 14894
rect 22296 14822 22324 15014
rect 22284 14816 22336 14822
rect 22284 14758 22336 14764
rect 22296 14414 22324 14758
rect 22388 14618 22416 15150
rect 22664 15042 22692 15574
rect 22572 15026 22692 15042
rect 22940 15026 22968 16594
rect 23216 16454 23244 18686
rect 23296 18634 23348 18640
rect 23400 18086 23428 20878
rect 23676 20602 23704 20878
rect 23664 20596 23716 20602
rect 23664 20538 23716 20544
rect 23388 18080 23440 18086
rect 23388 18022 23440 18028
rect 23204 16448 23256 16454
rect 23204 16390 23256 16396
rect 23216 16182 23244 16390
rect 23204 16176 23256 16182
rect 23204 16118 23256 16124
rect 23388 16176 23440 16182
rect 23388 16118 23440 16124
rect 23112 16040 23164 16046
rect 23112 15982 23164 15988
rect 23124 15706 23152 15982
rect 23204 15904 23256 15910
rect 23204 15846 23256 15852
rect 23296 15904 23348 15910
rect 23296 15846 23348 15852
rect 23112 15700 23164 15706
rect 23112 15642 23164 15648
rect 23216 15638 23244 15846
rect 23204 15632 23256 15638
rect 23204 15574 23256 15580
rect 23308 15502 23336 15846
rect 23400 15706 23428 16118
rect 23388 15700 23440 15706
rect 23388 15642 23440 15648
rect 23296 15496 23348 15502
rect 23216 15444 23296 15450
rect 23216 15438 23348 15444
rect 23216 15422 23336 15438
rect 23216 15094 23244 15422
rect 23296 15360 23348 15366
rect 23296 15302 23348 15308
rect 23204 15088 23256 15094
rect 23204 15030 23256 15036
rect 22560 15020 22692 15026
rect 22612 15014 22692 15020
rect 22928 15020 22980 15026
rect 22560 14962 22612 14968
rect 22928 14962 22980 14968
rect 22560 14884 22612 14890
rect 22612 14844 22692 14872
rect 22560 14826 22612 14832
rect 22376 14612 22428 14618
rect 22376 14554 22428 14560
rect 21916 14408 21968 14414
rect 22192 14408 22244 14414
rect 21968 14368 22048 14396
rect 21916 14350 21968 14356
rect 21916 13932 21968 13938
rect 21916 13874 21968 13880
rect 21928 13530 21956 13874
rect 21916 13524 21968 13530
rect 21916 13466 21968 13472
rect 21928 12782 21956 13466
rect 22020 13326 22048 14368
rect 22192 14350 22244 14356
rect 22284 14408 22336 14414
rect 22284 14350 22336 14356
rect 22664 13938 22692 14844
rect 22940 14074 22968 14962
rect 23020 14408 23072 14414
rect 23216 14362 23244 15030
rect 23308 14618 23336 15302
rect 23400 15042 23428 15642
rect 24492 15428 24544 15434
rect 24492 15370 24544 15376
rect 24308 15360 24360 15366
rect 24504 15337 24532 15370
rect 24308 15302 24360 15308
rect 24490 15328 24546 15337
rect 24320 15094 24348 15302
rect 24490 15263 24546 15272
rect 24308 15088 24360 15094
rect 23400 15026 23520 15042
rect 24308 15030 24360 15036
rect 23400 15020 23532 15026
rect 23400 15014 23480 15020
rect 23480 14962 23532 14968
rect 24860 14952 24912 14958
rect 24860 14894 24912 14900
rect 23296 14612 23348 14618
rect 23296 14554 23348 14560
rect 23020 14350 23072 14356
rect 22928 14068 22980 14074
rect 22928 14010 22980 14016
rect 23032 13954 23060 14350
rect 23124 14346 23244 14362
rect 23388 14408 23440 14414
rect 23388 14350 23440 14356
rect 23112 14340 23244 14346
rect 23164 14334 23244 14340
rect 23112 14282 23164 14288
rect 22192 13932 22244 13938
rect 22192 13874 22244 13880
rect 22652 13932 22704 13938
rect 22652 13874 22704 13880
rect 22756 13926 23060 13954
rect 22204 13569 22232 13874
rect 22756 13870 22784 13926
rect 22744 13864 22796 13870
rect 22744 13806 22796 13812
rect 22928 13864 22980 13870
rect 22928 13806 22980 13812
rect 22468 13796 22520 13802
rect 22468 13738 22520 13744
rect 22284 13728 22336 13734
rect 22284 13670 22336 13676
rect 22190 13560 22246 13569
rect 22296 13530 22324 13670
rect 22480 13530 22508 13738
rect 22560 13728 22612 13734
rect 22560 13670 22612 13676
rect 22836 13728 22888 13734
rect 22836 13670 22888 13676
rect 22190 13495 22246 13504
rect 22284 13524 22336 13530
rect 22100 13456 22152 13462
rect 22098 13424 22100 13433
rect 22152 13424 22154 13433
rect 22098 13359 22154 13368
rect 22008 13320 22060 13326
rect 22008 13262 22060 13268
rect 22100 13184 22152 13190
rect 22098 13152 22100 13161
rect 22152 13152 22154 13161
rect 22098 13087 22154 13096
rect 21916 12776 21968 12782
rect 21916 12718 21968 12724
rect 22006 12472 22062 12481
rect 22006 12407 22062 12416
rect 22100 12436 22152 12442
rect 22020 12306 22048 12407
rect 22100 12378 22152 12384
rect 22008 12300 22060 12306
rect 22008 12242 22060 12248
rect 21916 12232 21968 12238
rect 21916 12174 21968 12180
rect 21928 12102 21956 12174
rect 21916 12096 21968 12102
rect 21916 12038 21968 12044
rect 21916 11756 21968 11762
rect 21916 11698 21968 11704
rect 21824 11620 21876 11626
rect 21824 11562 21876 11568
rect 21364 11552 21416 11558
rect 21364 11494 21416 11500
rect 21376 11218 21404 11494
rect 21364 11212 21416 11218
rect 21364 11154 21416 11160
rect 20260 11144 20312 11150
rect 20260 11086 20312 11092
rect 20444 11144 20496 11150
rect 20444 11086 20496 11092
rect 20904 11144 20956 11150
rect 20904 11086 20956 11092
rect 21548 11144 21600 11150
rect 21548 11086 21600 11092
rect 20272 10130 20300 11086
rect 20444 11008 20496 11014
rect 20444 10950 20496 10956
rect 20352 10192 20404 10198
rect 20352 10134 20404 10140
rect 20260 10124 20312 10130
rect 20260 10066 20312 10072
rect 20076 10056 20128 10062
rect 20076 9998 20128 10004
rect 19800 9988 19852 9994
rect 19800 9930 19852 9936
rect 19812 9586 19840 9930
rect 20168 9920 20220 9926
rect 20168 9862 20220 9868
rect 20180 9722 20208 9862
rect 20168 9716 20220 9722
rect 20168 9658 20220 9664
rect 19800 9580 19852 9586
rect 19800 9522 19852 9528
rect 19892 9580 19944 9586
rect 19892 9522 19944 9528
rect 20076 9580 20128 9586
rect 20076 9522 20128 9528
rect 20260 9580 20312 9586
rect 20260 9522 20312 9528
rect 19904 9382 19932 9522
rect 19892 9376 19944 9382
rect 19892 9318 19944 9324
rect 19904 9042 19932 9318
rect 19892 9036 19944 9042
rect 19892 8978 19944 8984
rect 20088 8974 20116 9522
rect 20076 8968 20128 8974
rect 20076 8910 20128 8916
rect 20272 8634 20300 9522
rect 20364 9450 20392 10134
rect 20456 10062 20484 10950
rect 20916 10810 20944 11086
rect 21560 10810 21588 11086
rect 20904 10804 20956 10810
rect 20904 10746 20956 10752
rect 21548 10804 21600 10810
rect 21548 10746 21600 10752
rect 21836 10742 21864 11562
rect 21928 11354 21956 11698
rect 22112 11354 22140 12378
rect 22204 12374 22232 13495
rect 22284 13466 22336 13472
rect 22468 13524 22520 13530
rect 22468 13466 22520 13472
rect 22192 12368 22244 12374
rect 22192 12310 22244 12316
rect 22296 12102 22324 13466
rect 22376 13320 22428 13326
rect 22480 13308 22508 13466
rect 22428 13280 22508 13308
rect 22376 13262 22428 13268
rect 22480 12986 22508 13280
rect 22572 13025 22600 13670
rect 22650 13288 22706 13297
rect 22650 13223 22652 13232
rect 22704 13223 22706 13232
rect 22652 13194 22704 13200
rect 22558 13016 22614 13025
rect 22468 12980 22520 12986
rect 22558 12951 22614 12960
rect 22468 12922 22520 12928
rect 22848 12850 22876 13670
rect 22940 13161 22968 13806
rect 23032 13530 23060 13926
rect 23020 13524 23072 13530
rect 23020 13466 23072 13472
rect 23124 13394 23152 14282
rect 23400 14006 23428 14350
rect 23480 14068 23532 14074
rect 23480 14010 23532 14016
rect 23388 14000 23440 14006
rect 23388 13942 23440 13948
rect 23296 13932 23348 13938
rect 23296 13874 23348 13880
rect 23202 13560 23258 13569
rect 23202 13495 23204 13504
rect 23256 13495 23258 13504
rect 23204 13466 23256 13472
rect 23202 13424 23258 13433
rect 23112 13388 23164 13394
rect 23202 13359 23258 13368
rect 23112 13330 23164 13336
rect 23216 13326 23244 13359
rect 23308 13326 23336 13874
rect 23204 13320 23256 13326
rect 23296 13320 23348 13326
rect 23204 13262 23256 13268
rect 23294 13288 23296 13297
rect 23348 13288 23350 13297
rect 22926 13152 22982 13161
rect 22926 13087 22982 13096
rect 22560 12844 22612 12850
rect 22560 12786 22612 12792
rect 22836 12844 22888 12850
rect 22836 12786 22888 12792
rect 22376 12708 22428 12714
rect 22376 12650 22428 12656
rect 22388 12442 22416 12650
rect 22468 12640 22520 12646
rect 22468 12582 22520 12588
rect 22480 12442 22508 12582
rect 22376 12436 22428 12442
rect 22376 12378 22428 12384
rect 22468 12436 22520 12442
rect 22468 12378 22520 12384
rect 22376 12300 22428 12306
rect 22376 12242 22428 12248
rect 22468 12300 22520 12306
rect 22468 12242 22520 12248
rect 22284 12096 22336 12102
rect 22284 12038 22336 12044
rect 22192 11756 22244 11762
rect 22192 11698 22244 11704
rect 21916 11348 21968 11354
rect 21916 11290 21968 11296
rect 22100 11348 22152 11354
rect 22100 11290 22152 11296
rect 22204 11286 22232 11698
rect 22388 11694 22416 12242
rect 22376 11688 22428 11694
rect 22376 11630 22428 11636
rect 22480 11626 22508 12242
rect 22468 11620 22520 11626
rect 22468 11562 22520 11568
rect 22192 11280 22244 11286
rect 22192 11222 22244 11228
rect 22284 11212 22336 11218
rect 22284 11154 22336 11160
rect 22100 11144 22152 11150
rect 22100 11086 22152 11092
rect 21824 10736 21876 10742
rect 21824 10678 21876 10684
rect 21272 10668 21324 10674
rect 21272 10610 21324 10616
rect 21180 10464 21232 10470
rect 21180 10406 21232 10412
rect 20720 10124 20772 10130
rect 20720 10066 20772 10072
rect 20444 10056 20496 10062
rect 20444 9998 20496 10004
rect 20628 9512 20680 9518
rect 20628 9454 20680 9460
rect 20352 9444 20404 9450
rect 20352 9386 20404 9392
rect 20640 9178 20668 9454
rect 20628 9172 20680 9178
rect 20628 9114 20680 9120
rect 20732 9058 20760 10066
rect 21192 9586 21220 10406
rect 21284 9722 21312 10610
rect 21548 10600 21600 10606
rect 21548 10542 21600 10548
rect 21272 9716 21324 9722
rect 21272 9658 21324 9664
rect 21180 9580 21232 9586
rect 21180 9522 21232 9528
rect 21192 9450 21220 9522
rect 21560 9518 21588 10542
rect 21836 10266 21864 10678
rect 21824 10260 21876 10266
rect 21824 10202 21876 10208
rect 21548 9512 21600 9518
rect 21548 9454 21600 9460
rect 20996 9444 21048 9450
rect 20996 9386 21048 9392
rect 21180 9444 21232 9450
rect 21180 9386 21232 9392
rect 20640 9042 20760 9058
rect 20628 9036 20760 9042
rect 20680 9030 20760 9036
rect 20628 8978 20680 8984
rect 21008 8974 21036 9386
rect 20720 8968 20772 8974
rect 20720 8910 20772 8916
rect 20996 8968 21048 8974
rect 20996 8910 21048 8916
rect 20444 8900 20496 8906
rect 20444 8842 20496 8848
rect 20260 8628 20312 8634
rect 20260 8570 20312 8576
rect 20456 8498 20484 8842
rect 20732 8498 20760 8910
rect 21192 8838 21220 9386
rect 21560 9382 21588 9454
rect 21548 9376 21600 9382
rect 21548 9318 21600 9324
rect 21456 8968 21508 8974
rect 21456 8910 21508 8916
rect 21180 8832 21232 8838
rect 21180 8774 21232 8780
rect 21468 8634 21496 8910
rect 21456 8628 21508 8634
rect 21456 8570 21508 8576
rect 20444 8492 20496 8498
rect 20444 8434 20496 8440
rect 20720 8492 20772 8498
rect 20720 8434 20772 8440
rect 19616 7540 19668 7546
rect 19616 7482 19668 7488
rect 20732 7002 20760 8434
rect 21364 7268 21416 7274
rect 21364 7210 21416 7216
rect 19984 6996 20036 7002
rect 19984 6938 20036 6944
rect 20720 6996 20772 7002
rect 20720 6938 20772 6944
rect 19616 6792 19668 6798
rect 19616 6734 19668 6740
rect 19628 6458 19656 6734
rect 19996 6730 20024 6938
rect 19984 6724 20036 6730
rect 19984 6666 20036 6672
rect 19616 6452 19668 6458
rect 19616 6394 19668 6400
rect 19524 5704 19576 5710
rect 19524 5646 19576 5652
rect 19996 5642 20024 6666
rect 20732 6458 20760 6938
rect 20812 6860 20864 6866
rect 20812 6802 20864 6808
rect 20720 6452 20772 6458
rect 20720 6394 20772 6400
rect 20824 6254 20852 6802
rect 21376 6322 21404 7210
rect 21546 6488 21602 6497
rect 21546 6423 21548 6432
rect 21600 6423 21602 6432
rect 21548 6394 21600 6400
rect 21364 6316 21416 6322
rect 21364 6258 21416 6264
rect 20812 6248 20864 6254
rect 20812 6190 20864 6196
rect 21088 6248 21140 6254
rect 21088 6190 21140 6196
rect 20824 5778 20852 6190
rect 21100 5914 21128 6190
rect 21088 5908 21140 5914
rect 21088 5850 21140 5856
rect 20812 5772 20864 5778
rect 20812 5714 20864 5720
rect 18788 5636 18840 5642
rect 18788 5578 18840 5584
rect 19984 5636 20036 5642
rect 19984 5578 20036 5584
rect 18696 5568 18748 5574
rect 18696 5510 18748 5516
rect 16672 5364 16724 5370
rect 16672 5306 16724 5312
rect 16580 5296 16632 5302
rect 16580 5238 16632 5244
rect 15660 5228 15712 5234
rect 15660 5170 15712 5176
rect 15292 4276 15344 4282
rect 15292 4218 15344 4224
rect 15108 4208 15160 4214
rect 15108 4150 15160 4156
rect 13360 4140 13412 4146
rect 13360 4082 13412 4088
rect 13728 4140 13860 4146
rect 13780 4134 13860 4140
rect 13728 4082 13780 4088
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 13832 3534 13860 4134
rect 13912 4140 13964 4146
rect 13912 4082 13964 4088
rect 14924 4140 14976 4146
rect 14924 4082 14976 4088
rect 13924 3602 13952 4082
rect 14188 4072 14240 4078
rect 14188 4014 14240 4020
rect 14200 3738 14228 4014
rect 14936 3738 14964 4082
rect 14188 3732 14240 3738
rect 14188 3674 14240 3680
rect 14924 3732 14976 3738
rect 14924 3674 14976 3680
rect 15120 3602 15148 4150
rect 18708 4146 18736 5510
rect 19996 5370 20024 5578
rect 19984 5364 20036 5370
rect 19984 5306 20036 5312
rect 21560 5234 21588 6394
rect 21836 5778 21864 10202
rect 22112 10198 22140 11086
rect 22100 10192 22152 10198
rect 22100 10134 22152 10140
rect 22296 9450 22324 11154
rect 22376 11144 22428 11150
rect 22376 11086 22428 11092
rect 22388 10810 22416 11086
rect 22572 11082 22600 12786
rect 22834 12744 22890 12753
rect 22834 12679 22890 12688
rect 22848 12646 22876 12679
rect 22836 12640 22888 12646
rect 22836 12582 22888 12588
rect 22836 12164 22888 12170
rect 22940 12152 22968 13087
rect 23020 12844 23072 12850
rect 23020 12786 23072 12792
rect 23112 12844 23164 12850
rect 23112 12786 23164 12792
rect 22888 12124 22968 12152
rect 22836 12106 22888 12112
rect 23032 11082 23060 12786
rect 23124 11694 23152 12786
rect 23216 12628 23244 13262
rect 23294 13223 23350 13232
rect 23400 12850 23428 13942
rect 23492 13326 23520 14010
rect 23664 13864 23716 13870
rect 23664 13806 23716 13812
rect 23676 13530 23704 13806
rect 23664 13524 23716 13530
rect 23664 13466 23716 13472
rect 24492 13388 24544 13394
rect 24492 13330 24544 13336
rect 23480 13320 23532 13326
rect 23480 13262 23532 13268
rect 24032 13320 24084 13326
rect 24032 13262 24084 13268
rect 23492 12918 23520 13262
rect 23572 13252 23624 13258
rect 23572 13194 23624 13200
rect 23480 12912 23532 12918
rect 23480 12854 23532 12860
rect 23388 12844 23440 12850
rect 23388 12786 23440 12792
rect 23584 12646 23612 13194
rect 24044 12918 24072 13262
rect 24308 13184 24360 13190
rect 24308 13126 24360 13132
rect 24032 12912 24084 12918
rect 24032 12854 24084 12860
rect 23388 12640 23440 12646
rect 23216 12600 23388 12628
rect 23388 12582 23440 12588
rect 23572 12640 23624 12646
rect 23572 12582 23624 12588
rect 23202 12336 23258 12345
rect 23202 12271 23258 12280
rect 23216 12170 23244 12271
rect 23400 12209 23428 12582
rect 24044 12442 24072 12854
rect 24320 12850 24348 13126
rect 24504 12850 24532 13330
rect 24584 13320 24636 13326
rect 24584 13262 24636 13268
rect 24308 12844 24360 12850
rect 24308 12786 24360 12792
rect 24492 12844 24544 12850
rect 24492 12786 24544 12792
rect 24032 12436 24084 12442
rect 24032 12378 24084 12384
rect 23386 12200 23442 12209
rect 23204 12164 23256 12170
rect 23386 12135 23442 12144
rect 23204 12106 23256 12112
rect 23112 11688 23164 11694
rect 23112 11630 23164 11636
rect 22560 11076 22612 11082
rect 22560 11018 22612 11024
rect 23020 11076 23072 11082
rect 23020 11018 23072 11024
rect 22376 10804 22428 10810
rect 22376 10746 22428 10752
rect 23400 10674 23428 12135
rect 24596 11898 24624 13262
rect 24768 13184 24820 13190
rect 24768 13126 24820 13132
rect 24780 13025 24808 13126
rect 24766 13016 24822 13025
rect 24766 12951 24822 12960
rect 24872 12306 24900 14894
rect 24860 12300 24912 12306
rect 24860 12242 24912 12248
rect 24584 11892 24636 11898
rect 24584 11834 24636 11840
rect 22468 10668 22520 10674
rect 22468 10610 22520 10616
rect 23388 10668 23440 10674
rect 23388 10610 23440 10616
rect 22284 9444 22336 9450
rect 22284 9386 22336 9392
rect 22480 9110 22508 10610
rect 22652 10056 22704 10062
rect 22652 9998 22704 10004
rect 22664 9654 22692 9998
rect 22652 9648 22704 9654
rect 22652 9590 22704 9596
rect 22468 9104 22520 9110
rect 22468 9046 22520 9052
rect 24676 6316 24728 6322
rect 24676 6258 24728 6264
rect 21824 5772 21876 5778
rect 21824 5714 21876 5720
rect 21548 5228 21600 5234
rect 21548 5170 21600 5176
rect 18696 4140 18748 4146
rect 18696 4082 18748 4088
rect 15200 3936 15252 3942
rect 15200 3878 15252 3884
rect 13912 3596 13964 3602
rect 13912 3538 13964 3544
rect 15108 3596 15160 3602
rect 15108 3538 15160 3544
rect 15212 3534 15240 3878
rect 24688 3738 24716 6258
rect 24676 3732 24728 3738
rect 24676 3674 24728 3680
rect 13820 3528 13872 3534
rect 13820 3470 13872 3476
rect 15200 3528 15252 3534
rect 24860 3528 24912 3534
rect 15200 3470 15252 3476
rect 24858 3496 24860 3505
rect 24912 3496 24914 3505
rect 24858 3431 24914 3440
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
<< via2 >>
rect 4880 26138 4936 26140
rect 4960 26138 5016 26140
rect 5040 26138 5096 26140
rect 5120 26138 5176 26140
rect 4880 26086 4926 26138
rect 4926 26086 4936 26138
rect 4960 26086 4990 26138
rect 4990 26086 5002 26138
rect 5002 26086 5016 26138
rect 5040 26086 5054 26138
rect 5054 26086 5066 26138
rect 5066 26086 5096 26138
rect 5120 26086 5130 26138
rect 5130 26086 5176 26138
rect 4880 26084 4936 26086
rect 4960 26084 5016 26086
rect 5040 26084 5096 26086
rect 5120 26084 5176 26086
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 110 24248 166 24304
rect 1398 15000 1454 15056
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4880 25050 4936 25052
rect 4960 25050 5016 25052
rect 5040 25050 5096 25052
rect 5120 25050 5176 25052
rect 4880 24998 4926 25050
rect 4926 24998 4936 25050
rect 4960 24998 4990 25050
rect 4990 24998 5002 25050
rect 5002 24998 5016 25050
rect 5040 24998 5054 25050
rect 5054 24998 5066 25050
rect 5066 24998 5096 25050
rect 5120 24998 5130 25050
rect 5130 24998 5176 25050
rect 4880 24996 4936 24998
rect 4960 24996 5016 24998
rect 5040 24996 5096 24998
rect 5120 24996 5176 24998
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4880 23962 4936 23964
rect 4960 23962 5016 23964
rect 5040 23962 5096 23964
rect 5120 23962 5176 23964
rect 4880 23910 4926 23962
rect 4926 23910 4936 23962
rect 4960 23910 4990 23962
rect 4990 23910 5002 23962
rect 5002 23910 5016 23962
rect 5040 23910 5054 23962
rect 5054 23910 5066 23962
rect 5066 23910 5096 23962
rect 5120 23910 5130 23962
rect 5130 23910 5176 23962
rect 4880 23908 4936 23910
rect 4960 23908 5016 23910
rect 5040 23908 5096 23910
rect 5120 23908 5176 23910
rect 4880 22874 4936 22876
rect 4960 22874 5016 22876
rect 5040 22874 5096 22876
rect 5120 22874 5176 22876
rect 4880 22822 4926 22874
rect 4926 22822 4936 22874
rect 4960 22822 4990 22874
rect 4990 22822 5002 22874
rect 5002 22822 5016 22874
rect 5040 22822 5054 22874
rect 5054 22822 5066 22874
rect 5066 22822 5096 22874
rect 5120 22822 5130 22874
rect 5130 22822 5176 22874
rect 4880 22820 4936 22822
rect 4960 22820 5016 22822
rect 5040 22820 5096 22822
rect 5120 22820 5176 22822
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4880 21786 4936 21788
rect 4960 21786 5016 21788
rect 5040 21786 5096 21788
rect 5120 21786 5176 21788
rect 4880 21734 4926 21786
rect 4926 21734 4936 21786
rect 4960 21734 4990 21786
rect 4990 21734 5002 21786
rect 5002 21734 5016 21786
rect 5040 21734 5054 21786
rect 5054 21734 5066 21786
rect 5066 21734 5096 21786
rect 5120 21734 5130 21786
rect 5130 21734 5176 21786
rect 4880 21732 4936 21734
rect 4960 21732 5016 21734
rect 5040 21732 5096 21734
rect 5120 21732 5176 21734
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 7470 24384 7526 24440
rect 8206 24692 8208 24712
rect 8208 24692 8260 24712
rect 8260 24692 8262 24712
rect 8206 24656 8262 24692
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 846 14184 902 14240
rect 846 11500 848 11520
rect 848 11500 900 11520
rect 900 11500 902 11520
rect 846 11464 902 11500
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4880 20698 4936 20700
rect 4960 20698 5016 20700
rect 5040 20698 5096 20700
rect 5120 20698 5176 20700
rect 4880 20646 4926 20698
rect 4926 20646 4936 20698
rect 4960 20646 4990 20698
rect 4990 20646 5002 20698
rect 5002 20646 5016 20698
rect 5040 20646 5054 20698
rect 5054 20646 5066 20698
rect 5066 20646 5096 20698
rect 5120 20646 5130 20698
rect 5130 20646 5176 20698
rect 4880 20644 4936 20646
rect 4960 20644 5016 20646
rect 5040 20644 5096 20646
rect 5120 20644 5176 20646
rect 4880 19610 4936 19612
rect 4960 19610 5016 19612
rect 5040 19610 5096 19612
rect 5120 19610 5176 19612
rect 4880 19558 4926 19610
rect 4926 19558 4936 19610
rect 4960 19558 4990 19610
rect 4990 19558 5002 19610
rect 5002 19558 5016 19610
rect 5040 19558 5054 19610
rect 5054 19558 5066 19610
rect 5066 19558 5096 19610
rect 5120 19558 5130 19610
rect 5130 19558 5176 19610
rect 4880 19556 4936 19558
rect 4960 19556 5016 19558
rect 5040 19556 5096 19558
rect 5120 19556 5176 19558
rect 9034 24656 9090 24712
rect 9402 24384 9458 24440
rect 4880 18522 4936 18524
rect 4960 18522 5016 18524
rect 5040 18522 5096 18524
rect 5120 18522 5176 18524
rect 4880 18470 4926 18522
rect 4926 18470 4936 18522
rect 4960 18470 4990 18522
rect 4990 18470 5002 18522
rect 5002 18470 5016 18522
rect 5040 18470 5054 18522
rect 5054 18470 5066 18522
rect 5066 18470 5096 18522
rect 5120 18470 5130 18522
rect 5130 18470 5176 18522
rect 4880 18468 4936 18470
rect 4960 18468 5016 18470
rect 5040 18468 5096 18470
rect 5120 18468 5176 18470
rect 8850 21936 8906 21992
rect 9770 22480 9826 22536
rect 10138 22480 10194 22536
rect 4880 17434 4936 17436
rect 4960 17434 5016 17436
rect 5040 17434 5096 17436
rect 5120 17434 5176 17436
rect 4880 17382 4926 17434
rect 4926 17382 4936 17434
rect 4960 17382 4990 17434
rect 4990 17382 5002 17434
rect 5002 17382 5016 17434
rect 5040 17382 5054 17434
rect 5054 17382 5066 17434
rect 5066 17382 5096 17434
rect 5120 17382 5130 17434
rect 5130 17382 5176 17434
rect 4880 17380 4936 17382
rect 4960 17380 5016 17382
rect 5040 17380 5096 17382
rect 5120 17380 5176 17382
rect 4880 16346 4936 16348
rect 4960 16346 5016 16348
rect 5040 16346 5096 16348
rect 5120 16346 5176 16348
rect 4880 16294 4926 16346
rect 4926 16294 4936 16346
rect 4960 16294 4990 16346
rect 4990 16294 5002 16346
rect 5002 16294 5016 16346
rect 5040 16294 5054 16346
rect 5054 16294 5066 16346
rect 5066 16294 5096 16346
rect 5120 16294 5130 16346
rect 5130 16294 5176 16346
rect 4880 16292 4936 16294
rect 4960 16292 5016 16294
rect 5040 16292 5096 16294
rect 5120 16292 5176 16294
rect 4880 15258 4936 15260
rect 4960 15258 5016 15260
rect 5040 15258 5096 15260
rect 5120 15258 5176 15260
rect 4880 15206 4926 15258
rect 4926 15206 4936 15258
rect 4960 15206 4990 15258
rect 4990 15206 5002 15258
rect 5002 15206 5016 15258
rect 5040 15206 5054 15258
rect 5054 15206 5066 15258
rect 5066 15206 5096 15258
rect 5120 15206 5130 15258
rect 5130 15206 5176 15258
rect 4880 15204 4936 15206
rect 4960 15204 5016 15206
rect 5040 15204 5096 15206
rect 5120 15204 5176 15206
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4880 14170 4936 14172
rect 4960 14170 5016 14172
rect 5040 14170 5096 14172
rect 5120 14170 5176 14172
rect 4880 14118 4926 14170
rect 4926 14118 4936 14170
rect 4960 14118 4990 14170
rect 4990 14118 5002 14170
rect 5002 14118 5016 14170
rect 5040 14118 5054 14170
rect 5054 14118 5066 14170
rect 5066 14118 5096 14170
rect 5120 14118 5130 14170
rect 5130 14118 5176 14170
rect 4880 14116 4936 14118
rect 4960 14116 5016 14118
rect 5040 14116 5096 14118
rect 5120 14116 5176 14118
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4880 13082 4936 13084
rect 4960 13082 5016 13084
rect 5040 13082 5096 13084
rect 5120 13082 5176 13084
rect 4880 13030 4926 13082
rect 4926 13030 4936 13082
rect 4960 13030 4990 13082
rect 4990 13030 5002 13082
rect 5002 13030 5016 13082
rect 5040 13030 5054 13082
rect 5054 13030 5066 13082
rect 5066 13030 5096 13082
rect 5120 13030 5130 13082
rect 5130 13030 5176 13082
rect 4880 13028 4936 13030
rect 4960 13028 5016 13030
rect 5040 13028 5096 13030
rect 5120 13028 5176 13030
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 3330 9580 3386 9616
rect 3330 9560 3332 9580
rect 3332 9560 3384 9580
rect 3384 9560 3386 9580
rect 3238 8492 3294 8528
rect 3238 8472 3240 8492
rect 3240 8472 3292 8492
rect 3292 8472 3294 8492
rect 2870 7928 2926 7984
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4158 10104 4214 10160
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 3422 7928 3478 7984
rect 3606 8608 3662 8664
rect 3606 8472 3662 8528
rect 4158 8492 4214 8528
rect 4158 8472 4160 8492
rect 4160 8472 4212 8492
rect 4212 8472 4214 8492
rect 4434 8472 4490 8528
rect 3882 7928 3938 7984
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4250 7248 4306 7304
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 11058 21936 11114 21992
rect 11702 24112 11758 24168
rect 11886 22752 11942 22808
rect 12162 21936 12218 21992
rect 12162 21548 12218 21584
rect 12162 21528 12164 21548
rect 12164 21528 12216 21548
rect 12216 21528 12218 21548
rect 13358 24148 13360 24168
rect 13360 24148 13412 24168
rect 13412 24148 13414 24168
rect 12806 23704 12862 23760
rect 13358 24112 13414 24148
rect 13358 23740 13360 23760
rect 13360 23740 13412 23760
rect 13412 23740 13414 23760
rect 13358 23704 13414 23740
rect 12438 18808 12494 18864
rect 12714 18808 12770 18864
rect 14278 23432 14334 23488
rect 15934 24112 15990 24168
rect 15014 22752 15070 22808
rect 16118 24692 16120 24712
rect 16120 24692 16172 24712
rect 16172 24692 16174 24712
rect 16118 24656 16174 24692
rect 17406 23432 17462 23488
rect 18418 24792 18474 24848
rect 24858 25236 24860 25256
rect 24860 25236 24912 25256
rect 24912 25236 24914 25256
rect 24858 25200 24914 25236
rect 4710 9968 4766 10024
rect 4894 10104 4950 10160
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 5170 9580 5226 9616
rect 5170 9560 5172 9580
rect 5172 9560 5224 9580
rect 5224 9560 5226 9580
rect 4710 8608 4766 8664
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 5078 8472 5134 8528
rect 4710 8372 4712 8392
rect 4712 8372 4764 8392
rect 4764 8372 4766 8392
rect 4710 8336 4766 8372
rect 5170 7928 5226 7984
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 5722 8336 5778 8392
rect 5078 7248 5134 7304
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 12254 14340 12310 14376
rect 12254 14320 12256 14340
rect 12256 14320 12308 14340
rect 12308 14320 12310 14340
rect 13082 14356 13084 14376
rect 13084 14356 13136 14376
rect 13136 14356 13138 14376
rect 13082 14320 13138 14356
rect 19246 24112 19302 24168
rect 19798 22208 19854 22264
rect 21086 24656 21142 24712
rect 21270 24148 21272 24168
rect 21272 24148 21324 24168
rect 21324 24148 21326 24168
rect 21270 24112 21326 24148
rect 9862 6296 9918 6352
rect 20994 23432 21050 23488
rect 21730 24792 21786 24848
rect 20718 15408 20774 15464
rect 11886 6724 11942 6760
rect 11886 6704 11888 6724
rect 11888 6704 11940 6724
rect 11940 6704 11942 6724
rect 11702 6316 11758 6352
rect 11702 6296 11704 6316
rect 11704 6296 11756 6316
rect 11756 6296 11758 6316
rect 12622 6740 12624 6760
rect 12624 6740 12676 6760
rect 12676 6740 12678 6760
rect 12622 6704 12678 6740
rect 12898 6296 12954 6352
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 18510 12280 18566 12336
rect 22006 21528 22062 21584
rect 22374 21548 22430 21584
rect 22374 21528 22376 21548
rect 22376 21528 22428 21548
rect 22428 21528 22430 21548
rect 21454 15272 21510 15328
rect 20902 12180 20904 12200
rect 20904 12180 20956 12200
rect 20956 12180 20958 12200
rect 20902 12144 20958 12180
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 21086 12416 21142 12472
rect 21454 13096 21510 13152
rect 24490 15272 24546 15328
rect 22190 13504 22246 13560
rect 22098 13404 22100 13424
rect 22100 13404 22152 13424
rect 22152 13404 22154 13424
rect 22098 13368 22154 13404
rect 22098 13132 22100 13152
rect 22100 13132 22152 13152
rect 22152 13132 22154 13152
rect 22098 13096 22154 13132
rect 22006 12416 22062 12472
rect 22650 13252 22706 13288
rect 22650 13232 22652 13252
rect 22652 13232 22704 13252
rect 22704 13232 22706 13252
rect 22558 12960 22614 13016
rect 23202 13524 23258 13560
rect 23202 13504 23204 13524
rect 23204 13504 23256 13524
rect 23256 13504 23258 13524
rect 23202 13368 23258 13424
rect 23294 13268 23296 13288
rect 23296 13268 23348 13288
rect 23348 13268 23350 13288
rect 22926 13096 22982 13152
rect 21546 6452 21602 6488
rect 21546 6432 21548 6452
rect 21548 6432 21600 6452
rect 21600 6432 21602 6452
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 22834 12688 22890 12744
rect 23294 13232 23350 13268
rect 23202 12280 23258 12336
rect 23386 12144 23442 12200
rect 24766 12960 24822 13016
rect 24858 3476 24860 3496
rect 24860 3476 24912 3496
rect 24912 3476 24914 3496
rect 24858 3440 24914 3476
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
<< metal3 >>
rect 4870 26144 5186 26145
rect 4870 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5186 26144
rect 4870 26079 5186 26080
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 24853 25258 24919 25261
rect 25525 25258 26325 25288
rect 24853 25256 26325 25258
rect 24853 25200 24858 25256
rect 24914 25200 26325 25256
rect 24853 25198 26325 25200
rect 24853 25195 24919 25198
rect 25525 25168 26325 25198
rect 4870 25056 5186 25057
rect 4870 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5186 25056
rect 4870 24991 5186 24992
rect 18413 24850 18479 24853
rect 21725 24850 21791 24853
rect 18413 24848 21791 24850
rect 18413 24792 18418 24848
rect 18474 24792 21730 24848
rect 21786 24792 21791 24848
rect 18413 24790 21791 24792
rect 18413 24787 18479 24790
rect 21725 24787 21791 24790
rect 8201 24714 8267 24717
rect 9029 24714 9095 24717
rect 8201 24712 9095 24714
rect 8201 24656 8206 24712
rect 8262 24656 9034 24712
rect 9090 24656 9095 24712
rect 8201 24654 9095 24656
rect 8201 24651 8267 24654
rect 9029 24651 9095 24654
rect 16113 24714 16179 24717
rect 21081 24714 21147 24717
rect 16113 24712 21147 24714
rect 16113 24656 16118 24712
rect 16174 24656 21086 24712
rect 21142 24656 21147 24712
rect 16113 24654 21147 24656
rect 16113 24651 16179 24654
rect 21081 24651 21147 24654
rect 0 24578 800 24608
rect 0 24518 1042 24578
rect 0 24488 800 24518
rect 105 24306 171 24309
rect 982 24306 1042 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 7465 24442 7531 24445
rect 9397 24442 9463 24445
rect 7465 24440 9463 24442
rect 7465 24384 7470 24440
rect 7526 24384 9402 24440
rect 9458 24384 9463 24440
rect 7465 24382 9463 24384
rect 7465 24379 7531 24382
rect 9397 24379 9463 24382
rect 105 24304 1042 24306
rect 105 24248 110 24304
rect 166 24248 1042 24304
rect 105 24246 1042 24248
rect 105 24243 171 24246
rect 11697 24170 11763 24173
rect 13353 24170 13419 24173
rect 15929 24170 15995 24173
rect 11697 24168 15995 24170
rect 11697 24112 11702 24168
rect 11758 24112 13358 24168
rect 13414 24112 15934 24168
rect 15990 24112 15995 24168
rect 11697 24110 15995 24112
rect 11697 24107 11763 24110
rect 13353 24107 13419 24110
rect 15929 24107 15995 24110
rect 19241 24170 19307 24173
rect 21265 24170 21331 24173
rect 19241 24168 21331 24170
rect 19241 24112 19246 24168
rect 19302 24112 21270 24168
rect 21326 24112 21331 24168
rect 19241 24110 21331 24112
rect 19241 24107 19307 24110
rect 21265 24107 21331 24110
rect 4870 23968 5186 23969
rect 4870 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5186 23968
rect 4870 23903 5186 23904
rect 12801 23762 12867 23765
rect 13353 23762 13419 23765
rect 12801 23760 13419 23762
rect 12801 23704 12806 23760
rect 12862 23704 13358 23760
rect 13414 23704 13419 23760
rect 12801 23702 13419 23704
rect 12801 23699 12867 23702
rect 13353 23699 13419 23702
rect 14273 23490 14339 23493
rect 17401 23490 17467 23493
rect 20989 23490 21055 23493
rect 14273 23488 21055 23490
rect 14273 23432 14278 23488
rect 14334 23432 17406 23488
rect 17462 23432 20994 23488
rect 21050 23432 21055 23488
rect 14273 23430 21055 23432
rect 14273 23427 14339 23430
rect 17401 23427 17467 23430
rect 20989 23427 21055 23430
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 4870 22880 5186 22881
rect 4870 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5186 22880
rect 4870 22815 5186 22816
rect 11881 22810 11947 22813
rect 15009 22810 15075 22813
rect 11881 22808 15075 22810
rect 11881 22752 11886 22808
rect 11942 22752 15014 22808
rect 15070 22752 15075 22808
rect 11881 22750 15075 22752
rect 11881 22747 11947 22750
rect 15009 22747 15075 22750
rect 9765 22538 9831 22541
rect 10133 22538 10199 22541
rect 9765 22536 12450 22538
rect 9765 22480 9770 22536
rect 9826 22480 10138 22536
rect 10194 22480 12450 22536
rect 9765 22478 12450 22480
rect 9765 22475 9831 22478
rect 10133 22475 10199 22478
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 12390 22266 12450 22478
rect 19793 22266 19859 22269
rect 12390 22264 19859 22266
rect 12390 22208 19798 22264
rect 19854 22208 19859 22264
rect 12390 22206 19859 22208
rect 19793 22203 19859 22206
rect 8845 21994 8911 21997
rect 11053 21994 11119 21997
rect 12157 21994 12223 21997
rect 8845 21992 12223 21994
rect 8845 21936 8850 21992
rect 8906 21936 11058 21992
rect 11114 21936 12162 21992
rect 12218 21936 12223 21992
rect 8845 21934 12223 21936
rect 8845 21931 8911 21934
rect 11053 21931 11119 21934
rect 12157 21931 12223 21934
rect 4870 21792 5186 21793
rect 4870 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5186 21792
rect 4870 21727 5186 21728
rect 12157 21586 12223 21589
rect 22001 21586 22067 21589
rect 22369 21586 22435 21589
rect 12157 21584 22435 21586
rect 12157 21528 12162 21584
rect 12218 21528 22006 21584
rect 22062 21528 22374 21584
rect 22430 21528 22435 21584
rect 12157 21526 22435 21528
rect 12157 21523 12223 21526
rect 22001 21523 22067 21526
rect 22369 21523 22435 21526
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 4870 20704 5186 20705
rect 4870 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5186 20704
rect 4870 20639 5186 20640
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 4870 19616 5186 19617
rect 4870 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5186 19616
rect 4870 19551 5186 19552
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 12433 18866 12499 18869
rect 12709 18866 12775 18869
rect 12433 18864 12775 18866
rect 12433 18808 12438 18864
rect 12494 18808 12714 18864
rect 12770 18808 12775 18864
rect 12433 18806 12775 18808
rect 12433 18803 12499 18806
rect 12709 18803 12775 18806
rect 4870 18528 5186 18529
rect 4870 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5186 18528
rect 4870 18463 5186 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 4870 17440 5186 17441
rect 4870 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5186 17440
rect 4870 17375 5186 17376
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 4870 16352 5186 16353
rect 4870 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5186 16352
rect 4870 16287 5186 16288
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 20713 15466 20779 15469
rect 20713 15464 20914 15466
rect 20713 15408 20718 15464
rect 20774 15408 20914 15464
rect 20713 15406 20914 15408
rect 20713 15403 20779 15406
rect 20854 15330 20914 15406
rect 21449 15330 21515 15333
rect 21582 15330 21588 15332
rect 20854 15328 21588 15330
rect 20854 15272 21454 15328
rect 21510 15272 21588 15328
rect 20854 15270 21588 15272
rect 21449 15267 21515 15270
rect 21582 15268 21588 15270
rect 21652 15330 21658 15332
rect 24485 15330 24551 15333
rect 21652 15328 24551 15330
rect 21652 15272 24490 15328
rect 24546 15272 24551 15328
rect 21652 15270 24551 15272
rect 21652 15268 21658 15270
rect 24485 15267 24551 15270
rect 4870 15264 5186 15265
rect 4870 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5186 15264
rect 4870 15199 5186 15200
rect 0 15058 800 15088
rect 1393 15058 1459 15061
rect 0 15056 1459 15058
rect 0 15000 1398 15056
rect 1454 15000 1459 15056
rect 0 14998 1459 15000
rect 0 14968 800 14998
rect 1393 14995 1459 14998
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 0 14378 800 14408
rect 12249 14378 12315 14381
rect 13077 14378 13143 14381
rect 0 14288 858 14378
rect 12249 14376 13143 14378
rect 12249 14320 12254 14376
rect 12310 14320 13082 14376
rect 13138 14320 13143 14376
rect 12249 14318 13143 14320
rect 12249 14315 12315 14318
rect 13077 14315 13143 14318
rect 798 14245 858 14288
rect 798 14240 907 14245
rect 798 14184 846 14240
rect 902 14184 907 14240
rect 798 14182 907 14184
rect 841 14179 907 14182
rect 4870 14176 5186 14177
rect 4870 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5186 14176
rect 4870 14111 5186 14112
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 22185 13562 22251 13565
rect 23197 13562 23263 13565
rect 22185 13560 23263 13562
rect 22185 13504 22190 13560
rect 22246 13504 23202 13560
rect 23258 13504 23263 13560
rect 22185 13502 23263 13504
rect 22185 13499 22251 13502
rect 23197 13499 23263 13502
rect 22093 13426 22159 13429
rect 23197 13426 23263 13429
rect 22093 13424 23263 13426
rect 22093 13368 22098 13424
rect 22154 13368 23202 13424
rect 23258 13368 23263 13424
rect 22093 13366 23263 13368
rect 22093 13363 22159 13366
rect 23197 13363 23263 13366
rect 22645 13290 22711 13293
rect 23289 13290 23355 13293
rect 22645 13288 23355 13290
rect 22645 13232 22650 13288
rect 22706 13232 23294 13288
rect 23350 13232 23355 13288
rect 22645 13230 23355 13232
rect 22645 13227 22711 13230
rect 23289 13227 23355 13230
rect 21449 13154 21515 13157
rect 22093 13154 22159 13157
rect 22921 13154 22987 13157
rect 21449 13152 22987 13154
rect 21449 13096 21454 13152
rect 21510 13096 22098 13152
rect 22154 13096 22926 13152
rect 22982 13096 22987 13152
rect 21449 13094 22987 13096
rect 21449 13091 21515 13094
rect 22093 13091 22159 13094
rect 22921 13091 22987 13094
rect 4870 13088 5186 13089
rect 4870 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5186 13088
rect 4870 13023 5186 13024
rect 22553 13018 22619 13021
rect 24761 13018 24827 13021
rect 25525 13018 26325 13048
rect 22553 13016 22754 13018
rect 22553 12960 22558 13016
rect 22614 12960 22754 13016
rect 22553 12958 22754 12960
rect 22553 12955 22619 12958
rect 22694 12746 22754 12958
rect 24761 13016 26325 13018
rect 24761 12960 24766 13016
rect 24822 12960 26325 13016
rect 24761 12958 26325 12960
rect 24761 12955 24827 12958
rect 25525 12928 26325 12958
rect 22829 12746 22895 12749
rect 22694 12744 22895 12746
rect 22694 12688 22834 12744
rect 22890 12688 22895 12744
rect 22694 12686 22895 12688
rect 22829 12683 22895 12686
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 21081 12474 21147 12477
rect 22001 12474 22067 12477
rect 21081 12472 22067 12474
rect 21081 12416 21086 12472
rect 21142 12416 22006 12472
rect 22062 12416 22067 12472
rect 21081 12414 22067 12416
rect 21081 12411 21147 12414
rect 22001 12411 22067 12414
rect 18505 12338 18571 12341
rect 23197 12338 23263 12341
rect 18505 12336 23263 12338
rect 18505 12280 18510 12336
rect 18566 12280 23202 12336
rect 23258 12280 23263 12336
rect 18505 12278 23263 12280
rect 18505 12275 18571 12278
rect 23197 12275 23263 12278
rect 20897 12202 20963 12205
rect 23381 12202 23447 12205
rect 20897 12200 23447 12202
rect 20897 12144 20902 12200
rect 20958 12144 23386 12200
rect 23442 12144 23447 12200
rect 20897 12142 23447 12144
rect 20897 12139 20963 12142
rect 23381 12139 23447 12142
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 0 11658 800 11688
rect 0 11568 858 11658
rect 798 11525 858 11568
rect 798 11520 907 11525
rect 798 11464 846 11520
rect 902 11464 907 11520
rect 798 11462 907 11464
rect 841 11459 907 11462
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 4870 10847 5186 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 4153 10162 4219 10165
rect 4889 10162 4955 10165
rect 4153 10160 4955 10162
rect 4153 10104 4158 10160
rect 4214 10104 4894 10160
rect 4950 10104 4955 10160
rect 4153 10102 4955 10104
rect 4153 10099 4219 10102
rect 4889 10099 4955 10102
rect 4705 10026 4771 10029
rect 4662 10024 4771 10026
rect 4662 9968 4710 10024
rect 4766 9968 4771 10024
rect 4662 9963 4771 9968
rect 3325 9618 3391 9621
rect 4662 9618 4722 9963
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 5165 9618 5231 9621
rect 3325 9616 5231 9618
rect 3325 9560 3330 9616
rect 3386 9560 5170 9616
rect 5226 9560 5231 9616
rect 3325 9558 5231 9560
rect 3325 9555 3391 9558
rect 5165 9555 5231 9558
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 3601 8666 3667 8669
rect 4705 8666 4771 8669
rect 3601 8664 4771 8666
rect 3601 8608 3606 8664
rect 3662 8608 4710 8664
rect 4766 8608 4771 8664
rect 3601 8606 4771 8608
rect 3601 8603 3667 8606
rect 4705 8603 4771 8606
rect 3233 8530 3299 8533
rect 3601 8530 3667 8533
rect 4153 8530 4219 8533
rect 3233 8528 4219 8530
rect 3233 8472 3238 8528
rect 3294 8472 3606 8528
rect 3662 8472 4158 8528
rect 4214 8472 4219 8528
rect 3233 8470 4219 8472
rect 3233 8467 3299 8470
rect 3601 8467 3667 8470
rect 4153 8467 4219 8470
rect 4429 8530 4495 8533
rect 5073 8530 5139 8533
rect 4429 8528 5139 8530
rect 4429 8472 4434 8528
rect 4490 8472 5078 8528
rect 5134 8472 5139 8528
rect 4429 8470 5139 8472
rect 4429 8467 4495 8470
rect 5073 8467 5139 8470
rect 4705 8394 4771 8397
rect 5717 8394 5783 8397
rect 4705 8392 5783 8394
rect 4705 8336 4710 8392
rect 4766 8336 5722 8392
rect 5778 8336 5783 8392
rect 4705 8334 5783 8336
rect 4705 8331 4771 8334
rect 5717 8331 5783 8334
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 2865 7986 2931 7989
rect 3417 7986 3483 7989
rect 3877 7986 3943 7989
rect 5165 7986 5231 7989
rect 2865 7984 5231 7986
rect 2865 7928 2870 7984
rect 2926 7928 3422 7984
rect 3478 7928 3882 7984
rect 3938 7928 5170 7984
rect 5226 7928 5231 7984
rect 2865 7926 5231 7928
rect 2865 7923 2931 7926
rect 3417 7923 3483 7926
rect 3877 7923 3943 7926
rect 5165 7923 5231 7926
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 4245 7306 4311 7309
rect 5073 7306 5139 7309
rect 4245 7304 5139 7306
rect 4245 7248 4250 7304
rect 4306 7248 5078 7304
rect 5134 7248 5139 7304
rect 4245 7246 5139 7248
rect 4245 7243 4311 7246
rect 5073 7243 5139 7246
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 11881 6762 11947 6765
rect 12617 6762 12683 6765
rect 11881 6760 12683 6762
rect 11881 6704 11886 6760
rect 11942 6704 12622 6760
rect 12678 6704 12683 6760
rect 11881 6702 12683 6704
rect 11881 6699 11947 6702
rect 12617 6699 12683 6702
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 21541 6492 21607 6493
rect 21541 6490 21588 6492
rect 21496 6488 21588 6490
rect 21496 6432 21546 6488
rect 21496 6430 21588 6432
rect 21541 6428 21588 6430
rect 21652 6428 21658 6492
rect 21541 6427 21607 6428
rect 9857 6354 9923 6357
rect 11697 6354 11763 6357
rect 12893 6354 12959 6357
rect 9857 6352 12959 6354
rect 9857 6296 9862 6352
rect 9918 6296 11702 6352
rect 11758 6296 12898 6352
rect 12954 6296 12959 6352
rect 9857 6294 12959 6296
rect 9857 6291 9923 6294
rect 11697 6291 11763 6294
rect 12893 6291 12959 6294
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 4870 5407 5186 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 24853 3498 24919 3501
rect 25525 3498 26325 3528
rect 24853 3496 26325 3498
rect 24853 3440 24858 3496
rect 24914 3440 26325 3496
rect 24853 3438 26325 3440
rect 24853 3435 24919 3438
rect 25525 3408 26325 3438
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
<< via3 >>
rect 4876 26140 4940 26144
rect 4876 26084 4880 26140
rect 4880 26084 4936 26140
rect 4936 26084 4940 26140
rect 4876 26080 4940 26084
rect 4956 26140 5020 26144
rect 4956 26084 4960 26140
rect 4960 26084 5016 26140
rect 5016 26084 5020 26140
rect 4956 26080 5020 26084
rect 5036 26140 5100 26144
rect 5036 26084 5040 26140
rect 5040 26084 5096 26140
rect 5096 26084 5100 26140
rect 5036 26080 5100 26084
rect 5116 26140 5180 26144
rect 5116 26084 5120 26140
rect 5120 26084 5176 26140
rect 5176 26084 5180 26140
rect 5116 26080 5180 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 4876 25052 4940 25056
rect 4876 24996 4880 25052
rect 4880 24996 4936 25052
rect 4936 24996 4940 25052
rect 4876 24992 4940 24996
rect 4956 25052 5020 25056
rect 4956 24996 4960 25052
rect 4960 24996 5016 25052
rect 5016 24996 5020 25052
rect 4956 24992 5020 24996
rect 5036 25052 5100 25056
rect 5036 24996 5040 25052
rect 5040 24996 5096 25052
rect 5096 24996 5100 25052
rect 5036 24992 5100 24996
rect 5116 25052 5180 25056
rect 5116 24996 5120 25052
rect 5120 24996 5176 25052
rect 5176 24996 5180 25052
rect 5116 24992 5180 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 4876 23964 4940 23968
rect 4876 23908 4880 23964
rect 4880 23908 4936 23964
rect 4936 23908 4940 23964
rect 4876 23904 4940 23908
rect 4956 23964 5020 23968
rect 4956 23908 4960 23964
rect 4960 23908 5016 23964
rect 5016 23908 5020 23964
rect 4956 23904 5020 23908
rect 5036 23964 5100 23968
rect 5036 23908 5040 23964
rect 5040 23908 5096 23964
rect 5096 23908 5100 23964
rect 5036 23904 5100 23908
rect 5116 23964 5180 23968
rect 5116 23908 5120 23964
rect 5120 23908 5176 23964
rect 5176 23908 5180 23964
rect 5116 23904 5180 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 4876 22876 4940 22880
rect 4876 22820 4880 22876
rect 4880 22820 4936 22876
rect 4936 22820 4940 22876
rect 4876 22816 4940 22820
rect 4956 22876 5020 22880
rect 4956 22820 4960 22876
rect 4960 22820 5016 22876
rect 5016 22820 5020 22876
rect 4956 22816 5020 22820
rect 5036 22876 5100 22880
rect 5036 22820 5040 22876
rect 5040 22820 5096 22876
rect 5096 22820 5100 22876
rect 5036 22816 5100 22820
rect 5116 22876 5180 22880
rect 5116 22820 5120 22876
rect 5120 22820 5176 22876
rect 5176 22820 5180 22876
rect 5116 22816 5180 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 4876 21788 4940 21792
rect 4876 21732 4880 21788
rect 4880 21732 4936 21788
rect 4936 21732 4940 21788
rect 4876 21728 4940 21732
rect 4956 21788 5020 21792
rect 4956 21732 4960 21788
rect 4960 21732 5016 21788
rect 5016 21732 5020 21788
rect 4956 21728 5020 21732
rect 5036 21788 5100 21792
rect 5036 21732 5040 21788
rect 5040 21732 5096 21788
rect 5096 21732 5100 21788
rect 5036 21728 5100 21732
rect 5116 21788 5180 21792
rect 5116 21732 5120 21788
rect 5120 21732 5176 21788
rect 5176 21732 5180 21788
rect 5116 21728 5180 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 4876 20700 4940 20704
rect 4876 20644 4880 20700
rect 4880 20644 4936 20700
rect 4936 20644 4940 20700
rect 4876 20640 4940 20644
rect 4956 20700 5020 20704
rect 4956 20644 4960 20700
rect 4960 20644 5016 20700
rect 5016 20644 5020 20700
rect 4956 20640 5020 20644
rect 5036 20700 5100 20704
rect 5036 20644 5040 20700
rect 5040 20644 5096 20700
rect 5096 20644 5100 20700
rect 5036 20640 5100 20644
rect 5116 20700 5180 20704
rect 5116 20644 5120 20700
rect 5120 20644 5176 20700
rect 5176 20644 5180 20700
rect 5116 20640 5180 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 4876 19612 4940 19616
rect 4876 19556 4880 19612
rect 4880 19556 4936 19612
rect 4936 19556 4940 19612
rect 4876 19552 4940 19556
rect 4956 19612 5020 19616
rect 4956 19556 4960 19612
rect 4960 19556 5016 19612
rect 5016 19556 5020 19612
rect 4956 19552 5020 19556
rect 5036 19612 5100 19616
rect 5036 19556 5040 19612
rect 5040 19556 5096 19612
rect 5096 19556 5100 19612
rect 5036 19552 5100 19556
rect 5116 19612 5180 19616
rect 5116 19556 5120 19612
rect 5120 19556 5176 19612
rect 5176 19556 5180 19612
rect 5116 19552 5180 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 4876 18524 4940 18528
rect 4876 18468 4880 18524
rect 4880 18468 4936 18524
rect 4936 18468 4940 18524
rect 4876 18464 4940 18468
rect 4956 18524 5020 18528
rect 4956 18468 4960 18524
rect 4960 18468 5016 18524
rect 5016 18468 5020 18524
rect 4956 18464 5020 18468
rect 5036 18524 5100 18528
rect 5036 18468 5040 18524
rect 5040 18468 5096 18524
rect 5096 18468 5100 18524
rect 5036 18464 5100 18468
rect 5116 18524 5180 18528
rect 5116 18468 5120 18524
rect 5120 18468 5176 18524
rect 5176 18468 5180 18524
rect 5116 18464 5180 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 4876 17436 4940 17440
rect 4876 17380 4880 17436
rect 4880 17380 4936 17436
rect 4936 17380 4940 17436
rect 4876 17376 4940 17380
rect 4956 17436 5020 17440
rect 4956 17380 4960 17436
rect 4960 17380 5016 17436
rect 5016 17380 5020 17436
rect 4956 17376 5020 17380
rect 5036 17436 5100 17440
rect 5036 17380 5040 17436
rect 5040 17380 5096 17436
rect 5096 17380 5100 17436
rect 5036 17376 5100 17380
rect 5116 17436 5180 17440
rect 5116 17380 5120 17436
rect 5120 17380 5176 17436
rect 5176 17380 5180 17436
rect 5116 17376 5180 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 4876 16348 4940 16352
rect 4876 16292 4880 16348
rect 4880 16292 4936 16348
rect 4936 16292 4940 16348
rect 4876 16288 4940 16292
rect 4956 16348 5020 16352
rect 4956 16292 4960 16348
rect 4960 16292 5016 16348
rect 5016 16292 5020 16348
rect 4956 16288 5020 16292
rect 5036 16348 5100 16352
rect 5036 16292 5040 16348
rect 5040 16292 5096 16348
rect 5096 16292 5100 16348
rect 5036 16288 5100 16292
rect 5116 16348 5180 16352
rect 5116 16292 5120 16348
rect 5120 16292 5176 16348
rect 5176 16292 5180 16348
rect 5116 16288 5180 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 21588 15268 21652 15332
rect 4876 15260 4940 15264
rect 4876 15204 4880 15260
rect 4880 15204 4936 15260
rect 4936 15204 4940 15260
rect 4876 15200 4940 15204
rect 4956 15260 5020 15264
rect 4956 15204 4960 15260
rect 4960 15204 5016 15260
rect 5016 15204 5020 15260
rect 4956 15200 5020 15204
rect 5036 15260 5100 15264
rect 5036 15204 5040 15260
rect 5040 15204 5096 15260
rect 5096 15204 5100 15260
rect 5036 15200 5100 15204
rect 5116 15260 5180 15264
rect 5116 15204 5120 15260
rect 5120 15204 5176 15260
rect 5176 15204 5180 15260
rect 5116 15200 5180 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 4876 14172 4940 14176
rect 4876 14116 4880 14172
rect 4880 14116 4936 14172
rect 4936 14116 4940 14172
rect 4876 14112 4940 14116
rect 4956 14172 5020 14176
rect 4956 14116 4960 14172
rect 4960 14116 5016 14172
rect 5016 14116 5020 14172
rect 4956 14112 5020 14116
rect 5036 14172 5100 14176
rect 5036 14116 5040 14172
rect 5040 14116 5096 14172
rect 5096 14116 5100 14172
rect 5036 14112 5100 14116
rect 5116 14172 5180 14176
rect 5116 14116 5120 14172
rect 5120 14116 5176 14172
rect 5176 14116 5180 14172
rect 5116 14112 5180 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 4876 13084 4940 13088
rect 4876 13028 4880 13084
rect 4880 13028 4936 13084
rect 4936 13028 4940 13084
rect 4876 13024 4940 13028
rect 4956 13084 5020 13088
rect 4956 13028 4960 13084
rect 4960 13028 5016 13084
rect 5016 13028 5020 13084
rect 4956 13024 5020 13028
rect 5036 13084 5100 13088
rect 5036 13028 5040 13084
rect 5040 13028 5096 13084
rect 5096 13028 5100 13084
rect 5036 13024 5100 13028
rect 5116 13084 5180 13088
rect 5116 13028 5120 13084
rect 5120 13028 5176 13084
rect 5176 13028 5180 13084
rect 5116 13024 5180 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 21588 6488 21652 6492
rect 21588 6432 21602 6488
rect 21602 6432 21652 6488
rect 21588 6428 21652 6432
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
<< metal4 >>
rect 4208 25600 4528 26160
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 26144 5188 26160
rect 4868 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5188 26144
rect 4868 25056 5188 26080
rect 4868 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5188 25056
rect 4868 23968 5188 24992
rect 4868 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5188 23968
rect 4868 22880 5188 23904
rect 4868 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5188 22880
rect 4868 21792 5188 22816
rect 4868 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5188 21792
rect 4868 20704 5188 21728
rect 4868 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5188 20704
rect 4868 19616 5188 20640
rect 4868 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5188 19616
rect 4868 18528 5188 19552
rect 4868 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5188 18528
rect 4868 17440 5188 18464
rect 4868 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5188 17440
rect 4868 16352 5188 17376
rect 4868 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5188 16352
rect 4868 15264 5188 16288
rect 21587 15332 21653 15333
rect 21587 15268 21588 15332
rect 21652 15268 21653 15332
rect 21587 15267 21653 15268
rect 4868 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5188 15264
rect 4868 14176 5188 15200
rect 4868 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5188 14176
rect 4868 13088 5188 14112
rect 4868 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5188 13088
rect 4868 12000 5188 13024
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4868 10912 5188 11936
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 5472 5188 6496
rect 21590 6493 21650 15267
rect 21587 6492 21653 6493
rect 21587 6428 21588 6492
rect 21652 6428 21653 6492
rect 21587 6427 21653 6428
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
use sky130_fd_sc_hd__inv_2  _0442_
timestamp 1
transform -1 0 5980 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0443_
timestamp 1
transform 1 0 5612 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0444_
timestamp 1
transform -1 0 15180 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0445_
timestamp 1
transform -1 0 11132 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0446_
timestamp 1
transform 1 0 13156 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0447_
timestamp 1
transform -1 0 10488 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0448_
timestamp 1
transform 1 0 15456 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0449_
timestamp 1
transform 1 0 16652 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0450_
timestamp 1
transform 1 0 16928 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0451_
timestamp 1
transform 1 0 15916 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0452_
timestamp 1
transform -1 0 17480 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0453_
timestamp 1
transform 1 0 4324 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0454_
timestamp 1
transform 1 0 4876 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or4bb_1  _0455_
timestamp 1
transform 1 0 3772 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _0456_
timestamp 1
transform 1 0 5336 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a211oi_1  _0457_
timestamp 1
transform -1 0 5152 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _0458_
timestamp 1
transform 1 0 3404 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0459_
timestamp 1
transform 1 0 3404 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0460_
timestamp 1
transform 1 0 2852 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_2  _0461_
timestamp 1
transform -1 0 3404 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0462_
timestamp 1
transform -1 0 4876 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0463_
timestamp 1
transform -1 0 5336 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0464_
timestamp 1
transform -1 0 5428 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _0465_
timestamp 1
transform -1 0 5980 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0466_
timestamp 1
transform -1 0 3680 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0467_
timestamp 1
transform 1 0 3404 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _0468_
timestamp 1
transform -1 0 5796 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0469_
timestamp 1
transform -1 0 4968 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0470_
timestamp 1
transform -1 0 7636 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0471_
timestamp 1
transform -1 0 4692 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0472_
timestamp 1
transform -1 0 3496 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0473_
timestamp 1
transform 1 0 4784 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0474_
timestamp 1
transform 1 0 1932 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0475_
timestamp 1
transform -1 0 4784 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0476_
timestamp 1
transform 1 0 3772 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0477_
timestamp 1
transform 1 0 8280 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _0478_
timestamp 1
transform -1 0 12788 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0479_
timestamp 1
transform 1 0 10488 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0480_
timestamp 1
transform 1 0 7728 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _0481_
timestamp 1
transform 1 0 8372 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _0482_
timestamp 1
transform -1 0 13432 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _0483_
timestamp 1
transform 1 0 12328 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _0484_
timestamp 1
transform -1 0 11776 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _0485_
timestamp 1
transform 1 0 11040 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0486_
timestamp 1
transform 1 0 7820 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0487_
timestamp 1
transform 1 0 8372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0488_
timestamp 1
transform 1 0 10580 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0489_
timestamp 1
transform -1 0 9568 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _0490_
timestamp 1
transform 1 0 12052 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0491_
timestamp 1
transform 1 0 9568 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0492_
timestamp 1
transform 1 0 11500 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__a221oi_1  _0493_
timestamp 1
transform 1 0 11408 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0494_
timestamp 1
transform -1 0 12604 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o2111a_1  _0495_
timestamp 1
transform 1 0 11500 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__a2111oi_1  _0496_
timestamp 1
transform 1 0 10672 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a2111oi_1  _0497_
timestamp 1
transform -1 0 9384 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _0498_
timestamp 1
transform 1 0 9384 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _0499_
timestamp 1
transform -1 0 10488 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0500_
timestamp 1
transform -1 0 6808 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor3b_2  _0501_
timestamp 1
transform 1 0 3772 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__and4bb_1  _0502_
timestamp 1
transform 1 0 4232 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _0503_
timestamp 1
transform 1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _0504_
timestamp 1
transform 1 0 5428 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a31oi_2  _0505_
timestamp 1
transform 1 0 5612 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0506_
timestamp 1
transform 1 0 8096 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0507_
timestamp 1
transform 1 0 7636 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0508_
timestamp 1
transform 1 0 8556 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0509_
timestamp 1
transform -1 0 7636 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0510_
timestamp 1
transform 1 0 8280 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0511_
timestamp 1
transform 1 0 9200 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0512_
timestamp 1
transform -1 0 8004 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0513_
timestamp 1
transform 1 0 6900 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0514_
timestamp 1
transform 1 0 7360 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0515_
timestamp 1
transform -1 0 9384 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0516_
timestamp 1
transform -1 0 7084 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0517_
timestamp 1
transform -1 0 6256 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0518_
timestamp 1
transform -1 0 8464 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0519_
timestamp 1
transform -1 0 7728 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0520_
timestamp 1
transform -1 0 7728 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0521_
timestamp 1
transform 1 0 8188 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0522_
timestamp 1
transform 1 0 8372 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0523_
timestamp 1
transform 1 0 9568 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0524_
timestamp 1
transform -1 0 13616 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0525_
timestamp 1
transform 1 0 13432 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0526_
timestamp 1
transform 1 0 12420 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0527_
timestamp 1
transform -1 0 13156 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0528_
timestamp 1
transform 1 0 13708 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _0529_
timestamp 1
transform -1 0 12328 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0530_
timestamp 1
transform -1 0 11408 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0531_
timestamp 1
transform 1 0 11868 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0532_
timestamp 1
transform 1 0 12052 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0533_
timestamp 1
transform -1 0 13156 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0534_
timestamp 1
transform -1 0 12144 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0535_
timestamp 1
transform 1 0 12512 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0536_
timestamp 1
transform 1 0 13248 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0537_
timestamp 1
transform 1 0 13708 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0538_
timestamp 1
transform 1 0 12880 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0539_
timestamp 1
transform -1 0 13156 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0540_
timestamp 1
transform -1 0 12696 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0541_
timestamp 1
transform -1 0 15272 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0542_
timestamp 1
transform -1 0 13064 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0543_
timestamp 1
transform -1 0 13524 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0544_
timestamp 1
transform -1 0 14628 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _0545_
timestamp 1
transform -1 0 14168 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0546_
timestamp 1
transform -1 0 13892 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0547_
timestamp 1
transform 1 0 9660 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0548_
timestamp 1
transform 1 0 7360 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0549_
timestamp 1
transform 1 0 9108 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0550_
timestamp 1
transform 1 0 7636 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0551_
timestamp 1
transform 1 0 6716 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0552_
timestamp 1
transform 1 0 13064 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0553_
timestamp 1
transform 1 0 12604 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0554_
timestamp 1
transform -1 0 10488 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0555_
timestamp 1
transform -1 0 9568 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0556_
timestamp 1
transform 1 0 9476 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _0557_
timestamp 1
transform 1 0 10028 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _0558_
timestamp 1
transform 1 0 9384 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0559_
timestamp 1
transform 1 0 8280 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0560_
timestamp 1
transform 1 0 13064 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0561_
timestamp 1
transform 1 0 13156 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0562_
timestamp 1
transform -1 0 11316 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0563_
timestamp 1
transform 1 0 12420 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0564_
timestamp 1
transform 1 0 13064 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0565_
timestamp 1
transform 1 0 10212 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and4bb_1  _0566_
timestamp 1
transform 1 0 1932 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__nand2b_1  _0567_
timestamp 1
transform -1 0 3312 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _0568_
timestamp 1
transform 1 0 4232 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0569_
timestamp 1
transform -1 0 4416 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0570_
timestamp 1
transform -1 0 23000 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0571_
timestamp 1
transform 1 0 20976 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0572_
timestamp 1
transform 1 0 19320 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0573_
timestamp 1
transform 1 0 16468 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0574_
timestamp 1
transform -1 0 20424 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0575_
timestamp 1
transform 1 0 16928 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0576_
timestamp 1
transform 1 0 17756 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0577_
timestamp 1
transform -1 0 17204 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _0578_
timestamp 1
transform 1 0 21068 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0579_
timestamp 1
transform -1 0 18400 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _0580_
timestamp 1
transform 1 0 15180 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0581_
timestamp 1
transform -1 0 21620 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0582_
timestamp 1
transform 1 0 16008 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0583_
timestamp 1
transform -1 0 21344 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0584_
timestamp 1
transform -1 0 15732 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _0585_
timestamp 1
transform 1 0 21804 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _0586_
timestamp 1
transform 1 0 19964 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0587_
timestamp 1
transform 1 0 16560 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0588_
timestamp 1
transform -1 0 21712 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0589_
timestamp 1
transform 1 0 17848 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _0590_
timestamp 1
transform -1 0 17664 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0591_
timestamp 1
transform -1 0 19780 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _0592_
timestamp 1
transform 1 0 16100 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0593_
timestamp 1
transform 1 0 15088 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a2111o_1  _0594_
timestamp 1
transform 1 0 20516 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__o2111ai_1  _0595_
timestamp 1
transform 1 0 21804 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o2111a_1  _0596_
timestamp 1
transform -1 0 17480 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _0597_
timestamp 1
transform -1 0 20424 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _0598_
timestamp 1
transform 1 0 17940 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__a2111o_1  _0599_
timestamp 1
transform 1 0 17020 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__a2111o_1  _0600_
timestamp 1
transform 1 0 17664 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__a2111o_1  _0601_
timestamp 1
transform 1 0 15732 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _0602_
timestamp 1
transform 1 0 17112 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0603_
timestamp 1
transform -1 0 19136 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0604_
timestamp 1
transform 1 0 18584 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _0605_
timestamp 1
transform -1 0 19964 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0606_
timestamp 1
transform -1 0 16468 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0607_
timestamp 1
transform 1 0 17296 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0608_
timestamp 1
transform -1 0 16100 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0609_
timestamp 1
transform 1 0 15640 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0610_
timestamp 1
transform 1 0 14996 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0611_
timestamp 1
transform 1 0 15456 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0612_
timestamp 1
transform 1 0 16652 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0613_
timestamp 1
transform 1 0 16744 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0614_
timestamp 1
transform -1 0 17296 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0615_
timestamp 1
transform -1 0 19136 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0616_
timestamp 1
transform 1 0 18400 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0617_
timestamp 1
transform -1 0 19136 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0618_
timestamp 1
transform 1 0 20056 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0619_
timestamp 1
transform -1 0 21160 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0620_
timestamp 1
transform 1 0 20516 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0621_
timestamp 1
transform 1 0 21160 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0622_
timestamp 1
transform 1 0 21252 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0623_
timestamp 1
transform -1 0 22448 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0624_
timestamp 1
transform 1 0 23460 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0625_
timestamp 1
transform 1 0 22724 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0626_
timestamp 1
transform 1 0 22632 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0627_
timestamp 1
transform -1 0 22724 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0628_
timestamp 1
transform 1 0 21988 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0629_
timestamp 1
transform -1 0 22724 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0630_
timestamp 1
transform 1 0 22724 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0631_
timestamp 1
transform -1 0 22724 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0632_
timestamp 1
transform -1 0 22264 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0633_
timestamp 1
transform -1 0 21528 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0634_
timestamp 1
transform -1 0 21160 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0635_
timestamp 1
transform -1 0 20516 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0636_
timestamp 1
transform -1 0 20884 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0637_
timestamp 1
transform -1 0 20148 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0638_
timestamp 1
transform 1 0 19136 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0639_
timestamp 1
transform -1 0 19136 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0640_
timestamp 1
transform -1 0 20516 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0641_
timestamp 1
transform -1 0 18676 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0642_
timestamp 1
transform 1 0 17572 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0643_
timestamp 1
transform 1 0 16652 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0644_
timestamp 1
transform -1 0 15824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0645_
timestamp 1
transform -1 0 22448 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0646_
timestamp 1
transform -1 0 22724 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0647_
timestamp 1
transform 1 0 16100 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0648_
timestamp 1
transform 1 0 17296 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0649_
timestamp 1
transform 1 0 18032 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0650_
timestamp 1
transform -1 0 22448 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0651_
timestamp 1
transform 1 0 19228 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0652_
timestamp 1
transform -1 0 21068 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0653_
timestamp 1
transform 1 0 19412 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0654_
timestamp 1
transform 1 0 15364 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0655_
timestamp 1
transform 1 0 17848 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0656_
timestamp 1
transform 1 0 20056 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0657_
timestamp 1
transform -1 0 19964 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a211oi_1  _0658_
timestamp 1
transform 1 0 19136 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0659_
timestamp 1
transform 1 0 18032 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0660_
timestamp 1
transform 1 0 15824 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0661_
timestamp 1
transform 1 0 17204 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _0662_
timestamp 1
transform 1 0 17204 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__o2111a_1  _0663_
timestamp 1
transform -1 0 20056 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0664_
timestamp 1
transform -1 0 22356 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0665_
timestamp 1
transform -1 0 21712 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0666_
timestamp 1
transform -1 0 22448 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0667_
timestamp 1
transform 1 0 21712 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0668_
timestamp 1
transform -1 0 20148 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0669_
timestamp 1
transform -1 0 20700 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0670_
timestamp 1
transform 1 0 20332 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0671_
timestamp 1
transform 1 0 19504 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0672_
timestamp 1
transform -1 0 19872 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0673_
timestamp 1
transform -1 0 19504 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0674_
timestamp 1
transform 1 0 17572 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0675_
timestamp 1
transform 1 0 16652 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0676_
timestamp 1
transform 1 0 17296 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0677_
timestamp 1
transform 1 0 16928 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0678_
timestamp 1
transform 1 0 17204 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0679_
timestamp 1
transform -1 0 18768 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0680_
timestamp 1
transform -1 0 18216 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0681_
timestamp 1
transform 1 0 18676 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0682_
timestamp 1
transform -1 0 18676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _0683_
timestamp 1
transform -1 0 19136 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0684_
timestamp 1
transform -1 0 20424 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0685_
timestamp 1
transform 1 0 20332 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0686_
timestamp 1
transform 1 0 19872 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _0687_
timestamp 1
transform -1 0 21436 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _0688_
timestamp 1
transform 1 0 19228 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0689_
timestamp 1
transform -1 0 24196 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0690_
timestamp 1
transform 1 0 24288 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0691_
timestamp 1
transform -1 0 24288 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0692_
timestamp 1
transform -1 0 22908 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0693_
timestamp 1
transform -1 0 24012 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _0694_
timestamp 1
transform 1 0 21436 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0695_
timestamp 1
transform 1 0 20792 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0696_
timestamp 1
transform -1 0 22724 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor3b_1  _0697_
timestamp 1
transform 1 0 23092 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0698_
timestamp 1
transform 1 0 19136 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0699_
timestamp 1
transform -1 0 20240 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _0700_
timestamp 1
transform 1 0 21896 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0701_
timestamp 1
transform -1 0 23092 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0702_
timestamp 1
transform 1 0 23184 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0703_
timestamp 1
transform 1 0 22448 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0704_
timestamp 1
transform 1 0 21252 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0705_
timestamp 1
transform 1 0 21804 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0706_
timestamp 1
transform -1 0 20976 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0707_
timestamp 1
transform -1 0 21804 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0708_
timestamp 1
transform 1 0 20424 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _0709_
timestamp 1
transform 1 0 19964 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0710_
timestamp 1
transform 1 0 23644 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0711_
timestamp 1
transform -1 0 23184 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0712_
timestamp 1
transform -1 0 21344 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0713_
timestamp 1
transform -1 0 22448 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0714_
timestamp 1
transform -1 0 22816 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0715_
timestamp 1
transform -1 0 22356 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0716_
timestamp 1
transform 1 0 21988 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a2111oi_1  _0717_
timestamp 1
transform 1 0 22632 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0718_
timestamp 1
transform -1 0 18216 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0719_
timestamp 1
transform 1 0 18216 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0720_
timestamp 1
transform 1 0 18676 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _0721_
timestamp 1
transform 1 0 20976 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _0722_
timestamp 1
transform 1 0 17848 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0723_
timestamp 1
transform 1 0 18032 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0724_
timestamp 1
transform 1 0 20976 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0725_
timestamp 1
transform 1 0 19320 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0726_
timestamp 1
transform -1 0 20608 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0727_
timestamp 1
transform -1 0 21896 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0728_
timestamp 1
transform -1 0 22448 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0729_
timestamp 1
transform -1 0 6072 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _0730_
timestamp 1
transform -1 0 3680 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0731_
timestamp 1
transform -1 0 5888 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _0732_
timestamp 1
transform 1 0 2208 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_1  _0733_
timestamp 1
transform -1 0 3772 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__a211o_1  _0734_
timestamp 1
transform 1 0 2300 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0735_
timestamp 1
transform -1 0 5428 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0736_
timestamp 1
transform -1 0 3680 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0737_
timestamp 1
transform -1 0 23184 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0738_
timestamp 1
transform -1 0 22540 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0739_
timestamp 1
transform -1 0 20976 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0740_
timestamp 1
transform -1 0 20884 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _0741_
timestamp 1
transform 1 0 21344 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _0742_
timestamp 1
transform 1 0 23736 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a2111o_1  _0743_
timestamp 1
transform 1 0 21804 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0744_
timestamp 1
transform 1 0 20424 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0745_
timestamp 1
transform 1 0 22908 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_4  _0746_
timestamp 1
transform -1 0 5704 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _0747_
timestamp 1
transform 1 0 7636 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0748_
timestamp 1
transform 1 0 7636 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0749_
timestamp 1
transform 1 0 7176 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0750_
timestamp 1
transform 1 0 6348 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0751_
timestamp 1
transform 1 0 6348 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0752_
timestamp 1
transform 1 0 4784 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0753_
timestamp 1
transform -1 0 4232 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0754_
timestamp 1
transform 1 0 3772 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0755_
timestamp 1
transform 1 0 2116 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0756_
timestamp 1
transform 1 0 1748 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0757_
timestamp 1
transform -1 0 1656 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0758_
timestamp 1
transform -1 0 3680 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0759_
timestamp 1
transform 1 0 6900 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _0760_
timestamp 1
transform 1 0 5796 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0761_
timestamp 1
transform 1 0 6532 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0762_
timestamp 1
transform 1 0 12328 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0763_
timestamp 1
transform 1 0 16652 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__nand3_1  _0764_
timestamp 1
transform 1 0 12880 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0765_
timestamp 1
transform 1 0 12236 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0766_
timestamp 1
transform 1 0 13248 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0767_
timestamp 1
transform 1 0 17112 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0768_
timestamp 1
transform -1 0 13156 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0769_
timestamp 1
transform 1 0 11500 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22oi_1  _0770_
timestamp 1
transform -1 0 12696 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0771_
timestamp 1
transform 1 0 12328 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0772_
timestamp 1
transform 1 0 11684 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0773_
timestamp 1
transform -1 0 13892 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0774_
timestamp 1
transform -1 0 13524 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _0775_
timestamp 1
transform 1 0 14260 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0776_
timestamp 1
transform 1 0 11500 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0777_
timestamp 1
transform -1 0 10856 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0778_
timestamp 1
transform 1 0 10856 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0779_
timestamp 1
transform -1 0 12696 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0780_
timestamp 1
transform 1 0 11500 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0781_
timestamp 1
transform 1 0 12788 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _0782_
timestamp 1
transform 1 0 12972 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _0783_
timestamp 1
transform -1 0 12788 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0784_
timestamp 1
transform 1 0 12972 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0785_
timestamp 1
transform -1 0 12788 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0786_
timestamp 1
transform 1 0 13984 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0787_
timestamp 1
transform 1 0 15640 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0788_
timestamp 1
transform -1 0 16468 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0789_
timestamp 1
transform 1 0 16928 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0790_
timestamp 1
transform 1 0 12880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0791_
timestamp 1
transform 1 0 13156 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a22oi_1  _0792_
timestamp 1
transform 1 0 13800 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0793_
timestamp 1
transform 1 0 14076 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0794_
timestamp 1
transform 1 0 13892 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0795_
timestamp 1
transform -1 0 12144 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0796_
timestamp 1
transform 1 0 13248 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0797_
timestamp 1
transform 1 0 12696 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0798_
timestamp 1
transform 1 0 14720 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0799_
timestamp 1
transform 1 0 15364 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0800_
timestamp 1
transform 1 0 15824 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0801_
timestamp 1
transform -1 0 19136 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _0802_
timestamp 1
transform 1 0 14628 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_1  _0803_
timestamp 1
transform -1 0 13892 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0804_
timestamp 1
transform 1 0 14720 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0805_
timestamp 1
transform 1 0 14536 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _0806_
timestamp 1
transform 1 0 15640 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0807_
timestamp 1
transform 1 0 16376 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0808_
timestamp 1
transform 1 0 20516 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0809_
timestamp 1
transform 1 0 15732 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _0810_
timestamp 1
transform 1 0 15272 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0811_
timestamp 1
transform 1 0 15548 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0812_
timestamp 1
transform 1 0 15824 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a22oi_1  _0813_
timestamp 1
transform 1 0 17112 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0814_
timestamp 1
transform -1 0 3128 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0815_
timestamp 1
transform -1 0 3680 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0816_
timestamp 1
transform 1 0 4876 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0817_
timestamp 1
transform -1 0 4600 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _0818_
timestamp 1
transform 1 0 3588 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0819_
timestamp 1
transform 1 0 2760 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0820_
timestamp 1
transform 1 0 2484 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0821_
timestamp 1
transform 1 0 2852 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _0822_
timestamp 1
transform 1 0 2852 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _0823_
timestamp 1
transform -1 0 2852 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0824_
timestamp 1
transform 1 0 4600 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0825_
timestamp 1
transform -1 0 5336 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0826_
timestamp 1
transform -1 0 4876 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0827_
timestamp 1
transform 1 0 6992 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _0828_
timestamp 1
transform -1 0 6532 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0829_
timestamp 1
transform 1 0 4324 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0830_
timestamp 1
transform -1 0 5888 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0831_
timestamp 1
transform 1 0 5888 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0832_
timestamp 1
transform 1 0 6348 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0833_
timestamp 1
transform -1 0 4140 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _0834_
timestamp 1
transform 1 0 2852 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _0835_
timestamp 1
transform 1 0 4416 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0836_
timestamp 1
transform -1 0 4324 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0837_
timestamp 1
transform 1 0 3772 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0838_
timestamp 1
transform -1 0 3404 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0839_
timestamp 1
transform -1 0 4692 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_1  _0840_
timestamp 1
transform -1 0 4232 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0841_
timestamp 1
transform 1 0 3220 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__o311a_1  _0842_
timestamp 1
transform 1 0 6164 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o211ai_1  _0843_
timestamp 1
transform 1 0 5520 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0844_
timestamp 1
transform 1 0 6348 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0845_
timestamp 1
transform 1 0 3864 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0846_
timestamp 1
transform 1 0 2668 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _0847_
timestamp 1
transform -1 0 2852 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0848_
timestamp 1
transform 1 0 1932 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0849_
timestamp 1
transform 1 0 10028 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0850_
timestamp 1
transform -1 0 9752 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0851_
timestamp 1
transform 1 0 8924 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0852_
timestamp 1
transform 1 0 8004 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0853_
timestamp 1
transform 1 0 10028 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0854_
timestamp 1
transform 1 0 9108 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0855_
timestamp 1
transform 1 0 9752 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0856_
timestamp 1
transform 1 0 7728 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0857_
timestamp 1
transform 1 0 11500 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0858_
timestamp 1
transform 1 0 9568 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0859_
timestamp 1
transform 1 0 8556 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0860_
timestamp 1
transform 1 0 8004 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0861_
timestamp 1
transform 1 0 10396 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0862_
timestamp 1
transform 1 0 8924 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0863_
timestamp 1
transform 1 0 9752 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0864_
timestamp 1
transform 1 0 7176 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _0865_
timestamp 1
transform 1 0 14076 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0866_
timestamp 1
transform 1 0 16928 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nand4_1  _0867_
timestamp 1
transform 1 0 12880 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0868_
timestamp 1
transform 1 0 13064 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0869_
timestamp 1
transform 1 0 15272 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0870_
timestamp 1
transform 1 0 15548 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0871_
timestamp 1
transform -1 0 15272 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0872_
timestamp 1
transform 1 0 12236 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22oi_1  _0873_
timestamp 1
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0874_
timestamp 1
transform 1 0 13524 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0875_
timestamp 1
transform 1 0 13984 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0876_
timestamp 1
transform -1 0 15824 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0877_
timestamp 1
transform -1 0 15272 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _0878_
timestamp 1
transform 1 0 15732 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0879_
timestamp 1
transform -1 0 13064 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0880_
timestamp 1
transform 1 0 11500 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0881_
timestamp 1
transform 1 0 11500 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0882_
timestamp 1
transform 1 0 11684 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0883_
timestamp 1
transform 1 0 12144 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0884_
timestamp 1
transform -1 0 13892 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0885_
timestamp 1
transform 1 0 14076 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0886_
timestamp 1
transform -1 0 15732 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _0887_
timestamp 1
transform -1 0 14812 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0888_
timestamp 1
transform 1 0 14812 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0889_
timestamp 1
transform 1 0 15456 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0890_
timestamp 1
transform 1 0 17296 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0891_
timestamp 1
transform 1 0 12052 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0892_
timestamp 1
transform 1 0 11132 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22oi_1  _0893_
timestamp 1
transform 1 0 11592 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0894_
timestamp 1
transform 1 0 12144 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0895_
timestamp 1
transform 1 0 11960 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0896_
timestamp 1
transform -1 0 12420 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0897_
timestamp 1
transform 1 0 14720 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0898_
timestamp 1
transform 1 0 12420 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0899_
timestamp 1
transform -1 0 13432 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0900_
timestamp 1
transform 1 0 13340 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0901_
timestamp 1
transform 1 0 13708 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0902_
timestamp 1
transform 1 0 18032 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _0903_
timestamp 1
transform 1 0 12696 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0904_
timestamp 1
transform -1 0 13984 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _0905_
timestamp 1
transform -1 0 13432 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o21bai_1  _0906_
timestamp 1
transform -1 0 13156 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0907_
timestamp 1
transform 1 0 12420 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0908_
timestamp 1
transform 1 0 13340 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0909_
timestamp 1
transform 1 0 17020 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0910_
timestamp 1
transform 1 0 13432 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _0911_
timestamp 1
transform 1 0 14076 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0912_
timestamp 1
transform -1 0 13340 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0913_
timestamp 1
transform 1 0 14076 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _0914_
timestamp 1
transform 1 0 15456 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0915_
timestamp 1
transform 1 0 6348 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0916_
timestamp 1
transform 1 0 5428 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0917_
timestamp 1
transform 1 0 6348 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0918_
timestamp 1
transform 1 0 6900 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0919_
timestamp 1
transform 1 0 4140 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0920_
timestamp 1
transform 1 0 2760 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0921_
timestamp 1
transform 1 0 2392 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0922_
timestamp 1
transform 1 0 2392 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0923_
timestamp 1
transform 1 0 1840 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_1  _0924_
timestamp 1
transform 1 0 20884 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0925_
timestamp 1
transform -1 0 24932 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0926_
timestamp 1
transform 1 0 19228 0 -1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0927_
timestamp 1
transform 1 0 22448 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0928_
timestamp 1
transform 1 0 22816 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _0929_
timestamp 1
transform 1 0 7452 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _0930_
timestamp 1
transform 1 0 7452 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _0931_
timestamp 1
transform 1 0 6808 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _0932_
timestamp 1
transform 1 0 4968 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _0933_
timestamp 1
transform 1 0 6348 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _0934_
timestamp 1
transform 1 0 4324 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _0935_
timestamp 1
transform 1 0 3772 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _0936_
timestamp 1
transform 1 0 3220 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _0937_
timestamp 1
transform 1 0 1380 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _0938_
timestamp 1
transform -1 0 5796 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _0939_
timestamp 1
transform -1 0 4600 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0940_
timestamp 1
transform 1 0 1380 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0941_
timestamp 1
transform 1 0 1656 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _0942_
timestamp 1
transform 1 0 16100 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _0943_
timestamp 1
transform 1 0 15180 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _0944_
timestamp 1
transform 1 0 14260 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _0945_
timestamp 1
transform 1 0 17848 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _0946_
timestamp 1
transform -1 0 21160 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _0947_
timestamp 1
transform 1 0 19228 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _0948_
timestamp 1
transform 1 0 16652 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _0949_
timestamp 1
transform -1 0 20516 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0950_
timestamp 1
transform 1 0 1380 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0951_
timestamp 1
transform 1 0 2944 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0952_
timestamp 1
transform 1 0 1380 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0953_
timestamp 1
transform 1 0 3404 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0954_
timestamp 1
transform -1 0 6992 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0955_
timestamp 1
transform -1 0 6808 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0956_
timestamp 1
transform 1 0 8924 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0957_
timestamp 1
transform -1 0 8556 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0958_
timestamp 1
transform -1 0 8188 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0959_
timestamp 1
transform 1 0 6532 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0960_
timestamp 1
transform 1 0 6348 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0961_
timestamp 1
transform 1 0 8648 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0962_
timestamp 1
transform 1 0 12144 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0963_
timestamp 1
transform 1 0 10304 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0964_
timestamp 1
transform 1 0 9568 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0965_
timestamp 1
transform -1 0 13984 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0966_
timestamp 1
transform -1 0 13064 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0967_
timestamp 1
transform 1 0 13064 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0968_
timestamp 1
transform -1 0 15916 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _0969_
timestamp 1
transform 1 0 1380 0 1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _0970_
timestamp 1
transform 1 0 1840 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0971_
timestamp 1
transform 1 0 1472 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0972_
timestamp 1
transform 1 0 1748 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0973_
timestamp 1
transform 1 0 4140 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _0974_
timestamp 1
transform -1 0 8372 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _0975_
timestamp 1
transform 1 0 1472 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0976_
timestamp 1
transform -1 0 6900 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0977_
timestamp 1
transform 1 0 3680 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _0978_
timestamp 1
transform 1 0 1380 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _0979_
timestamp 1
transform 1 0 9752 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _0980_
timestamp 1
transform 1 0 9384 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _0981_
timestamp 1
transform 1 0 8096 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _0982_
timestamp 1
transform 1 0 7360 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _0983_
timestamp 1
transform 1 0 9200 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _0984_
timestamp 1
transform 1 0 8924 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _0985_
timestamp 1
transform 1 0 9200 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_2  _0986_
timestamp 1
transform 1 0 6900 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _0987_
timestamp 1
transform 1 0 9476 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_2  _0988_
timestamp 1
transform 1 0 8924 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _0989_
timestamp 1
transform 1 0 7912 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_2  _0990_
timestamp 1
transform 1 0 7728 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _0991_
timestamp 1
transform 1 0 10212 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_2  _0992_
timestamp 1
transform 1 0 6992 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _0993_
timestamp 1
transform 1 0 9200 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_2  _0994_
timestamp 1
transform 1 0 6900 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _0995_
timestamp 1
transform 1 0 14812 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _0996_
timestamp 1
transform 1 0 14628 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _0997_
timestamp 1
transform 1 0 15916 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _0998_
timestamp 1
transform 1 0 16928 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _0999_
timestamp 1
transform 1 0 17480 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _1000_
timestamp 1
transform 1 0 16928 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _1001_
timestamp 1
transform 1 0 13524 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _1002_
timestamp 1
transform 1 0 14996 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _1003_
timestamp 1
transform 1 0 5336 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _1004_
timestamp 1
transform 1 0 4968 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _1005_
timestamp 1
transform -1 0 6900 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _1006_
timestamp 1
transform 1 0 4876 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _1007_
timestamp 1
transform 1 0 4048 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _1008_
timestamp 1
transform 1 0 1932 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _1009_
timestamp 1
transform 1 0 1380 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _1010_
timestamp 1
transform 1 0 1656 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _1011_
timestamp 1
transform 1 0 1380 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1012_
timestamp 1
transform 1 0 17756 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1013_
timestamp 1
transform -1 0 16376 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1014_
timestamp 1
transform -1 0 16284 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1015_
timestamp 1
transform 1 0 16744 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1016_
timestamp 1
transform 1 0 19228 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1017_
timestamp 1
transform -1 0 21712 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1018_
timestamp 1
transform 1 0 21988 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1019_
timestamp 1
transform 1 0 23000 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1020_
timestamp 1
transform 1 0 22632 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1021_
timestamp 1
transform -1 0 23368 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1022_
timestamp 1
transform 1 0 15364 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1023_
timestamp 1
transform 1 0 19228 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1024_
timestamp 1
transform 1 0 19504 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1025_
timestamp 1
transform 1 0 15548 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1026_
timestamp 1
transform 1 0 18400 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 1
transform 1 0 12880 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_clk
timestamp 1
transform -1 0 5520 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_clk
timestamp 1
transform -1 0 8832 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_clk
timestamp 1
transform 1 0 3772 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_clk
timestamp 1
transform 1 0 7820 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_clk
timestamp 1
transform -1 0 18952 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_clk
timestamp 1
transform 1 0 20424 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_clk
timestamp 1
transform -1 0 17480 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_clk
timestamp 1
transform 1 0 20516 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_4  clkload0
timestamp 1
transform 1 0 3772 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_8  clkload1
timestamp 1
transform 1 0 3772 0 1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_2  clkload2
timestamp 1
transform 1 0 6716 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_4  clkload3
timestamp 1
transform 1 0 15456 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__inv_8  clkload4
timestamp 1
transform 1 0 20424 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__inv_6  clkload5
timestamp 1
transform 1 0 15640 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__inv_6  clkload6
timestamp 1
transform 1 0 20516 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  fanout20
timestamp 1
transform -1 0 18952 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout21
timestamp 1
transform -1 0 8832 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout22
timestamp 1
transform 1 0 13432 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout23
timestamp 1
transform -1 0 4324 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout25
timestamp 1
transform -1 0 4324 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout26
timestamp 1
transform -1 0 6900 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout27
timestamp 1
transform -1 0 8096 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout28
timestamp 1
transform 1 0 10304 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout29
timestamp 1
transform -1 0 10948 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout30
timestamp 1
transform 1 0 7728 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout31
timestamp 1
transform 1 0 6900 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout32
timestamp 1
transform -1 0 9476 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout33
timestamp 1
transform 1 0 11684 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout34
timestamp 1
transform -1 0 10948 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout35
timestamp 1
transform 1 0 18400 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout36
timestamp 1
transform -1 0 20148 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout37
timestamp 1
transform 1 0 24380 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout38
timestamp 1
transform -1 0 18400 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout39
timestamp 1
transform 1 0 21344 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3
timestamp 1636968456
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1636968456
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp 1
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1636968456
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1636968456
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp 1
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1636968456
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1636968456
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1636968456
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1636968456
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1636968456
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1636968456
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1636968456
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1636968456
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1636968456
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1636968456
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1636968456
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1636968456
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1636968456
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1636968456
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_253
timestamp 1
transform 1 0 24380 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1636968456
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1636968456
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1636968456
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1636968456
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1636968456
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1636968456
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1636968456
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1636968456
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1636968456
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1636968456
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1636968456
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1636968456
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1636968456
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1636968456
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1636968456
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1636968456
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1636968456
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1636968456
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_249
timestamp 1
transform 1 0 24012 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_257
timestamp 1
transform 1 0 24748 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1636968456
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1636968456
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1636968456
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1636968456
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1636968456
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1636968456
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1636968456
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1636968456
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1636968456
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1636968456
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_144
timestamp 1
transform 1 0 14352 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_151
timestamp 1636968456
transform 1 0 14996 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_163
timestamp 1636968456
transform 1 0 16100 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_175
timestamp 1636968456
transform 1 0 17204 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_187
timestamp 1
transform 1 0 18308 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1636968456
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1636968456
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1636968456
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1636968456
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_253
timestamp 1
transform 1 0 24380 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1636968456
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1636968456
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1636968456
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1636968456
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1636968456
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1636968456
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1636968456
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1636968456
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1636968456
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_125
timestamp 1
transform 1 0 12604 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_146
timestamp 1
transform 1 0 14536 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_165
timestamp 1
transform 1 0 16284 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1636968456
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1636968456
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1636968456
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1636968456
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1636968456
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1636968456
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_249
timestamp 1
transform 1 0 24012 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_257
timestamp 1
transform 1 0 24748 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1636968456
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1636968456
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1636968456
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1636968456
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1636968456
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1636968456
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1636968456
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1636968456
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1636968456
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_121
timestamp 1
transform 1 0 12236 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_125
timestamp 1
transform 1 0 12604 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1636968456
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1636968456
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1636968456
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1636968456
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1636968456
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1636968456
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1636968456
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1636968456
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_253
timestamp 1
transform 1 0 24380 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1636968456
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1636968456
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_27
timestamp 1
transform 1 0 3588 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_48
timestamp 1
transform 1 0 5520 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_63
timestamp 1
transform 1 0 6900 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_71
timestamp 1
transform 1 0 7636 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_95
timestamp 1636968456
transform 1 0 9844 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_107
timestamp 1
transform 1 0 10948 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_120
timestamp 1
transform 1 0 12144 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_144
timestamp 1636968456
transform 1 0 14352 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_156
timestamp 1
transform 1 0 15456 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_163
timestamp 1
transform 1 0 16100 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1636968456
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1636968456
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_193
timestamp 1
transform 1 0 18860 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_201
timestamp 1
transform 1 0 19596 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_207
timestamp 1636968456
transform 1 0 20148 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_219
timestamp 1
transform 1 0 21252 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1636968456
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1636968456
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_249
timestamp 1
transform 1 0 24012 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_257
timestamp 1
transform 1 0 24748 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3
timestamp 1
transform 1 0 1380 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_24
timestamp 1
transform 1 0 3312 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1636968456
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_41
timestamp 1
transform 1 0 4876 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1636968456
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_97
timestamp 1
transform 1 0 10028 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_126
timestamp 1
transform 1 0 12696 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_141
timestamp 1
transform 1 0 14076 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_145
timestamp 1
transform 1 0 14444 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_153
timestamp 1
transform 1 0 15180 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_173
timestamp 1
transform 1 0 17020 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_180
timestamp 1
transform 1 0 17664 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_186
timestamp 1
transform 1 0 18216 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_218
timestamp 1636968456
transform 1 0 21160 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_230
timestamp 1636968456
transform 1 0 22264 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_242
timestamp 1
transform 1 0 23368 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_250
timestamp 1
transform 1 0 24104 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_253
timestamp 1
transform 1 0 24380 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_32
timestamp 1636968456
transform 1 0 4048 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_44
timestamp 1636968456
transform 1 0 5152 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_66
timestamp 1
transform 1 0 7176 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_7_93
timestamp 1
transform 1 0 9660 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_99
timestamp 1
transform 1 0 10212 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_106
timestamp 1
transform 1 0 10856 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_7_116
timestamp 1
transform 1 0 11776 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_122
timestamp 1
transform 1 0 12328 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_138
timestamp 1
transform 1 0 13800 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_145
timestamp 1
transform 1 0 14444 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_154
timestamp 1
transform 1 0 15272 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1636968456
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1636968456
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_249
timestamp 1
transform 1 0 24012 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_257
timestamp 1
transform 1 0 24748 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3
timestamp 1
transform 1 0 1380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_29
timestamp 1
transform 1 0 3772 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_40
timestamp 1
transform 1 0 4784 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_56
timestamp 1
transform 1 0 6256 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_64
timestamp 1
transform 1 0 6992 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_85
timestamp 1
transform 1 0 8924 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_109
timestamp 1
transform 1 0 11132 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_131
timestamp 1
transform 1 0 13156 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1636968456
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_153
timestamp 1
transform 1 0 15180 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_157
timestamp 1
transform 1 0 15548 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_167
timestamp 1
transform 1 0 16468 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_186
timestamp 1
transform 1 0 18216 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_218
timestamp 1636968456
transform 1 0 21160 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_230
timestamp 1636968456
transform 1 0 22264 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_242
timestamp 1
transform 1 0 23368 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_250
timestamp 1
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_253
timestamp 1
transform 1 0 24380 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1636968456
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_15
timestamp 1
transform 1 0 2484 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_24
timestamp 1
transform 1 0 3312 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_46
timestamp 1
transform 1 0 5336 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_64
timestamp 1636968456
transform 1 0 6992 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_76
timestamp 1
transform 1 0 8096 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_80
timestamp 1
transform 1 0 8464 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_90
timestamp 1
transform 1 0 9384 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_107
timestamp 1
transform 1 0 10948 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_113
timestamp 1
transform 1 0 11500 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_127
timestamp 1
transform 1 0 12788 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_136
timestamp 1
transform 1 0 13616 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_142
timestamp 1
transform 1 0 14168 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_151
timestamp 1636968456
transform 1 0 14996 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_163
timestamp 1
transform 1 0 16100 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_169
timestamp 1
transform 1 0 16652 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_179
timestamp 1
transform 1 0 17572 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_203
timestamp 1636968456
transform 1 0 19780 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_215
timestamp 1
transform 1 0 20884 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1636968456
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1636968456
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_249
timestamp 1
transform 1 0 24012 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_257
timestamp 1
transform 1 0 24748 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1636968456
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_36
timestamp 1
transform 1 0 4416 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_44
timestamp 1
transform 1 0 5152 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_71
timestamp 1636968456
transform 1 0 7636 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1636968456
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1636968456
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1636968456
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_121
timestamp 1
transform 1 0 12236 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_127
timestamp 1
transform 1 0 12788 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_141
timestamp 1
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_164
timestamp 1636968456
transform 1 0 16192 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_176
timestamp 1636968456
transform 1 0 17296 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1636968456
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1636968456
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1636968456
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1636968456
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_253
timestamp 1
transform 1 0 24380 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_11_3
timestamp 1
transform 1 0 1380 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_11
timestamp 1
transform 1 0 2116 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_41
timestamp 1
transform 1 0 4876 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_47
timestamp 1
transform 1 0 5428 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_52
timestamp 1
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_57
timestamp 1
transform 1 0 6348 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_63
timestamp 1
transform 1 0 6900 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_106
timestamp 1
transform 1 0 10856 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_11_113
timestamp 1
transform 1 0 11500 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_121
timestamp 1
transform 1 0 12236 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_127
timestamp 1
transform 1 0 12788 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_133
timestamp 1
transform 1 0 13340 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_138
timestamp 1636968456
transform 1 0 13800 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_150
timestamp 1636968456
transform 1 0 14904 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_162
timestamp 1
transform 1 0 16008 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_169
timestamp 1
transform 1 0 16652 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_182
timestamp 1636968456
transform 1 0 17848 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_194
timestamp 1636968456
transform 1 0 18952 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_206
timestamp 1
transform 1 0 20056 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_213
timestamp 1
transform 1 0 20700 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_221
timestamp 1
transform 1 0 21436 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1636968456
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1636968456
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_249
timestamp 1
transform 1 0 24012 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_257
timestamp 1
transform 1 0 24748 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1636968456
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_15
timestamp 1
transform 1 0 2484 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_39
timestamp 1
transform 1 0 4692 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_57
timestamp 1
transform 1 0 6348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_79
timestamp 1
transform 1 0 8372 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_94
timestamp 1
transform 1 0 9752 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_98
timestamp 1
transform 1 0 10120 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_120
timestamp 1
transform 1 0 12144 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_137
timestamp 1
transform 1 0 13708 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_141
timestamp 1
transform 1 0 14076 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_149
timestamp 1
transform 1 0 14812 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_193
timestamp 1
transform 1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_226
timestamp 1636968456
transform 1 0 21896 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_238
timestamp 1636968456
transform 1 0 23000 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_250
timestamp 1
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_253
timestamp 1
transform 1 0 24380 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1636968456
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_15
timestamp 1
transform 1 0 2484 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_53
timestamp 1
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_69
timestamp 1
transform 1 0 7452 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_13_84
timestamp 1
transform 1 0 8832 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_90
timestamp 1
transform 1 0 9384 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_122
timestamp 1636968456
transform 1 0 12328 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_134
timestamp 1
transform 1 0 13432 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_164
timestamp 1
transform 1 0 16192 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_199
timestamp 1
transform 1 0 19412 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_207
timestamp 1
transform 1 0 20148 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_221
timestamp 1
transform 1 0 21436 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_230
timestamp 1636968456
transform 1 0 22264 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_242
timestamp 1636968456
transform 1 0 23368 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_254
timestamp 1
transform 1 0 24472 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_258
timestamp 1
transform 1 0 24840 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_3
timestamp 1
transform 1 0 1380 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp 1
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_42
timestamp 1636968456
transform 1 0 4968 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_59
timestamp 1
transform 1 0 6532 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_63
timestamp 1
transform 1 0 6900 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_85
timestamp 1
transform 1 0 8924 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_91
timestamp 1
transform 1 0 9476 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_110
timestamp 1636968456
transform 1 0 11224 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_122
timestamp 1
transform 1 0 12328 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_149
timestamp 1
transform 1 0 14812 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_160
timestamp 1
transform 1 0 15824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_193
timestamp 1
transform 1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_205
timestamp 1
transform 1 0 19964 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_237
timestamp 1636968456
transform 1 0 22908 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_249
timestamp 1
transform 1 0 24012 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_14_253
timestamp 1
transform 1 0 24380 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1636968456
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_15
timestamp 1
transform 1 0 2484 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_24
timestamp 1
transform 1 0 3312 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_48
timestamp 1
transform 1 0 5520 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_57
timestamp 1
transform 1 0 6348 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_65
timestamp 1
transform 1 0 7084 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_89
timestamp 1636968456
transform 1 0 9292 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_101
timestamp 1
transform 1 0 10396 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_109
timestamp 1
transform 1 0 11132 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1636968456
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_125
timestamp 1
transform 1 0 12604 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_146
timestamp 1
transform 1 0 14536 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_154
timestamp 1
transform 1 0 15272 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_163
timestamp 1
transform 1 0 16100 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_169
timestamp 1
transform 1 0 16652 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_173
timestamp 1
transform 1 0 17020 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_183
timestamp 1636968456
transform 1 0 17940 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_195
timestamp 1636968456
transform 1 0 19044 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_207
timestamp 1
transform 1 0 20148 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_225
timestamp 1
transform 1 0 21804 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_229
timestamp 1
transform 1 0 22172 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_235
timestamp 1636968456
transform 1 0 22724 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_247
timestamp 1636968456
transform 1 0 23828 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_39
timestamp 1
transform 1 0 4692 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_85
timestamp 1
transform 1 0 8924 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_93
timestamp 1
transform 1 0 9660 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_107
timestamp 1636968456
transform 1 0 10948 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_119
timestamp 1
transform 1 0 12052 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_125
timestamp 1
transform 1 0 12604 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1636968456
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_197
timestamp 1
transform 1 0 19228 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_216
timestamp 1
transform 1 0 20976 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_233
timestamp 1636968456
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_253
timestamp 1
transform 1 0 24380 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_17
timestamp 1
transform 1 0 2668 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_66
timestamp 1
transform 1 0 7176 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_17_81
timestamp 1
transform 1 0 8556 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_87
timestamp 1
transform 1 0 9108 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_109
timestamp 1
transform 1 0 11132 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_113
timestamp 1
transform 1 0 11500 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_130
timestamp 1
transform 1 0 13064 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_134
timestamp 1
transform 1 0 13432 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_142
timestamp 1636968456
transform 1 0 14168 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_154
timestamp 1636968456
transform 1 0 15272 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1636968456
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_181
timestamp 1
transform 1 0 17756 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_201
timestamp 1
transform 1 0 19596 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_212
timestamp 1636968456
transform 1 0 20608 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_225
timestamp 1
transform 1 0 21804 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_232
timestamp 1636968456
transform 1 0 22448 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_244
timestamp 1636968456
transform 1 0 23552 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_256
timestamp 1
transform 1 0 24656 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_26
timestamp 1
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_50
timestamp 1636968456
transform 1 0 5704 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_62
timestamp 1636968456
transform 1 0 6808 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_74
timestamp 1
transform 1 0 7912 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_106
timestamp 1
transform 1 0 10856 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_116
timestamp 1
transform 1 0 11776 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_131
timestamp 1
transform 1 0 13156 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_141
timestamp 1
transform 1 0 14076 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_170
timestamp 1
transform 1 0 16744 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_174
timestamp 1
transform 1 0 17112 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_208
timestamp 1
transform 1 0 20240 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_253
timestamp 1
transform 1 0 24380 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1636968456
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_15
timestamp 1
transform 1 0 2484 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_23
timestamp 1
transform 1 0 3220 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_34
timestamp 1
transform 1 0 4232 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_19_49
timestamp 1
transform 1 0 5612 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_78
timestamp 1
transform 1 0 8280 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_86
timestamp 1
transform 1 0 9016 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_96
timestamp 1636968456
transform 1 0 9936 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_108
timestamp 1
transform 1 0 11040 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_113
timestamp 1
transform 1 0 11500 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_122
timestamp 1636968456
transform 1 0 12328 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_134
timestamp 1636968456
transform 1 0 13432 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_146
timestamp 1
transform 1 0 14536 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_205
timestamp 1
transform 1 0 19964 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_213
timestamp 1
transform 1 0 20700 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_255
timestamp 1
transform 1 0 24564 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1636968456
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_15
timestamp 1
transform 1 0 2484 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1636968456
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_94
timestamp 1636968456
transform 1 0 9752 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_106
timestamp 1
transform 1 0 10856 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_112
timestamp 1
transform 1 0 11408 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_120
timestamp 1636968456
transform 1 0 12144 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_132
timestamp 1
transform 1 0 13248 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_146
timestamp 1
transform 1 0 14536 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_154
timestamp 1
transform 1 0 15272 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_163
timestamp 1
transform 1 0 16100 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_178
timestamp 1
transform 1 0 17480 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_192
timestamp 1
transform 1 0 18768 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1636968456
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_209
timestamp 1
transform 1 0 20332 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_215
timestamp 1
transform 1 0 20884 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_6
timestamp 1
transform 1 0 1656 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_30
timestamp 1
transform 1 0 3864 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_53
timestamp 1
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_75
timestamp 1
transform 1 0 8004 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_106
timestamp 1
transform 1 0 10856 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_21_113
timestamp 1
transform 1 0 11500 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_130
timestamp 1
transform 1 0 13064 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_134
timestamp 1
transform 1 0 13432 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_139
timestamp 1636968456
transform 1 0 13892 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_151
timestamp 1636968456
transform 1 0 14996 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_163
timestamp 1
transform 1 0 16100 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_169
timestamp 1
transform 1 0 16652 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_175
timestamp 1
transform 1 0 17204 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_179
timestamp 1
transform 1 0 17572 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_188
timestamp 1636968456
transform 1 0 18400 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_200
timestamp 1636968456
transform 1 0 19504 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_212
timestamp 1636968456
transform 1 0 20608 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_240
timestamp 1636968456
transform 1 0 23184 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_252
timestamp 1
transform 1 0 24288 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_258
timestamp 1
transform 1 0 24840 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_24
timestamp 1
transform 1 0 3312 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_29
timestamp 1
transform 1 0 3772 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_76
timestamp 1
transform 1 0 8096 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_85
timestamp 1
transform 1 0 8924 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_109
timestamp 1
transform 1 0 11132 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_137
timestamp 1
transform 1 0 13708 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_146
timestamp 1
transform 1 0 14536 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_159
timestamp 1636968456
transform 1 0 15732 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_171
timestamp 1
transform 1 0 16836 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_175
timestamp 1
transform 1 0 17204 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_185
timestamp 1
transform 1 0 18124 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_193
timestamp 1
transform 1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1636968456
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_209
timestamp 1
transform 1 0 20332 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_219
timestamp 1
transform 1 0 21252 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_223
timestamp 1
transform 1 0 21620 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_232
timestamp 1
transform 1 0 22448 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_243
timestamp 1
transform 1 0 23460 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_253
timestamp 1
transform 1 0 24380 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_23_3
timestamp 1
transform 1 0 1380 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_11
timestamp 1
transform 1 0 2116 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_44
timestamp 1636968456
transform 1 0 5152 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_66
timestamp 1
transform 1 0 7176 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_113
timestamp 1
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_169
timestamp 1
transform 1 0 16652 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_193
timestamp 1
transform 1 0 18860 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_220
timestamp 1
transform 1 0 21344 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_225
timestamp 1
transform 1 0 21804 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_231
timestamp 1
transform 1 0 22356 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_238
timestamp 1
transform 1 0 23000 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_38
timestamp 1
transform 1 0 4600 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_69
timestamp 1
transform 1 0 7452 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_80
timestamp 1
transform 1 0 8464 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_119
timestamp 1
transform 1 0 12052 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_127
timestamp 1
transform 1 0 12788 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_160
timestamp 1
transform 1 0 15824 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_188
timestamp 1
transform 1 0 18400 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_197
timestamp 1
transform 1 0 19228 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_204
timestamp 1
transform 1 0 19872 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_235
timestamp 1
transform 1 0 22724 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_3
timestamp 1
transform 1 0 1380 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_11
timestamp 1
transform 1 0 2116 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_23
timestamp 1636968456
transform 1 0 3220 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_35
timestamp 1636968456
transform 1 0 4324 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_66
timestamp 1
transform 1 0 7176 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_25_90
timestamp 1
transform 1 0 9384 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_96
timestamp 1
transform 1 0 9936 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_106
timestamp 1
transform 1 0 10856 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1636968456
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_125
timestamp 1
transform 1 0 12604 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_133
timestamp 1
transform 1 0 13340 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_144
timestamp 1
transform 1 0 14352 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_154
timestamp 1
transform 1 0 15272 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_163
timestamp 1
transform 1 0 16100 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1636968456
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_181
timestamp 1
transform 1 0 17756 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_187
timestamp 1
transform 1 0 18308 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_208
timestamp 1
transform 1 0 20240 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_212
timestamp 1
transform 1 0 20608 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_219
timestamp 1
transform 1 0 21252 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_233
timestamp 1
transform 1 0 22540 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_256
timestamp 1
transform 1 0 24656 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_24
timestamp 1
transform 1 0 3312 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1636968456
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_41
timestamp 1
transform 1 0 4876 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_45
timestamp 1
transform 1 0 5244 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_67
timestamp 1
transform 1 0 7268 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_80
timestamp 1
transform 1 0 8464 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_91
timestamp 1636968456
transform 1 0 9476 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_103
timestamp 1636968456
transform 1 0 10580 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_115
timestamp 1636968456
transform 1 0 11684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_127
timestamp 1636968456
transform 1 0 12788 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1636968456
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1636968456
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1636968456
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1636968456
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1636968456
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1636968456
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_221
timestamp 1
transform 1 0 21436 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_233
timestamp 1636968456
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_253
timestamp 1
transform 1 0 24380 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1
transform 1 0 1380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_7
timestamp 1
transform 1 0 1748 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_38
timestamp 1636968456
transform 1 0 4600 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_50
timestamp 1
transform 1 0 5704 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1636968456
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1636968456
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_81
timestamp 1
transform 1 0 8556 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_89
timestamp 1
transform 1 0 9292 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1636968456
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1636968456
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1636968456
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_149
timestamp 1
transform 1 0 14812 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_157
timestamp 1
transform 1 0 15548 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_163
timestamp 1
transform 1 0 16100 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_169
timestamp 1
transform 1 0 16652 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_194
timestamp 1636968456
transform 1 0 18952 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_206
timestamp 1636968456
transform 1 0 20056 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_218
timestamp 1
transform 1 0 21160 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1636968456
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_237
timestamp 1636968456
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_249
timestamp 1
transform 1 0 24012 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_257
timestamp 1
transform 1 0 24748 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_24
timestamp 1
transform 1 0 3312 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_37
timestamp 1636968456
transform 1 0 4508 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_49
timestamp 1636968456
transform 1 0 5612 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_61
timestamp 1636968456
transform 1 0 6716 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_73
timestamp 1
transform 1 0 7820 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_81
timestamp 1
transform 1 0 8556 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1636968456
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_97
timestamp 1
transform 1 0 10028 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_141
timestamp 1
transform 1 0 14076 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_145
timestamp 1
transform 1 0 14444 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_166
timestamp 1
transform 1 0 16376 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_176
timestamp 1636968456
transform 1 0 17296 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_217
timestamp 1636968456
transform 1 0 21068 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_229
timestamp 1636968456
transform 1 0 22172 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_241
timestamp 1
transform 1 0 23276 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_249
timestamp 1
transform 1 0 24012 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_28_253
timestamp 1
transform 1 0 24380 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1636968456
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_15
timestamp 1
transform 1 0 2484 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_22
timestamp 1
transform 1 0 3128 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_57
timestamp 1
transform 1 0 6348 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_65
timestamp 1
transform 1 0 7084 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_78
timestamp 1
transform 1 0 8280 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_102
timestamp 1
transform 1 0 10488 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_106
timestamp 1
transform 1 0 10856 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_113
timestamp 1
transform 1 0 11500 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_122
timestamp 1
transform 1 0 12328 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_140
timestamp 1
transform 1 0 13984 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_144
timestamp 1
transform 1 0 14352 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_165
timestamp 1
transform 1 0 16284 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_202
timestamp 1
transform 1 0 19688 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_232
timestamp 1636968456
transform 1 0 22448 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_244
timestamp 1636968456
transform 1 0 23552 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_256
timestamp 1
transform 1 0 24656 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1636968456
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_15
timestamp 1
transform 1 0 2484 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_19
timestamp 1
transform 1 0 2852 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_29
timestamp 1
transform 1 0 3772 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_51
timestamp 1
transform 1 0 5796 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_95
timestamp 1636968456
transform 1 0 9844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_107
timestamp 1
transform 1 0 10948 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_115
timestamp 1
transform 1 0 11684 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_136
timestamp 1
transform 1 0 13616 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_141
timestamp 1
transform 1 0 14076 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_149
timestamp 1
transform 1 0 14812 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_175
timestamp 1
transform 1 0 17204 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_183
timestamp 1
transform 1 0 17940 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_203
timestamp 1
transform 1 0 19780 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_225
timestamp 1
transform 1 0 21804 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_247
timestamp 1
transform 1 0 23828 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_253
timestamp 1
transform 1 0 24380 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_31_3
timestamp 1
transform 1 0 1380 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_11
timestamp 1
transform 1 0 2116 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_52
timestamp 1
transform 1 0 5888 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_57
timestamp 1
transform 1 0 6348 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_72
timestamp 1
transform 1 0 7728 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_100
timestamp 1636968456
transform 1 0 10304 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_113
timestamp 1
transform 1 0 11500 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_129
timestamp 1636968456
transform 1 0 12972 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_141
timestamp 1636968456
transform 1 0 14076 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_153
timestamp 1
transform 1 0 15180 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_157
timestamp 1
transform 1 0 15548 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1636968456
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1636968456
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_193
timestamp 1
transform 1 0 18860 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_199
timestamp 1
transform 1 0 19412 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_205
timestamp 1
transform 1 0 19964 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_211
timestamp 1
transform 1 0 20516 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_218
timestamp 1
transform 1 0 21160 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_232
timestamp 1636968456
transform 1 0 22448 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_244
timestamp 1636968456
transform 1 0 23552 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_256
timestamp 1
transform 1 0 24656 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_32_50
timestamp 1
transform 1 0 5704 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_56
timestamp 1
transform 1 0 6256 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_90
timestamp 1
transform 1 0 9384 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_99
timestamp 1636968456
transform 1 0 10212 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_111
timestamp 1
transform 1 0 11316 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_115
timestamp 1
transform 1 0 11684 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1636968456
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_153
timestamp 1
transform 1 0 15180 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_161
timestamp 1
transform 1 0 15916 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_168
timestamp 1636968456
transform 1 0 16560 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_180
timestamp 1636968456
transform 1 0 17664 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_192
timestamp 1
transform 1 0 18768 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_205
timestamp 1
transform 1 0 19964 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_212
timestamp 1636968456
transform 1 0 20608 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_224
timestamp 1636968456
transform 1 0 21712 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_236
timestamp 1636968456
transform 1 0 22816 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_248
timestamp 1
transform 1 0 23920 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_253
timestamp 1
transform 1 0 24380 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_33_3
timestamp 1
transform 1 0 1380 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_11
timestamp 1
transform 1 0 2116 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_57
timestamp 1
transform 1 0 6348 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_65
timestamp 1
transform 1 0 7084 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_84
timestamp 1
transform 1 0 8832 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_92
timestamp 1
transform 1 0 9568 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_102
timestamp 1
transform 1 0 10488 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1636968456
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_140
timestamp 1636968456
transform 1 0 13984 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_152
timestamp 1
transform 1 0 15088 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_180
timestamp 1
transform 1 0 17664 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_189
timestamp 1
transform 1 0 18492 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_194
timestamp 1
transform 1 0 18952 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_198
timestamp 1
transform 1 0 19320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_206
timestamp 1
transform 1 0 20056 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_210
timestamp 1
transform 1 0 20424 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_220
timestamp 1
transform 1 0 21344 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_225
timestamp 1
transform 1 0 21804 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_235
timestamp 1
transform 1 0 22724 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_33_258
timestamp 1
transform 1 0 24840 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_34_39
timestamp 1
transform 1 0 4692 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_62
timestamp 1636968456
transform 1 0 6808 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_74
timestamp 1
transform 1 0 7912 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_85
timestamp 1
transform 1 0 8924 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_89
timestamp 1
transform 1 0 9292 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_111
timestamp 1636968456
transform 1 0 11316 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_123
timestamp 1
transform 1 0 12420 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_129
timestamp 1
transform 1 0 12972 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_34_137
timestamp 1
transform 1 0 13708 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1636968456
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_178
timestamp 1
transform 1 0 17480 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_187
timestamp 1
transform 1 0 18308 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_210
timestamp 1
transform 1 0 20424 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_231
timestamp 1
transform 1 0 22356 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_246
timestamp 1
transform 1 0 23736 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_34_253
timestamp 1
transform 1 0 24380 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1636968456
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1636968456
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_27
timestamp 1
transform 1 0 3588 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_33
timestamp 1
transform 1 0 4140 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_44
timestamp 1
transform 1 0 5152 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_57
timestamp 1
transform 1 0 6348 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_68
timestamp 1
transform 1 0 7360 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_84
timestamp 1636968456
transform 1 0 8832 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_96
timestamp 1636968456
transform 1 0 9936 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_108
timestamp 1
transform 1 0 11040 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_130
timestamp 1
transform 1 0 13064 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_138
timestamp 1636968456
transform 1 0 13800 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_150
timestamp 1
transform 1 0 14904 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_165
timestamp 1
transform 1 0 16284 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_178
timestamp 1
transform 1 0 17480 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_182
timestamp 1
transform 1 0 17848 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_192
timestamp 1
transform 1 0 18768 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_200
timestamp 1
transform 1 0 19504 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_35_210
timestamp 1
transform 1 0 20424 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_232
timestamp 1
transform 1 0 22448 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_254
timestamp 1
transform 1 0 24472 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_258
timestamp 1
transform 1 0 24840 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1636968456
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1636968456
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1636968456
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_41
timestamp 1
transform 1 0 4876 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_36_62
timestamp 1
transform 1 0 6808 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_70
timestamp 1
transform 1 0 7544 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_79
timestamp 1
transform 1 0 8372 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_85
timestamp 1
transform 1 0 8924 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_94
timestamp 1636968456
transform 1 0 9752 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_106
timestamp 1
transform 1 0 10856 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_36_133
timestamp 1
transform 1 0 13340 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_141
timestamp 1
transform 1 0 14076 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_149
timestamp 1
transform 1 0 14812 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_203
timestamp 1
transform 1 0 19780 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_223
timestamp 1
transform 1 0 21620 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_240
timestamp 1636968456
transform 1 0 23184 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_253
timestamp 1
transform 1 0 24380 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_3
timestamp 1
transform 1 0 1380 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_7
timestamp 1
transform 1 0 1748 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_28
timestamp 1636968456
transform 1 0 3680 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_40
timestamp 1636968456
transform 1 0 4784 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_52
timestamp 1
transform 1 0 5888 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_77
timestamp 1
transform 1 0 8188 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_81
timestamp 1
transform 1 0 8556 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_102
timestamp 1
transform 1 0 10488 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_113
timestamp 1
transform 1 0 11500 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_117
timestamp 1
transform 1 0 11868 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_125
timestamp 1
transform 1 0 12604 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_37_147
timestamp 1
transform 1 0 14628 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_155
timestamp 1
transform 1 0 15364 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_159
timestamp 1
transform 1 0 15732 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_37_169
timestamp 1
transform 1 0 16652 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_178
timestamp 1636968456
transform 1 0 17480 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_190
timestamp 1636968456
transform 1 0 18584 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_202
timestamp 1636968456
transform 1 0 19688 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_214
timestamp 1
transform 1 0 20792 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_222
timestamp 1
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_235
timestamp 1636968456
transform 1 0 22724 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_247
timestamp 1636968456
transform 1 0 23828 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_26
timestamp 1
transform 1 0 3496 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_40
timestamp 1636968456
transform 1 0 4784 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_52
timestamp 1636968456
transform 1 0 5888 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_64
timestamp 1
transform 1 0 6992 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_38_75
timestamp 1
transform 1 0 8004 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_38_85
timestamp 1
transform 1 0 8924 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_92
timestamp 1
transform 1 0 9568 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_38_102
timestamp 1
transform 1 0 10488 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_109
timestamp 1
transform 1 0 11132 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_116
timestamp 1636968456
transform 1 0 11776 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_128
timestamp 1
transform 1 0 12880 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_134
timestamp 1
transform 1 0 13432 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_38_164
timestamp 1
transform 1 0 16192 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_188
timestamp 1
transform 1 0 18400 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1636968456
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1636968456
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_221
timestamp 1636968456
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_233
timestamp 1636968456
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_245
timestamp 1
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_253
timestamp 1
transform 1 0 24380 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_39_3
timestamp 1
transform 1 0 1380 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_23
timestamp 1
transform 1 0 3220 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_53
timestamp 1
transform 1 0 5980 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_39_57
timestamp 1
transform 1 0 6348 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_75
timestamp 1
transform 1 0 8004 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_85
timestamp 1636968456
transform 1 0 8924 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_97
timestamp 1
transform 1 0 10028 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_103
timestamp 1
transform 1 0 10580 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_131
timestamp 1636968456
transform 1 0 13156 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_143
timestamp 1636968456
transform 1 0 14260 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_155
timestamp 1636968456
transform 1 0 15364 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_175
timestamp 1
transform 1 0 17204 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_181
timestamp 1
transform 1 0 17756 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_188
timestamp 1
transform 1 0 18400 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_211
timestamp 1
transform 1 0 20516 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_220
timestamp 1
transform 1 0 21344 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_239
timestamp 1636968456
transform 1 0 23092 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_251
timestamp 1
transform 1 0 24196 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_40_3
timestamp 1
transform 1 0 1380 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_40_64
timestamp 1
transform 1 0 6992 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_82
timestamp 1
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1636968456
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_97
timestamp 1
transform 1 0 10028 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_113
timestamp 1
transform 1 0 11500 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_121
timestamp 1
transform 1 0 12236 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_137
timestamp 1
transform 1 0 13708 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1636968456
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_153
timestamp 1
transform 1 0 15180 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_183
timestamp 1
transform 1 0 17940 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_187
timestamp 1
transform 1 0 18308 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_242
timestamp 1
transform 1 0 23368 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_250
timestamp 1
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_253
timestamp 1
transform 1 0 24380 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_3
timestamp 1
transform 1 0 1380 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_41_32
timestamp 1
transform 1 0 4048 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_41_53
timestamp 1
transform 1 0 5980 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_57
timestamp 1
transform 1 0 6348 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_98
timestamp 1636968456
transform 1 0 10120 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_110
timestamp 1
transform 1 0 11224 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_113
timestamp 1
transform 1 0 11500 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_121
timestamp 1
transform 1 0 12236 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_154
timestamp 1
transform 1 0 15272 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_187
timestamp 1
transform 1 0 18308 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_195
timestamp 1
transform 1 0 19044 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_41_199
timestamp 1
transform 1 0 19412 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_220
timestamp 1
transform 1 0 21344 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_235
timestamp 1636968456
transform 1 0 22724 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_247
timestamp 1636968456
transform 1 0 23828 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_3
timestamp 1
transform 1 0 1380 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_43
timestamp 1
transform 1 0 5060 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_55
timestamp 1636968456
transform 1 0 6164 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_67
timestamp 1
transform 1 0 7268 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_42_81
timestamp 1
transform 1 0 8556 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_42_105
timestamp 1
transform 1 0 10764 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_109
timestamp 1
transform 1 0 11132 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_42_137
timestamp 1
transform 1 0 13708 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1636968456
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_153
timestamp 1
transform 1 0 15180 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1636968456
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_217
timestamp 1636968456
transform 1 0 21068 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_229
timestamp 1636968456
transform 1 0 22172 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_241
timestamp 1
transform 1 0 23276 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_249
timestamp 1
transform 1 0 24012 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_42_253
timestamp 1
transform 1 0 24380 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1636968456
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1636968456
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_27
timestamp 1
transform 1 0 3588 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_35
timestamp 1636968456
transform 1 0 4324 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_47
timestamp 1
transform 1 0 5428 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1636968456
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1636968456
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_81
timestamp 1
transform 1 0 8556 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_85
timestamp 1
transform 1 0 8924 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_91
timestamp 1
transform 1 0 9476 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_43_98
timestamp 1
transform 1 0 10120 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_43_105
timestamp 1
transform 1 0 10764 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_113
timestamp 1
transform 1 0 11500 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_118
timestamp 1
transform 1 0 11960 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_43_126
timestamp 1
transform 1 0 12696 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_132
timestamp 1
transform 1 0 13248 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_141
timestamp 1
transform 1 0 14076 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_147
timestamp 1
transform 1 0 14628 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_43_154
timestamp 1
transform 1 0 15272 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_160
timestamp 1
transform 1 0 15824 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_169
timestamp 1
transform 1 0 16652 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_177
timestamp 1
transform 1 0 17388 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_43_182
timestamp 1
transform 1 0 17848 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_43_189
timestamp 1
transform 1 0 18492 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_195
timestamp 1
transform 1 0 19044 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_197
timestamp 1636968456
transform 1 0 19228 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_209
timestamp 1636968456
transform 1 0 20332 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_221
timestamp 1
transform 1 0 21436 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1636968456
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1636968456
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_249
timestamp 1
transform 1 0 24012 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_43_253
timestamp 1
transform 1 0 24380 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 1
transform 1 0 3772 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1
transform -1 0 6072 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1
transform -1 0 3588 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1
transform -1 0 6164 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1
transform -1 0 19136 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1
transform -1 0 22540 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1
transform -1 0 15824 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1
transform -1 0 4324 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1
transform -1 0 18216 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1
transform -1 0 4876 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1
transform -1 0 3220 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1
transform 1 0 3772 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1
transform -1 0 19964 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1
transform -1 0 16928 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1
transform -1 0 4048 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1
transform -1 0 6164 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1
transform 1 0 13616 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1
transform 1 0 12972 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1
transform 1 0 15548 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1
transform 1 0 16192 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1
transform 1 0 14904 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 1
transform 1 0 12328 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1
transform 1 0 9108 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1
transform 1 0 11684 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1
transform 1 0 14260 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1
transform 1 0 10396 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1
transform 1 0 11040 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1
transform 1 0 18124 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1
transform 1 0 9752 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1
transform 1 0 17480 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1
transform -1 0 1656 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1
transform -1 0 24932 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 1
transform 1 0 1380 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  matrix_mult_40
timestamp 1
transform 1 0 24656 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  max_cap24
timestamp 1
transform -1 0 21804 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output18
timestamp 1
transform -1 0 1748 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp 1
transform 1 0 24564 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_44
timestamp 1
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1
transform -1 0 25208 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_45
timestamp 1
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1
transform -1 0 25208 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_46
timestamp 1
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1
transform -1 0 25208 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_47
timestamp 1
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1
transform -1 0 25208 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_48
timestamp 1
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1
transform -1 0 25208 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_49
timestamp 1
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1
transform -1 0 25208 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_50
timestamp 1
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1
transform -1 0 25208 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_51
timestamp 1
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1
transform -1 0 25208 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_52
timestamp 1
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1
transform -1 0 25208 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_53
timestamp 1
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1
transform -1 0 25208 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_54
timestamp 1
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1
transform -1 0 25208 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_55
timestamp 1
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1
transform -1 0 25208 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_56
timestamp 1
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1
transform -1 0 25208 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_57
timestamp 1
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1
transform -1 0 25208 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_58
timestamp 1
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1
transform -1 0 25208 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_59
timestamp 1
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1
transform -1 0 25208 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_60
timestamp 1
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1
transform -1 0 25208 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_61
timestamp 1
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1
transform -1 0 25208 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_62
timestamp 1
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1
transform -1 0 25208 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_63
timestamp 1
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1
transform -1 0 25208 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_64
timestamp 1
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1
transform -1 0 25208 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_65
timestamp 1
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1
transform -1 0 25208 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_66
timestamp 1
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1
transform -1 0 25208 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_67
timestamp 1
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1
transform -1 0 25208 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_68
timestamp 1
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1
transform -1 0 25208 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_69
timestamp 1
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1
transform -1 0 25208 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_70
timestamp 1
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1
transform -1 0 25208 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_71
timestamp 1
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1
transform -1 0 25208 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_72
timestamp 1
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1
transform -1 0 25208 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_73
timestamp 1
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1
transform -1 0 25208 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_74
timestamp 1
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1
transform -1 0 25208 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_75
timestamp 1
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1
transform -1 0 25208 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_76
timestamp 1
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1
transform -1 0 25208 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_77
timestamp 1
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1
transform -1 0 25208 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_78
timestamp 1
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 1
transform -1 0 25208 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_79
timestamp 1
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 1
transform -1 0 25208 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_80
timestamp 1
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 1
transform -1 0 25208 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_81
timestamp 1
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 1
transform -1 0 25208 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_82
timestamp 1
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 1
transform -1 0 25208 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_83
timestamp 1
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp 1
transform -1 0 25208 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_84
timestamp 1
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp 1
transform -1 0 25208 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_85
timestamp 1
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp 1
transform -1 0 25208 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Left_86
timestamp 1
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Right_42
timestamp 1
transform -1 0 25208 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Left_87
timestamp 1
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Right_43
timestamp 1
transform -1 0 25208 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_88
timestamp 1
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_89
timestamp 1
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_90
timestamp 1
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_91
timestamp 1
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_92
timestamp 1
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_93
timestamp 1
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_94
timestamp 1
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_95
timestamp 1
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_96
timestamp 1
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_97
timestamp 1
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_98
timestamp 1
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_99
timestamp 1
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_100
timestamp 1
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_101
timestamp 1
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_102
timestamp 1
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_103
timestamp 1
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_104
timestamp 1
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_105
timestamp 1
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_106
timestamp 1
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_107
timestamp 1
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_108
timestamp 1
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_109
timestamp 1
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_110
timestamp 1
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_111
timestamp 1
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_112
timestamp 1
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_113
timestamp 1
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_114
timestamp 1
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_115
timestamp 1
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_116
timestamp 1
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_117
timestamp 1
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_118
timestamp 1
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_119
timestamp 1
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_120
timestamp 1
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_121
timestamp 1
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_122
timestamp 1
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_123
timestamp 1
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_124
timestamp 1
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_125
timestamp 1
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_126
timestamp 1
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_127
timestamp 1
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_128
timestamp 1
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_129
timestamp 1
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_130
timestamp 1
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_131
timestamp 1
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_132
timestamp 1
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_133
timestamp 1
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_134
timestamp 1
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_135
timestamp 1
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_136
timestamp 1
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_137
timestamp 1
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_138
timestamp 1
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_139
timestamp 1
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_140
timestamp 1
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_141
timestamp 1
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_142
timestamp 1
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_143
timestamp 1
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_144
timestamp 1
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_145
timestamp 1
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_146
timestamp 1
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_147
timestamp 1
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_148
timestamp 1
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_149
timestamp 1
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_150
timestamp 1
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_151
timestamp 1
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_152
timestamp 1
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_153
timestamp 1
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_154
timestamp 1
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_155
timestamp 1
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_156
timestamp 1
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_157
timestamp 1
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_158
timestamp 1
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_159
timestamp 1
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_160
timestamp 1
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_161
timestamp 1
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_162
timestamp 1
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_163
timestamp 1
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_164
timestamp 1
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_165
timestamp 1
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_166
timestamp 1
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_167
timestamp 1
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_168
timestamp 1
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_169
timestamp 1
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_170
timestamp 1
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_171
timestamp 1
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_172
timestamp 1
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_173
timestamp 1
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_174
timestamp 1
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_175
timestamp 1
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_176
timestamp 1
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_177
timestamp 1
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_178
timestamp 1
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_179
timestamp 1
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_180
timestamp 1
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_181
timestamp 1
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_182
timestamp 1
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_183
timestamp 1
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_184
timestamp 1
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_185
timestamp 1
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_186
timestamp 1
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_187
timestamp 1
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_188
timestamp 1
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_189
timestamp 1
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_190
timestamp 1
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_191
timestamp 1
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_192
timestamp 1
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_193
timestamp 1
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_194
timestamp 1
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_195
timestamp 1
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_196
timestamp 1
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_197
timestamp 1
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_198
timestamp 1
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_199
timestamp 1
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_200
timestamp 1
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_201
timestamp 1
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_202
timestamp 1
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_203
timestamp 1
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_204
timestamp 1
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_205
timestamp 1
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_206
timestamp 1
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_207
timestamp 1
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_208
timestamp 1
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_209
timestamp 1
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_210
timestamp 1
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_211
timestamp 1
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_212
timestamp 1
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_213
timestamp 1
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_214
timestamp 1
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_215
timestamp 1
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_216
timestamp 1
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_217
timestamp 1
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_218
timestamp 1
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_219
timestamp 1
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_220
timestamp 1
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_221
timestamp 1
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_222
timestamp 1
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_223
timestamp 1
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_224
timestamp 1
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_225
timestamp 1
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_226
timestamp 1
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_227
timestamp 1
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_228
timestamp 1
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_229
timestamp 1
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_230
timestamp 1
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_231
timestamp 1
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_232
timestamp 1
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_233
timestamp 1
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_234
timestamp 1
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_235
timestamp 1
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_236
timestamp 1
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_237
timestamp 1
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_238
timestamp 1
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_239
timestamp 1
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_240
timestamp 1
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_241
timestamp 1
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_242
timestamp 1
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_243
timestamp 1
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_244
timestamp 1
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_245
timestamp 1
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_246
timestamp 1
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_247
timestamp 1
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_248
timestamp 1
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_249
timestamp 1
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_250
timestamp 1
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_251
timestamp 1
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_252
timestamp 1
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_253
timestamp 1
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_254
timestamp 1
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_255
timestamp 1
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_256
timestamp 1
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_257
timestamp 1
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_258
timestamp 1
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_259
timestamp 1
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_260
timestamp 1
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_261
timestamp 1
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_262
timestamp 1
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_263
timestamp 1
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_264
timestamp 1
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_265
timestamp 1
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_266
timestamp 1
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_267
timestamp 1
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_268
timestamp 1
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_269
timestamp 1
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_270
timestamp 1
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_271
timestamp 1
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_272
timestamp 1
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_273
timestamp 1
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_274
timestamp 1
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_275
timestamp 1
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_276
timestamp 1
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_277
timestamp 1
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_278
timestamp 1
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_279
timestamp 1
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_280
timestamp 1
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_281
timestamp 1
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_282
timestamp 1
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_283
timestamp 1
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_284
timestamp 1
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_285
timestamp 1
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_286
timestamp 1
transform 1 0 3680 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_287
timestamp 1
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_288
timestamp 1
transform 1 0 8832 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_289
timestamp 1
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_290
timestamp 1
transform 1 0 13984 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_291
timestamp 1
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_292
timestamp 1
transform 1 0 19136 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_293
timestamp 1
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_294
timestamp 1
transform 1 0 24288 0 -1 26112
box -38 -48 130 592
<< labels >>
flabel metal4 s 4868 2128 5188 26160 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4208 2128 4528 26160 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 13542 27669 13598 28469 0 FreeSans 224 90 0 0 bit_period[0]
port 2 nsew signal input
flabel metal2 s 12898 27669 12954 28469 0 FreeSans 224 90 0 0 bit_period[10]
port 3 nsew signal input
flabel metal2 s 15474 27669 15530 28469 0 FreeSans 224 90 0 0 bit_period[11]
port 4 nsew signal input
flabel metal2 s 16118 27669 16174 28469 0 FreeSans 224 90 0 0 bit_period[12]
port 5 nsew signal input
flabel metal2 s 14830 27669 14886 28469 0 FreeSans 224 90 0 0 bit_period[13]
port 6 nsew signal input
flabel metal2 s 12254 27669 12310 28469 0 FreeSans 224 90 0 0 bit_period[1]
port 7 nsew signal input
flabel metal2 s 9034 27669 9090 28469 0 FreeSans 224 90 0 0 bit_period[2]
port 8 nsew signal input
flabel metal2 s 11610 27669 11666 28469 0 FreeSans 224 90 0 0 bit_period[3]
port 9 nsew signal input
flabel metal2 s 14186 27669 14242 28469 0 FreeSans 224 90 0 0 bit_period[4]
port 10 nsew signal input
flabel metal2 s 10322 27669 10378 28469 0 FreeSans 224 90 0 0 bit_period[5]
port 11 nsew signal input
flabel metal2 s 10966 27669 11022 28469 0 FreeSans 224 90 0 0 bit_period[6]
port 12 nsew signal input
flabel metal2 s 18050 27669 18106 28469 0 FreeSans 224 90 0 0 bit_period[7]
port 13 nsew signal input
flabel metal2 s 9678 27669 9734 28469 0 FreeSans 224 90 0 0 bit_period[8]
port 14 nsew signal input
flabel metal2 s 17406 27669 17462 28469 0 FreeSans 224 90 0 0 bit_period[9]
port 15 nsew signal input
flabel metal3 s 0 24488 800 24608 0 FreeSans 480 0 0 0 clk
port 16 nsew signal input
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 confirmation
port 17 nsew signal input
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 data_read
port 18 nsew signal output
flabel metal3 s 25525 3408 26325 3528 0 FreeSans 480 0 0 0 n_rst
port 19 nsew signal input
flabel metal3 s 0 14288 800 14408 0 FreeSans 480 0 0 0 serial_in
port 20 nsew signal input
flabel metal3 s 25525 12928 26325 13048 0 FreeSans 480 0 0 0 serial_out
port 21 nsew signal output
flabel metal3 s 25525 25168 26325 25288 0 FreeSans 480 0 0 0 tx_busy
port 22 nsew signal output
rlabel metal1 13156 26112 13156 26112 0 VGND
rlabel metal1 13156 25568 13156 25568 0 VPWR
rlabel metal2 21206 15640 21206 15640 0 _0000_
rlabel metal1 24472 15062 24472 15062 0 _0001_
rlabel metal1 20010 14586 20010 14586 0 _0002_
rlabel metal2 22862 12665 22862 12665 0 _0003_
rlabel metal1 23046 15674 23046 15674 0 _0004_
rlabel metal2 7866 16252 7866 16252 0 _0005_
rlabel metal2 7866 15130 7866 15130 0 _0006_
rlabel metal2 7222 13532 7222 13532 0 _0007_
rlabel metal1 5888 11186 5888 11186 0 _0008_
rlabel metal2 6762 13260 6762 13260 0 _0009_
rlabel metal1 4784 11730 4784 11730 0 _0010_
rlabel metal1 4140 12614 4140 12614 0 _0011_
rlabel metal2 3634 15164 3634 15164 0 _0012_
rlabel metal1 1932 11866 1932 11866 0 _0013_
rlabel metal1 1748 11050 1748 11050 0 _0014_
rlabel metal1 16652 9690 16652 9690 0 _0015_
rlabel metal2 17158 11050 17158 11050 0 _0016_
rlabel metal1 14490 7514 14490 7514 0 _0017_
rlabel metal1 17894 7378 17894 7378 0 _0018_
rlabel metal1 19918 5746 19918 5746 0 _0019_
rlabel metal1 20102 6426 20102 6426 0 _0020_
rlabel metal1 16836 6222 16836 6222 0 _0021_
rlabel metal1 17342 5882 17342 5882 0 _0022_
rlabel metal2 3726 18462 3726 18462 0 _0023_
rlabel metal1 8004 8874 8004 8874 0 _0024_
rlabel metal2 3266 5984 3266 5984 0 _0025_
rlabel metal2 6578 5916 6578 5916 0 _0026_
rlabel metal1 3956 5270 3956 5270 0 _0027_
rlabel metal2 1702 6494 1702 6494 0 _0028_
rlabel metal2 10166 15708 10166 15708 0 _0029_
rlabel metal1 9752 14994 9752 14994 0 _0030_
rlabel metal1 8740 13498 8740 13498 0 _0031_
rlabel metal1 7912 9418 7912 9418 0 _0032_
rlabel metal1 9890 14042 9890 14042 0 _0033_
rlabel metal1 9246 12274 9246 12274 0 _0034_
rlabel metal2 9798 11492 9798 11492 0 _0035_
rlabel metal2 7314 11356 7314 11356 0 _0036_
rlabel metal1 10718 9486 10718 9486 0 _0037_
rlabel metal2 9338 9180 9338 9180 0 _0038_
rlabel metal2 8326 6188 8326 6188 0 _0039_
rlabel metal2 8142 6460 8142 6460 0 _0040_
rlabel metal1 10534 9010 10534 9010 0 _0041_
rlabel metal2 7406 8636 7406 8636 0 _0042_
rlabel metal1 9706 6834 9706 6834 0 _0043_
rlabel metal2 7314 6154 7314 6154 0 _0044_
rlabel metal1 16100 12274 16100 12274 0 _0045_
rlabel metal2 15042 12988 15042 12988 0 _0046_
rlabel metal1 16054 15130 16054 15130 0 _0047_
rlabel metal2 17342 14756 17342 14756 0 _0048_
rlabel metal1 17710 9486 17710 9486 0 _0049_
rlabel metal2 17066 8772 17066 8772 0 _0050_
rlabel metal2 13938 9758 13938 9758 0 _0051_
rlabel metal1 15456 8942 15456 8942 0 _0052_
rlabel metal1 6072 16218 6072 16218 0 _0053_
rlabel metal2 5382 15708 5382 15708 0 _0054_
rlabel metal2 6486 14620 6486 14620 0 _0055_
rlabel metal1 5428 13362 5428 13362 0 _0056_
rlabel metal2 4462 14076 4462 14076 0 _0057_
rlabel metal2 2346 13668 2346 13668 0 _0058_
rlabel metal2 1794 14620 1794 14620 0 _0059_
rlabel metal2 2070 15674 2070 15674 0 _0060_
rlabel metal2 1794 16796 1794 16796 0 _0061_
rlabel metal1 3634 23732 3634 23732 0 _0062_
rlabel metal1 2990 10030 2990 10030 0 _0063_
rlabel metal1 18262 21964 18262 21964 0 _0064_
rlabel metal2 22034 21063 22034 21063 0 _0065_
rlabel metal1 13018 21556 13018 21556 0 _0066_
rlabel metal1 9706 22508 9706 22508 0 _0067_
rlabel metal1 12972 21998 12972 21998 0 _0068_
rlabel metal1 17250 23562 17250 23562 0 _0069_
rlabel metal1 18584 21658 18584 21658 0 _0070_
rlabel via2 13386 24157 13386 24157 0 _0071_
rlabel metal1 17434 5712 17434 5712 0 _0072_
rlabel metal2 4830 25466 4830 25466 0 _0073_
rlabel metal1 4922 24106 4922 24106 0 _0074_
rlabel metal1 5566 23698 5566 23698 0 _0075_
rlabel metal1 5106 23562 5106 23562 0 _0076_
rlabel metal2 3450 23902 3450 23902 0 _0077_
rlabel metal1 3082 24208 3082 24208 0 _0078_
rlabel metal1 6440 7990 6440 7990 0 _0079_
rlabel metal1 2714 7990 2714 7990 0 _0080_
rlabel metal2 4462 8687 4462 8687 0 _0081_
rlabel metal1 5244 8942 5244 8942 0 _0082_
rlabel metal1 9154 15606 9154 15606 0 _0083_
rlabel metal1 4554 7412 4554 7412 0 _0084_
rlabel metal1 4140 9554 4140 9554 0 _0085_
rlabel metal2 4278 7327 4278 7327 0 _0086_
rlabel metal1 7406 6834 7406 6834 0 _0087_
rlabel metal1 6670 7888 6670 7888 0 _0088_
rlabel metal2 3358 11900 3358 11900 0 _0089_
rlabel metal1 2162 23630 2162 23630 0 _0090_
rlabel metal2 4738 25670 4738 25670 0 _0091_
rlabel metal1 10902 21998 10902 21998 0 _0092_
rlabel metal1 12190 23698 12190 23698 0 _0093_
rlabel metal2 11086 23868 11086 23868 0 _0094_
rlabel metal1 8878 21658 8878 21658 0 _0095_
rlabel metal1 9568 21590 9568 21590 0 _0096_
rlabel metal2 13018 23494 13018 23494 0 _0097_
rlabel metal1 12512 22474 12512 22474 0 _0098_
rlabel metal2 11270 23392 11270 23392 0 _0099_
rlabel metal2 11822 23868 11822 23868 0 _0100_
rlabel metal1 8648 22202 8648 22202 0 _0101_
rlabel metal2 9062 23052 9062 23052 0 _0102_
rlabel metal2 11086 23426 11086 23426 0 _0103_
rlabel metal2 9154 22780 9154 22780 0 _0104_
rlabel metal1 12696 22066 12696 22066 0 _0105_
rlabel metal1 10856 19958 10856 19958 0 _0106_
rlabel metal2 12282 22134 12282 22134 0 _0107_
rlabel metal1 12098 22066 12098 22066 0 _0108_
rlabel metal2 6578 21692 6578 21692 0 _0109_
rlabel metal1 10764 23154 10764 23154 0 _0110_
rlabel metal1 10488 23086 10488 23086 0 _0111_
rlabel metal1 9522 22678 9522 22678 0 _0112_
rlabel metal1 10120 22746 10120 22746 0 _0113_
rlabel metal1 7360 21998 7360 21998 0 _0114_
rlabel metal2 5658 21692 5658 21692 0 _0115_
rlabel metal1 2530 20502 2530 20502 0 _0116_
rlabel metal1 5290 21590 5290 21590 0 _0117_
rlabel metal1 5888 21386 5888 21386 0 _0118_
rlabel metal1 7774 22066 7774 22066 0 _0119_
rlabel metal1 8510 24378 8510 24378 0 _0120_
rlabel metal1 8740 24582 8740 24582 0 _0121_
rlabel metal1 7222 24072 7222 24072 0 _0122_
rlabel metal1 8878 24310 8878 24310 0 _0123_
rlabel metal1 7176 20298 7176 20298 0 _0124_
rlabel metal1 7544 23290 7544 23290 0 _0125_
rlabel metal1 7820 18326 7820 18326 0 _0126_
rlabel metal2 6210 19924 6210 19924 0 _0127_
rlabel metal2 7682 19720 7682 19720 0 _0128_
rlabel metal1 7360 18394 7360 18394 0 _0129_
rlabel metal1 9246 19686 9246 19686 0 _0130_
rlabel metal1 9614 18700 9614 18700 0 _0131_
rlabel metal1 12696 18054 12696 18054 0 _0132_
rlabel viali 13110 18257 13110 18257 0 _0133_
rlabel metal1 12420 18394 12420 18394 0 _0134_
rlabel metal1 13087 18122 13087 18122 0 _0135_
rlabel metal2 10994 18496 10994 18496 0 _0136_
rlabel metal2 12742 20774 12742 20774 0 _0137_
rlabel metal1 12612 19482 12612 19482 0 _0138_
rlabel metal2 13478 20230 13478 20230 0 _0139_
rlabel metal1 13202 20502 13202 20502 0 _0140_
rlabel metal1 13524 20570 13524 20570 0 _0141_
rlabel metal1 14063 22746 14063 22746 0 _0142_
rlabel metal1 12742 23834 12742 23834 0 _0143_
rlabel metal1 14030 24106 14030 24106 0 _0144_
rlabel metal1 13754 22542 13754 22542 0 _0145_
rlabel metal1 14122 22406 14122 22406 0 _0146_
rlabel metal1 13846 21964 13846 21964 0 _0147_
rlabel metal1 10396 19278 10396 19278 0 _0148_
rlabel metal1 8280 20366 8280 20366 0 _0149_
rlabel metal2 9706 21488 9706 21488 0 _0150_
rlabel metal1 8280 24378 8280 24378 0 _0151_
rlabel metal2 7314 21182 7314 21182 0 _0152_
rlabel metal2 13570 24650 13570 24650 0 _0153_
rlabel metal1 13432 20366 13432 20366 0 _0154_
rlabel metal1 9982 20570 9982 20570 0 _0155_
rlabel metal1 8648 18870 8648 18870 0 _0156_
rlabel metal1 10304 20978 10304 20978 0 _0157_
rlabel metal1 10856 20910 10856 20910 0 _0158_
rlabel metal1 10488 21046 10488 21046 0 _0159_
rlabel metal1 10764 20978 10764 20978 0 _0160_
rlabel metal1 13662 21114 13662 21114 0 _0161_
rlabel metal2 13018 21114 13018 21114 0 _0162_
rlabel metal1 10626 21114 10626 21114 0 _0163_
rlabel metal1 13662 24208 13662 24208 0 _0164_
rlabel metal1 11086 24276 11086 24276 0 _0165_
rlabel metal1 3496 7514 3496 7514 0 _0166_
rlabel metal1 20194 15436 20194 15436 0 _0167_
rlabel metal2 4002 8058 4002 8058 0 _0168_
rlabel metal1 20470 15368 20470 15368 0 _0169_
rlabel via1 20365 15470 20365 15470 0 _0170_
rlabel metal2 19734 20128 19734 20128 0 _0171_
rlabel metal1 17250 23154 17250 23154 0 _0172_
rlabel metal1 19044 22202 19044 22202 0 _0173_
rlabel metal2 17434 22916 17434 22916 0 _0174_
rlabel metal1 18170 22134 18170 22134 0 _0175_
rlabel metal1 16468 20570 16468 20570 0 _0176_
rlabel metal1 21804 22474 21804 22474 0 _0177_
rlabel metal2 17986 22576 17986 22576 0 _0178_
rlabel metal1 16284 21046 16284 21046 0 _0179_
rlabel metal2 21022 21148 21022 21148 0 _0180_
rlabel metal1 19826 20298 19826 20298 0 _0181_
rlabel metal1 19090 23290 19090 23290 0 _0182_
rlabel metal1 15686 22066 15686 22066 0 _0183_
rlabel metal1 22126 21658 22126 21658 0 _0184_
rlabel metal1 21160 21046 21160 21046 0 _0185_
rlabel metal1 17986 21454 17986 21454 0 _0186_
rlabel metal1 21022 20366 21022 20366 0 _0187_
rlabel metal2 18354 22508 18354 22508 0 _0188_
rlabel metal1 17158 20570 17158 20570 0 _0189_
rlabel metal1 18262 21556 18262 21556 0 _0190_
rlabel metal1 16836 19890 16836 19890 0 _0191_
rlabel metal1 15824 21658 15824 21658 0 _0192_
rlabel metal1 20332 20570 20332 20570 0 _0193_
rlabel metal1 20608 21318 20608 21318 0 _0194_
rlabel metal1 19688 21522 19688 21522 0 _0195_
rlabel metal2 19274 21114 19274 21114 0 _0196_
rlabel metal2 17986 21828 17986 21828 0 _0197_
rlabel metal2 17158 22576 17158 22576 0 _0198_
rlabel metal1 17526 22066 17526 22066 0 _0199_
rlabel metal1 17112 22134 17112 22134 0 _0200_
rlabel metal2 19090 21352 19090 21352 0 _0201_
rlabel metal1 18906 20468 18906 20468 0 _0202_
rlabel metal1 19688 20774 19688 20774 0 _0203_
rlabel metal1 16054 16966 16054 16966 0 _0204_
rlabel metal1 16782 17306 16782 17306 0 _0205_
rlabel metal2 15870 18904 15870 18904 0 _0206_
rlabel metal1 15502 18904 15502 18904 0 _0207_
rlabel metal2 20654 19074 20654 19074 0 _0208_
rlabel metal2 16882 18224 16882 18224 0 _0209_
rlabel metal2 18998 18394 18998 18394 0 _0210_
rlabel metal1 18860 17850 18860 17850 0 _0211_
rlabel metal1 20930 18870 20930 18870 0 _0212_
rlabel metal2 20930 19040 20930 19040 0 _0213_
rlabel metal1 22808 22746 22808 22746 0 _0214_
rlabel metal1 22034 19176 22034 19176 0 _0215_
rlabel metal1 23230 20944 23230 20944 0 _0216_
rlabel metal1 22540 21862 22540 21862 0 _0217_
rlabel metal1 22402 23698 22402 23698 0 _0218_
rlabel metal1 22356 23834 22356 23834 0 _0219_
rlabel metal1 22862 23834 22862 23834 0 _0220_
rlabel metal2 20930 23902 20930 23902 0 _0221_
rlabel metal1 21160 24174 21160 24174 0 _0222_
rlabel metal2 19918 23902 19918 23902 0 _0223_
rlabel metal1 20148 23766 20148 23766 0 _0224_
rlabel metal1 19182 24752 19182 24752 0 _0225_
rlabel metal1 17388 24310 17388 24310 0 _0226_
rlabel metal1 19642 23562 19642 23562 0 _0227_
rlabel metal1 17572 24378 17572 24378 0 _0228_
rlabel metal1 16238 24582 16238 24582 0 _0229_
rlabel metal1 19458 23766 19458 23766 0 _0230_
rlabel metal2 21022 19754 21022 19754 0 _0231_
rlabel metal1 19550 18802 19550 18802 0 _0232_
rlabel metal1 19182 18938 19182 18938 0 _0233_
rlabel metal1 18998 18802 18998 18802 0 _0234_
rlabel metal1 20930 18394 20930 18394 0 _0235_
rlabel metal2 19734 19040 19734 19040 0 _0236_
rlabel metal2 20470 20944 20470 20944 0 _0237_
rlabel metal2 20010 20128 20010 20128 0 _0238_
rlabel metal2 15962 20094 15962 20094 0 _0239_
rlabel metal1 20102 19856 20102 19856 0 _0240_
rlabel metal2 19918 19516 19918 19516 0 _0241_
rlabel metal2 19550 20781 19550 20781 0 _0242_
rlabel metal2 19642 23902 19642 23902 0 _0243_
rlabel metal1 19642 24208 19642 24208 0 _0244_
rlabel metal1 17204 24174 17204 24174 0 _0245_
rlabel metal2 17250 24582 17250 24582 0 _0246_
rlabel metal2 19734 24225 19734 24225 0 _0247_
rlabel metal2 21942 14586 21942 14586 0 _0248_
rlabel metal1 21712 14790 21712 14790 0 _0249_
rlabel metal1 21528 14314 21528 14314 0 _0250_
rlabel metal1 21896 14586 21896 14586 0 _0251_
rlabel metal1 20654 9554 20654 9554 0 _0252_
rlabel metal1 20332 9554 20332 9554 0 _0253_
rlabel metal1 20700 9146 20700 9146 0 _0254_
rlabel metal1 20056 11118 20056 11118 0 _0255_
rlabel metal1 19964 9690 19964 9690 0 _0256_
rlabel metal1 20378 10064 20378 10064 0 _0257_
rlabel metal1 18216 12614 18216 12614 0 _0258_
rlabel metal1 17526 12682 17526 12682 0 _0259_
rlabel metal1 18814 12818 18814 12818 0 _0260_
rlabel metal1 17480 12614 17480 12614 0 _0261_
rlabel metal1 17756 12410 17756 12410 0 _0262_
rlabel metal1 18400 13362 18400 13362 0 _0263_
rlabel metal1 18868 11798 18868 11798 0 _0264_
rlabel metal2 19090 12036 19090 12036 0 _0265_
rlabel metal1 18538 12240 18538 12240 0 _0266_
rlabel metal1 20010 12172 20010 12172 0 _0267_
rlabel metal1 20424 9418 20424 9418 0 _0268_
rlabel metal1 21712 9350 21712 9350 0 _0269_
rlabel metal2 21206 9180 21206 9180 0 _0270_
rlabel metal2 22678 9826 22678 9826 0 _0271_
rlabel metal1 20240 9078 20240 9078 0 _0272_
rlabel metal2 24334 12988 24334 12988 0 _0273_
rlabel metal1 24242 12852 24242 12852 0 _0274_
rlabel via1 22586 12817 22586 12817 0 _0275_
rlabel metal1 22218 10166 22218 10166 0 _0276_
rlabel metal2 23414 11628 23414 11628 0 _0277_
rlabel metal1 21482 9010 21482 9010 0 _0278_
rlabel metal2 22494 9860 22494 9860 0 _0279_
rlabel metal1 22356 10778 22356 10778 0 _0280_
rlabel metal2 22218 13124 22218 13124 0 _0281_
rlabel metal1 19734 11866 19734 11866 0 _0282_
rlabel metal2 22126 11866 22126 11866 0 _0283_
rlabel metal2 21942 11526 21942 11526 0 _0284_
rlabel metal2 22770 13889 22770 13889 0 _0285_
rlabel metal2 23322 14960 23322 14960 0 _0286_
rlabel metal1 21482 11084 21482 11084 0 _0287_
rlabel metal2 21574 10948 21574 10948 0 _0288_
rlabel metal1 22264 9418 22264 9418 0 _0289_
rlabel metal1 20516 11322 20516 11322 0 _0290_
rlabel metal1 21022 13158 21022 13158 0 _0291_
rlabel metal2 20470 11594 20470 11594 0 _0292_
rlabel metal1 20102 11322 20102 11322 0 _0293_
rlabel metal1 23276 13838 23276 13838 0 _0294_
rlabel metal1 21390 13294 21390 13294 0 _0295_
rlabel metal2 21942 12138 21942 12138 0 _0296_
rlabel metal1 22586 12682 22586 12682 0 _0297_
rlabel metal1 22264 13702 22264 13702 0 _0298_
rlabel metal1 21896 13498 21896 13498 0 _0299_
rlabel metal1 21206 12852 21206 12852 0 _0300_
rlabel metal1 18952 12342 18952 12342 0 _0301_
rlabel metal1 18584 12410 18584 12410 0 _0302_
rlabel metal1 20332 12682 20332 12682 0 _0303_
rlabel metal1 20562 11866 20562 11866 0 _0304_
rlabel metal2 18354 13226 18354 13226 0 _0305_
rlabel metal1 18630 12818 18630 12818 0 _0306_
rlabel metal1 19366 12784 19366 12784 0 _0307_
rlabel metal1 19964 12614 19964 12614 0 _0308_
rlabel metal2 21390 11356 21390 11356 0 _0309_
rlabel metal2 22218 11492 22218 11492 0 _0310_
rlabel metal1 3036 18734 3036 18734 0 _0311_
rlabel metal1 2691 19142 2691 19142 0 _0312_
rlabel via1 2806 19958 2806 19958 0 _0313_
rlabel metal2 2898 19958 2898 19958 0 _0314_
rlabel metal2 3634 20026 3634 20026 0 _0315_
rlabel metal2 22310 16252 22310 16252 0 _0316_
rlabel metal2 21114 16048 21114 16048 0 _0317_
rlabel metal2 20654 15674 20654 15674 0 _0318_
rlabel metal1 20930 15334 20930 15334 0 _0319_
rlabel metal1 21758 12954 21758 12954 0 _0320_
rlabel metal1 4876 19754 4876 19754 0 _0321_
rlabel metal2 1610 11322 1610 11322 0 _0322_
rlabel via2 3266 8483 3266 8483 0 _0323_
rlabel metal2 6762 7582 6762 7582 0 _0324_
rlabel metal1 5382 6630 5382 6630 0 _0325_
rlabel metal1 15364 8466 15364 8466 0 _0326_
rlabel metal2 12926 9112 12926 9112 0 _0327_
rlabel metal1 13110 7820 13110 7820 0 _0328_
rlabel metal1 13478 8976 13478 8976 0 _0329_
rlabel metal1 15226 8806 15226 8806 0 _0330_
rlabel metal1 12098 7344 12098 7344 0 _0331_
rlabel metal2 12282 7718 12282 7718 0 _0332_
rlabel metal1 12742 7378 12742 7378 0 _0333_
rlabel metal1 13202 7956 13202 7956 0 _0334_
rlabel metal2 13294 7684 13294 7684 0 _0335_
rlabel metal1 13202 7344 13202 7344 0 _0336_
rlabel metal1 14030 7378 14030 7378 0 _0337_
rlabel metal2 11730 5882 11730 5882 0 _0338_
rlabel metal1 12535 5610 12535 5610 0 _0339_
rlabel metal2 11914 5338 11914 5338 0 _0340_
rlabel metal1 12006 5746 12006 5746 0 _0341_
rlabel metal1 13018 5576 13018 5576 0 _0342_
rlabel metal1 13708 6358 13708 6358 0 _0343_
rlabel metal1 13478 5882 13478 5882 0 _0344_
rlabel metal1 12926 7310 12926 7310 0 _0345_
rlabel metal2 13754 6766 13754 6766 0 _0346_
rlabel metal1 13478 6256 13478 6256 0 _0347_
rlabel metal2 15686 6562 15686 6562 0 _0348_
rlabel metal1 16606 6834 16606 6834 0 _0349_
rlabel metal2 16974 7174 16974 7174 0 _0350_
rlabel metal2 13386 4556 13386 4556 0 _0351_
rlabel metal1 13892 4114 13892 4114 0 _0352_
rlabel metal1 13662 4114 13662 4114 0 _0353_
rlabel metal1 14168 3706 14168 3706 0 _0354_
rlabel metal1 14996 3910 14996 3910 0 _0355_
rlabel metal2 12926 4794 12926 4794 0 _0356_
rlabel metal1 13156 4658 13156 4658 0 _0357_
rlabel metal1 15272 4182 15272 4182 0 _0358_
rlabel metal1 15226 4114 15226 4114 0 _0359_
rlabel metal1 15916 4114 15916 4114 0 _0360_
rlabel metal1 17480 4114 17480 4114 0 _0361_
rlabel metal1 15640 6290 15640 6290 0 _0362_
rlabel metal1 14214 3978 14214 3978 0 _0363_
rlabel metal1 15364 5542 15364 5542 0 _0364_
rlabel metal1 15318 5644 15318 5644 0 _0365_
rlabel metal1 16376 5338 16376 5338 0 _0366_
rlabel metal1 17756 5542 17756 5542 0 _0367_
rlabel metal1 16284 5882 16284 5882 0 _0368_
rlabel metal1 16008 5542 16008 5542 0 _0369_
rlabel metal1 16054 6256 16054 6256 0 _0370_
rlabel metal1 3082 18394 3082 18394 0 _0371_
rlabel metal1 6578 9962 6578 9962 0 _0372_
rlabel metal2 4370 9894 4370 9894 0 _0373_
rlabel metal1 2852 9622 2852 9622 0 _0374_
rlabel metal2 3358 10234 3358 10234 0 _0375_
rlabel metal1 2990 8058 2990 8058 0 _0376_
rlabel metal1 2346 9996 2346 9996 0 _0377_
rlabel metal1 2852 9894 2852 9894 0 _0378_
rlabel metal1 2346 6834 2346 6834 0 _0379_
rlabel metal2 5934 9112 5934 9112 0 _0380_
rlabel metal1 4370 7344 4370 7344 0 _0381_
rlabel metal1 4646 8602 4646 8602 0 _0382_
rlabel metal1 15318 14416 15318 14416 0 _0383_
rlabel metal1 16284 14994 16284 14994 0 _0384_
rlabel metal1 5842 7412 5842 7412 0 _0385_
rlabel metal1 5988 8806 5988 8806 0 _0386_
rlabel metal2 6302 9316 6302 9316 0 _0387_
rlabel metal2 3266 8126 3266 8126 0 _0388_
rlabel metal2 3358 8704 3358 8704 0 _0389_
rlabel metal1 4692 6970 4692 6970 0 _0390_
rlabel metal1 4278 7514 4278 7514 0 _0391_
rlabel metal1 3358 7820 3358 7820 0 _0392_
rlabel metal1 2806 8500 2806 8500 0 _0393_
rlabel metal1 4462 8942 4462 8942 0 _0394_
rlabel metal1 3726 6426 3726 6426 0 _0395_
rlabel metal2 5934 7548 5934 7548 0 _0396_
rlabel metal1 6394 6426 6394 6426 0 _0397_
rlabel metal2 2530 8636 2530 8636 0 _0398_
rlabel metal1 2300 6766 2300 6766 0 _0399_
rlabel metal1 17158 13260 17158 13260 0 _0400_
rlabel metal2 14858 15844 14858 15844 0 _0401_
rlabel metal1 15234 14246 15234 14246 0 _0402_
rlabel metal2 15778 13770 15778 13770 0 _0403_
rlabel metal2 14122 14994 14122 14994 0 _0404_
rlabel metal1 13202 15878 13202 15878 0 _0405_
rlabel metal1 14076 15538 14076 15538 0 _0406_
rlabel metal1 14950 15980 14950 15980 0 _0407_
rlabel metal1 15042 16150 15042 16150 0 _0408_
rlabel metal2 15778 15300 15778 15300 0 _0409_
rlabel metal2 16054 15470 16054 15470 0 _0410_
rlabel metal1 12374 14348 12374 14348 0 _0411_
rlabel metal1 11822 13906 11822 13906 0 _0412_
rlabel metal2 12098 14688 12098 14688 0 _0413_
rlabel metal2 12466 14620 12466 14620 0 _0414_
rlabel metal1 13294 13974 13294 13974 0 _0415_
rlabel metal2 15502 14518 15502 14518 0 _0416_
rlabel metal2 14950 14790 14950 14790 0 _0417_
rlabel metal1 15640 15130 15640 15130 0 _0418_
rlabel metal1 14858 15538 14858 15538 0 _0419_
rlabel metal2 15410 15810 15410 15810 0 _0420_
rlabel metal2 17802 15164 17802 15164 0 _0421_
rlabel metal2 12190 12410 12190 12410 0 _0422_
rlabel metal2 12374 12036 12374 12036 0 _0423_
rlabel metal2 12834 12002 12834 12002 0 _0424_
rlabel metal2 12282 12070 12282 12070 0 _0425_
rlabel metal1 13064 12138 13064 12138 0 _0426_
rlabel metal1 12374 13872 12374 13872 0 _0427_
rlabel metal1 13018 13838 13018 13838 0 _0428_
rlabel metal1 13202 13770 13202 13770 0 _0429_
rlabel metal1 13524 11662 13524 11662 0 _0430_
rlabel metal2 13938 11900 13938 11900 0 _0431_
rlabel metal1 18262 10098 18262 10098 0 _0432_
rlabel metal2 13386 10880 13386 10880 0 _0433_
rlabel via1 13293 10642 13293 10642 0 _0434_
rlabel metal2 13570 10234 13570 10234 0 _0435_
rlabel metal2 12742 11866 12742 11866 0 _0436_
rlabel metal2 13478 11118 13478 11118 0 _0437_
rlabel metal1 16790 8534 16790 8534 0 _0438_
rlabel metal1 14490 10064 14490 10064 0 _0439_
rlabel metal1 14812 10438 14812 10438 0 _0440_
rlabel metal1 14260 10030 14260 10030 0 _0441_
rlabel metal2 13754 26877 13754 26877 0 bit_period[0]
rlabel metal2 13018 26843 13018 26843 0 bit_period[10]
rlabel metal2 15594 26843 15594 26843 0 bit_period[11]
rlabel metal2 16238 26843 16238 26843 0 bit_period[12]
rlabel metal2 15042 26877 15042 26877 0 bit_period[13]
rlabel metal2 12374 26877 12374 26877 0 bit_period[1]
rlabel metal2 9246 26877 9246 26877 0 bit_period[2]
rlabel metal2 11730 26843 11730 26843 0 bit_period[3]
rlabel metal2 14398 26877 14398 26877 0 bit_period[4]
rlabel metal2 10534 26877 10534 26877 0 bit_period[5]
rlabel metal1 11086 25874 11086 25874 0 bit_period[6]
rlabel metal2 18262 26877 18262 26877 0 bit_period[7]
rlabel metal2 9890 26877 9890 26877 0 bit_period[8]
rlabel metal2 17618 26877 17618 26877 0 bit_period[9]
rlabel metal1 12926 15096 12926 15096 0 clk
rlabel metal1 18308 20910 18308 20910 0 clknet_0_clk
rlabel metal1 1840 13906 1840 13906 0 clknet_3_0__leaf_clk
rlabel metal2 8142 14144 8142 14144 0 clknet_3_1__leaf_clk
rlabel metal2 1426 20434 1426 20434 0 clknet_3_2__leaf_clk
rlabel metal1 7452 20978 7452 20978 0 clknet_3_3__leaf_clk
rlabel metal1 16790 14926 16790 14926 0 clknet_3_4__leaf_clk
rlabel metal1 21390 15538 21390 15538 0 clknet_3_5__leaf_clk
rlabel metal2 13938 18768 13938 18768 0 clknet_3_6__leaf_clk
rlabel metal1 23322 24106 23322 24106 0 clknet_3_7__leaf_clk
rlabel metal1 3312 11662 3312 11662 0 cntrl.data_ready
rlabel metal2 2254 18938 2254 18938 0 cntrl.framing_error
rlabel metal1 3220 9010 3220 9010 0 cntrl.overrun_error
rlabel metal2 4738 8517 4738 8517 0 cntrl.state\[0\]
rlabel metal1 3680 6222 3680 6222 0 cntrl.state\[1\]
rlabel metal1 5842 6732 5842 6732 0 cntrl.state\[2\]
rlabel metal2 5290 6086 5290 6086 0 cntrl.state\[3\]
rlabel metal1 3818 6766 3818 6766 0 cntrl.state\[4\]
rlabel metal3 1050 15028 1050 15028 0 confirmation
rlabel metal3 751 11628 751 11628 0 data_read
rlabel via2 24886 3485 24886 3485 0 n_rst
rlabel viali 16238 19822 16238 19822 0 net1
rlabel metal1 19918 20910 19918 20910 0 net10
rlabel metal2 11086 25466 11086 25466 0 net11
rlabel metal1 21942 21352 21942 21352 0 net12
rlabel metal2 19964 21692 19964 21692 0 net13
rlabel metal1 17572 25670 17572 25670 0 net14
rlabel metal1 2300 15334 2300 15334 0 net15
rlabel metal2 21390 6766 21390 6766 0 net16
rlabel metal1 1702 14042 1702 14042 0 net17
rlabel metal1 1426 11220 1426 11220 0 net18
rlabel metal1 23506 11866 23506 11866 0 net19
rlabel metal1 13570 20910 13570 20910 0 net2
rlabel metal2 22448 22202 22448 22202 0 net20
rlabel metal2 14122 22950 14122 22950 0 net21
rlabel metal1 18584 5746 18584 5746 0 net22
rlabel metal2 4002 10370 4002 10370 0 net23
rlabel metal2 21574 12857 21574 12857 0 net24
rlabel metal2 3450 17153 3450 17153 0 net25
rlabel metal1 6171 12138 6171 12138 0 net26
rlabel metal1 6302 13267 6302 13267 0 net27
rlabel metal2 8234 13634 8234 13634 0 net28
rlabel metal2 8326 10880 8326 10880 0 net29
rlabel metal2 17802 25262 17802 25262 0 net3
rlabel metal1 3089 19822 3089 19822 0 net30
rlabel metal2 6118 17714 6118 17714 0 net31
rlabel metal2 10120 18258 10120 18258 0 net32
rlabel metal1 11185 17170 11185 17170 0 net33
rlabel metal1 11408 15470 11408 15470 0 net34
rlabel metal1 18584 6358 18584 6358 0 net35
rlabel metal1 19182 15062 19182 15062 0 net36
rlabel metal1 19734 18326 19734 18326 0 net37
rlabel metal1 17625 15402 17625 15402 0 net38
rlabel metal1 18262 15504 18262 15504 0 net39
rlabel metal2 16974 24684 16974 24684 0 net4
rlabel via2 24886 25245 24886 25245 0 net40
rlabel metal2 4186 17340 4186 17340 0 net41
rlabel metal2 5382 18564 5382 18564 0 net42
rlabel metal1 2254 11798 2254 11798 0 net43
rlabel metal1 5152 24174 5152 24174 0 net44
rlabel metal1 17434 6732 17434 6732 0 net45
rlabel metal1 21758 16014 21758 16014 0 net46
rlabel metal1 14950 10030 14950 10030 0 net47
rlabel metal1 1794 11662 1794 11662 0 net48
rlabel metal1 16560 6290 16560 6290 0 net49
rlabel metal1 13478 23086 13478 23086 0 net5
rlabel metal1 3726 23834 3726 23834 0 net50
rlabel metal1 2300 22678 2300 22678 0 net51
rlabel metal1 4554 25466 4554 25466 0 net52
rlabel metal1 19044 20026 19044 20026 0 net53
rlabel metal1 16100 13158 16100 13158 0 net54
rlabel metal1 2438 23732 2438 23732 0 net55
rlabel metal2 4278 6562 4278 6562 0 net56
rlabel metal1 15717 20910 15717 20910 0 net6
rlabel metal1 15548 21386 15548 21386 0 net7
rlabel metal1 15088 21998 15088 21998 0 net8
rlabel metal1 17618 20400 17618 20400 0 net9
rlabel via1 12282 15538 12282 15538 0 parallel_out1\[0\]
rlabel metal1 9338 15368 9338 15368 0 parallel_out1\[1\]
rlabel metal1 12834 14314 12834 14314 0 parallel_out1\[2\]
rlabel metal1 13519 13896 13519 13896 0 parallel_out1\[3\]
rlabel metal1 13294 14382 13294 14382 0 parallel_out1\[4\]
rlabel metal2 13018 14212 13018 14212 0 parallel_out1\[5\]
rlabel metal2 12466 15300 12466 15300 0 parallel_out1\[6\]
rlabel metal2 8694 11526 8694 11526 0 parallel_out1\[7\]
rlabel metal1 11086 5678 11086 5678 0 parallel_out2\[0\]
rlabel metal1 10074 9894 10074 9894 0 parallel_out2\[1\]
rlabel metal1 9821 5270 9821 5270 0 parallel_out2\[2\]
rlabel metal1 9016 6630 9016 6630 0 parallel_out2\[3\]
rlabel metal2 12834 6018 12834 6018 0 parallel_out2\[4\]
rlabel metal2 8878 8704 8878 8704 0 parallel_out2\[5\]
rlabel metal1 10603 6970 10603 6970 0 parallel_out2\[6\]
rlabel metal1 8142 5882 8142 5882 0 parallel_out2\[7\]
rlabel metal1 17020 12818 17020 12818 0 prod_adder.gen_for_loop\[0\].adder_n.a
rlabel metal1 17342 12886 17342 12886 0 prod_adder.gen_for_loop\[0\].adder_n.b
rlabel metal1 16583 12818 16583 12818 0 prod_adder.gen_for_loop\[1\].adder_n.a
rlabel metal1 17319 11050 17319 11050 0 prod_adder.gen_for_loop\[1\].adder_n.b
rlabel metal1 17503 15334 17503 15334 0 prod_adder.gen_for_loop\[2\].adder_n.a
rlabel metal1 18262 12852 18262 12852 0 prod_adder.gen_for_loop\[2\].adder_n.b
rlabel metal1 17894 14382 17894 14382 0 prod_adder.gen_for_loop\[3\].adder_n.a
rlabel metal1 18837 7514 18837 7514 0 prod_adder.gen_for_loop\[3\].adder_n.b
rlabel metal1 19458 9996 19458 9996 0 prod_adder.gen_for_loop\[4\].adder_n.a
rlabel metal1 18975 5678 18975 5678 0 prod_adder.gen_for_loop\[4\].adder_n.b
rlabel metal1 18101 8806 18101 8806 0 prod_adder.gen_for_loop\[5\].adder_n.a
rlabel metal1 20700 8466 20700 8466 0 prod_adder.gen_for_loop\[5\].adder_n.b
rlabel metal2 20102 9248 20102 9248 0 prod_adder.gen_for_loop\[6\].adder_n.a
rlabel metal2 19918 9282 19918 9282 0 prod_adder.gen_for_loop\[6\].adder_n.b
rlabel metal1 18101 9146 18101 9146 0 prod_adder.gen_for_loop\[7\].adder_n.a
rlabel metal2 19090 7854 19090 7854 0 prod_adder.gen_for_loop\[7\].adder_n.b
rlabel metal1 11270 16150 11270 16150 0 rx_data\[0\]
rlabel metal1 8648 15334 8648 15334 0 rx_data\[1\]
rlabel metal1 8533 13430 8533 13430 0 rx_data\[2\]
rlabel metal2 8510 8160 8510 8160 0 rx_data\[3\]
rlabel metal1 7843 12954 7843 12954 0 rx_data\[4\]
rlabel metal1 5934 12954 5934 12954 0 rx_data\[5\]
rlabel metal1 5060 12818 5060 12818 0 rx_data\[6\]
rlabel metal1 5819 14858 5819 14858 0 rx_data\[7\]
rlabel metal3 751 14348 751 14348 0 serial_in
rlabel metal2 24794 13073 24794 13073 0 serial_out
rlabel metal1 2024 20570 2024 20570 0 uart_rcv.control.next_state\[0\]
rlabel metal2 3266 20638 3266 20638 0 uart_rcv.control.next_state\[1\]
rlabel metal1 1702 19720 1702 19720 0 uart_rcv.control.next_state\[2\]
rlabel metal1 2622 20468 2622 20468 0 uart_rcv.control.packet_done
rlabel metal1 3818 20944 3818 20944 0 uart_rcv.control.state\[0\]
rlabel metal1 5566 20434 5566 20434 0 uart_rcv.control.state\[1\]
rlabel metal2 3174 19584 3174 19584 0 uart_rcv.control.state\[2\]
rlabel metal1 7659 16626 7659 16626 0 uart_rcv.data_buff.packet_data\[0\]
rlabel metal1 6348 16082 6348 16082 0 uart_rcv.data_buff.packet_data\[1\]
rlabel metal1 6716 14994 6716 14994 0 uart_rcv.data_buff.packet_data\[2\]
rlabel metal1 6647 13158 6647 13158 0 uart_rcv.data_buff.packet_data\[3\]
rlabel metal1 5221 14042 5221 14042 0 uart_rcv.data_buff.packet_data\[4\]
rlabel metal1 4692 14246 4692 14246 0 uart_rcv.data_buff.packet_data\[5\]
rlabel metal1 3013 14586 3013 14586 0 uart_rcv.data_buff.packet_data\[6\]
rlabel metal2 2898 15572 2898 15572 0 uart_rcv.data_buff.packet_data\[7\]
rlabel metal2 2898 17782 2898 17782 0 uart_rcv.sbc.stop_bit
rlabel metal1 3542 19414 3542 19414 0 uart_rcv.sbd.new_sample
rlabel metal1 3565 18938 3565 18938 0 uart_rcv.sbd.old_sample
rlabel metal1 3519 17646 3519 17646 0 uart_rcv.sbd.sync_phase
rlabel metal1 4922 23698 4922 23698 0 uart_rcv.shift_strobe
rlabel metal2 3910 23222 3910 23222 0 uart_rcv.tim.bit_cnt\[0\]
rlabel metal1 3588 24718 3588 24718 0 uart_rcv.tim.bit_cnt\[1\]
rlabel metal1 3680 25330 3680 25330 0 uart_rcv.tim.bit_cnt\[2\]
rlabel metal1 5980 24922 5980 24922 0 uart_rcv.tim.bit_cnt\[3\]
rlabel metal2 2898 23868 2898 23868 0 uart_rcv.tim.bit_count.next_cnt_out\[0\]
rlabel metal1 1932 24310 1932 24310 0 uart_rcv.tim.bit_count.next_cnt_out\[1\]
rlabel metal2 2070 25500 2070 25500 0 uart_rcv.tim.bit_count.next_cnt_out\[2\]
rlabel metal1 2530 24276 2530 24276 0 uart_rcv.tim.bit_count.next_cnt_out\[3\]
rlabel metal1 2231 23154 2231 23154 0 uart_rcv.tim.bit_count.next_roflag
rlabel metal2 8418 21828 8418 21828 0 uart_rcv.tim.clk_cnt\[0\]
rlabel metal2 12558 19686 12558 19686 0 uart_rcv.tim.clk_cnt\[10\]
rlabel metal2 12558 23018 12558 23018 0 uart_rcv.tim.clk_cnt\[11\]
rlabel metal1 15042 24922 15042 24922 0 uart_rcv.tim.clk_cnt\[12\]
rlabel metal1 13202 22678 13202 22678 0 uart_rcv.tim.clk_cnt\[13\]
rlabel metal2 10534 24650 10534 24650 0 uart_rcv.tim.clk_cnt\[1\]
rlabel metal1 7314 24378 7314 24378 0 uart_rcv.tim.clk_cnt\[2\]
rlabel metal2 7130 23222 7130 23222 0 uart_rcv.tim.clk_cnt\[3\]
rlabel metal1 8418 20536 8418 20536 0 uart_rcv.tim.clk_cnt\[4\]
rlabel metal1 7820 19686 7820 19686 0 uart_rcv.tim.clk_cnt\[5\]
rlabel metal1 9384 21318 9384 21318 0 uart_rcv.tim.clk_cnt\[6\]
rlabel metal1 13800 17850 13800 17850 0 uart_rcv.tim.clk_cnt\[7\]
rlabel metal2 12098 18292 12098 18292 0 uart_rcv.tim.clk_cnt\[8\]
rlabel metal1 11270 17306 11270 17306 0 uart_rcv.tim.clk_cnt\[9\]
rlabel metal1 6394 21454 6394 21454 0 uart_rcv.tim.clock_count.next_cnt_out\[0\]
rlabel metal1 13754 19890 13754 19890 0 uart_rcv.tim.clock_count.next_cnt_out\[10\]
rlabel metal2 12742 24956 12742 24956 0 uart_rcv.tim.clock_count.next_cnt_out\[11\]
rlabel metal2 13386 24548 13386 24548 0 uart_rcv.tim.clock_count.next_cnt_out\[12\]
rlabel metal1 13570 22066 13570 22066 0 uart_rcv.tim.clock_count.next_cnt_out\[13\]
rlabel metal1 9200 24922 9200 24922 0 uart_rcv.tim.clock_count.next_cnt_out\[1\]
rlabel via2 8234 24701 8234 24701 0 uart_rcv.tim.clock_count.next_cnt_out\[2\]
rlabel metal1 8556 22542 8556 22542 0 uart_rcv.tim.clock_count.next_cnt_out\[3\]
rlabel via1 6854 19210 6854 19210 0 uart_rcv.tim.clock_count.next_cnt_out\[4\]
rlabel metal1 6900 19890 6900 19890 0 uart_rcv.tim.clock_count.next_cnt_out\[5\]
rlabel metal2 9246 18564 9246 18564 0 uart_rcv.tim.clock_count.next_cnt_out\[6\]
rlabel metal1 12926 18054 12926 18054 0 uart_rcv.tim.clock_count.next_cnt_out\[7\]
rlabel metal2 10626 19040 10626 19040 0 uart_rcv.tim.clock_count.next_cnt_out\[8\]
rlabel metal1 9798 20978 9798 20978 0 uart_rcv.tim.clock_count.next_cnt_out\[9\]
rlabel metal1 7774 24140 7774 24140 0 uart_rcv.tim.clock_count.next_roflag
rlabel metal1 19596 18394 19596 18394 0 uart_tx.clk_cnt\[0\]
rlabel metal1 16882 24038 16882 24038 0 uart_tx.clk_cnt\[10\]
rlabel metal2 17894 23885 17894 23885 0 uart_tx.clk_cnt\[11\]
rlabel metal1 18814 21522 18814 21522 0 uart_tx.clk_cnt\[12\]
rlabel metal1 17020 22474 17020 22474 0 uart_tx.clk_cnt\[13\]
rlabel metal1 15226 20944 15226 20944 0 uart_tx.clk_cnt\[1\]
rlabel metal1 15732 20298 15732 20298 0 uart_tx.clk_cnt\[2\]
rlabel metal2 18446 21828 18446 21828 0 uart_tx.clk_cnt\[3\]
rlabel metal1 18308 17646 18308 17646 0 uart_tx.clk_cnt\[4\]
rlabel via1 20179 20910 20179 20910 0 uart_tx.clk_cnt\[5\]
rlabel metal1 21850 18632 21850 18632 0 uart_tx.clk_cnt\[6\]
rlabel metal2 23690 20740 23690 20740 0 uart_tx.clk_cnt\[7\]
rlabel metal1 22678 22406 22678 22406 0 uart_tx.clk_cnt\[8\]
rlabel metal1 22218 23800 22218 23800 0 uart_tx.clk_cnt\[9\]
rlabel metal2 18170 19346 18170 19346 0 uart_tx.count.next_cnt_out\[0\]
rlabel via2 16146 24701 16146 24701 0 uart_tx.count.next_cnt_out\[10\]
rlabel metal1 19366 24786 19366 24786 0 uart_tx.count.next_cnt_out\[11\]
rlabel metal1 19596 24378 19596 24378 0 uart_tx.count.next_cnt_out\[12\]
rlabel metal1 15778 24922 15778 24922 0 uart_tx.count.next_cnt_out\[13\]
rlabel metal1 16100 17578 16100 17578 0 uart_tx.count.next_cnt_out\[1\]
rlabel metal1 15870 18870 15870 18870 0 uart_tx.count.next_cnt_out\[2\]
rlabel via1 17066 17782 17066 17782 0 uart_tx.count.next_cnt_out\[3\]
rlabel metal1 18722 18632 18722 18632 0 uart_tx.count.next_cnt_out\[4\]
rlabel metal1 21114 18632 21114 18632 0 uart_tx.count.next_cnt_out\[5\]
rlabel metal2 22310 19142 22310 19142 0 uart_tx.count.next_cnt_out\[6\]
rlabel metal1 22954 20366 22954 20366 0 uart_tx.count.next_cnt_out\[7\]
rlabel metal1 22770 22066 22770 22066 0 uart_tx.count.next_cnt_out\[8\]
rlabel metal1 22862 24582 22862 24582 0 uart_tx.count.next_cnt_out\[9\]
rlabel metal2 20056 21556 20056 21556 0 uart_tx.count.next_roflag
rlabel metal1 20746 16048 20746 16048 0 uart_tx.count.roflag_ff
rlabel metal1 21482 14960 21482 14960 0 uart_tx.tx_ctrl.state\[0\]
rlabel metal1 22172 14994 22172 14994 0 uart_tx.tx_ctrl.state\[1\]
rlabel metal1 20930 14484 20930 14484 0 uart_tx.tx_ctrl.state\[2\]
rlabel metal2 22954 15810 22954 15810 0 uart_tx.tx_ctrl.state\[3\]
rlabel metal1 23368 15470 23368 15470 0 uart_tx.tx_ctrl.state\[4\]
<< properties >>
string FIXED_BBOX 0 0 26325 28469
<< end >>
