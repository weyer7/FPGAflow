VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sample_proj
  CLASS BLOCK ;
  FOREIGN sample_proj ;
  ORIGIN 0.000 0.000 ;
  SIZE 146.660 BY 157.380 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 144.400 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 144.400 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 142.660 23.840 146.660 24.440 ;
    END
  END clk
  PIN done
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 142.660 95.240 146.660 95.840 ;
    END
  END done
  PIN enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 142.660 30.640 146.660 31.240 ;
    END
  END enable
  PIN nrst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 142.660 27.240 146.660 27.840 ;
    END
  END nrst
  PIN out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 116.010 153.380 116.290 157.380 ;
    END
  END out[0]
  PIN out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 119.230 153.380 119.510 157.380 ;
    END
  END out[10]
  PIN out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 144.990 153.380 145.270 157.380 ;
    END
  END out[11]
  PIN out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 58.050 153.380 58.330 157.380 ;
    END
  END out[12]
  PIN out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 77.370 153.380 77.650 157.380 ;
    END
  END out[13]
  PIN out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 64.490 153.380 64.770 157.380 ;
    END
  END out[14]
  PIN out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 90.250 153.380 90.530 157.380 ;
    END
  END out[15]
  PIN out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 109.570 153.380 109.850 157.380 ;
    END
  END out[16]
  PIN out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 112.790 153.380 113.070 157.380 ;
    END
  END out[17]
  PIN out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 74.150 153.380 74.430 157.380 ;
    END
  END out[18]
  PIN out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 135.330 153.380 135.610 157.380 ;
    END
  END out[19]
  PIN out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 142.660 122.440 146.660 123.040 ;
    END
  END out[1]
  PIN out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 80.590 153.380 80.870 157.380 ;
    END
  END out[20]
  PIN out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 106.350 153.380 106.630 157.380 ;
    END
  END out[21]
  PIN out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 99.910 153.380 100.190 157.380 ;
    END
  END out[22]
  PIN out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 128.890 153.380 129.170 157.380 ;
    END
  END out[23]
  PIN out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 87.030 153.380 87.310 157.380 ;
    END
  END out[24]
  PIN out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 132.110 153.380 132.390 157.380 ;
    END
  END out[25]
  PIN out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 142.660 129.240 146.660 129.840 ;
    END
  END out[26]
  PIN out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 125.670 153.380 125.950 157.380 ;
    END
  END out[27]
  PIN out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 70.930 153.380 71.210 157.380 ;
    END
  END out[28]
  PIN out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 83.810 153.380 84.090 157.380 ;
    END
  END out[29]
  PIN out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 96.690 153.380 96.970 157.380 ;
    END
  END out[2]
  PIN out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 142.660 125.840 146.660 126.440 ;
    END
  END out[30]
  PIN out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 142.660 119.040 146.660 119.640 ;
    END
  END out[31]
  PIN out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 142.660 115.640 146.660 116.240 ;
    END
  END out[32]
  PIN out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 142.660 112.240 146.660 112.840 ;
    END
  END out[33]
  PIN out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 141.770 153.380 142.050 157.380 ;
    END
  END out[3]
  PIN out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 61.270 153.380 61.550 157.380 ;
    END
  END out[4]
  PIN out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 93.470 153.380 93.750 157.380 ;
    END
  END out[5]
  PIN out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 67.710 153.380 67.990 157.380 ;
    END
  END out[6]
  PIN out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 122.450 153.380 122.730 157.380 ;
    END
  END out[7]
  PIN out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 103.130 153.380 103.410 157.380 ;
    END
  END out[8]
  PIN out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 138.550 153.380 138.830 157.380 ;
    END
  END out[9]
  PIN prescaler[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END prescaler[0]
  PIN prescaler[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END prescaler[10]
  PIN prescaler[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END prescaler[11]
  PIN prescaler[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END prescaler[12]
  PIN prescaler[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END prescaler[13]
  PIN prescaler[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END prescaler[1]
  PIN prescaler[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END prescaler[2]
  PIN prescaler[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END prescaler[3]
  PIN prescaler[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END prescaler[4]
  PIN prescaler[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END prescaler[5]
  PIN prescaler[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END prescaler[6]
  PIN prescaler[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END prescaler[7]
  PIN prescaler[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END prescaler[8]
  PIN prescaler[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END prescaler[9]
  PIN stop
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 142.660 71.440 146.660 72.040 ;
    END
  END stop
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 140.950 144.350 ;
      LAYER li1 ;
        RECT 5.520 10.795 140.760 144.245 ;
      LAYER met1 ;
        RECT 4.210 10.640 143.910 144.400 ;
      LAYER met2 ;
        RECT 4.230 153.100 57.770 154.090 ;
        RECT 58.610 153.100 60.990 154.090 ;
        RECT 61.830 153.100 64.210 154.090 ;
        RECT 65.050 153.100 67.430 154.090 ;
        RECT 68.270 153.100 70.650 154.090 ;
        RECT 71.490 153.100 73.870 154.090 ;
        RECT 74.710 153.100 77.090 154.090 ;
        RECT 77.930 153.100 80.310 154.090 ;
        RECT 81.150 153.100 83.530 154.090 ;
        RECT 84.370 153.100 86.750 154.090 ;
        RECT 87.590 153.100 89.970 154.090 ;
        RECT 90.810 153.100 93.190 154.090 ;
        RECT 94.030 153.100 96.410 154.090 ;
        RECT 97.250 153.100 99.630 154.090 ;
        RECT 100.470 153.100 102.850 154.090 ;
        RECT 103.690 153.100 106.070 154.090 ;
        RECT 106.910 153.100 109.290 154.090 ;
        RECT 110.130 153.100 112.510 154.090 ;
        RECT 113.350 153.100 115.730 154.090 ;
        RECT 116.570 153.100 118.950 154.090 ;
        RECT 119.790 153.100 122.170 154.090 ;
        RECT 123.010 153.100 125.390 154.090 ;
        RECT 126.230 153.100 128.610 154.090 ;
        RECT 129.450 153.100 131.830 154.090 ;
        RECT 132.670 153.100 135.050 154.090 ;
        RECT 135.890 153.100 138.270 154.090 ;
        RECT 139.110 153.100 141.490 154.090 ;
        RECT 142.330 153.100 144.710 154.090 ;
        RECT 4.230 4.280 144.990 153.100 ;
        RECT 4.230 4.000 28.790 4.280 ;
        RECT 29.630 4.000 44.890 4.280 ;
        RECT 45.730 4.000 144.990 4.280 ;
      LAYER met3 ;
        RECT 3.990 130.240 142.660 144.325 ;
        RECT 3.990 128.840 142.260 130.240 ;
        RECT 3.990 126.840 142.660 128.840 ;
        RECT 3.990 125.440 142.260 126.840 ;
        RECT 3.990 123.440 142.660 125.440 ;
        RECT 3.990 122.040 142.260 123.440 ;
        RECT 3.990 120.040 142.660 122.040 ;
        RECT 4.400 118.640 142.260 120.040 ;
        RECT 3.990 116.640 142.660 118.640 ;
        RECT 4.400 115.240 142.260 116.640 ;
        RECT 3.990 113.240 142.660 115.240 ;
        RECT 4.400 111.840 142.260 113.240 ;
        RECT 3.990 109.840 142.660 111.840 ;
        RECT 4.400 108.440 142.660 109.840 ;
        RECT 3.990 106.440 142.660 108.440 ;
        RECT 4.400 105.040 142.660 106.440 ;
        RECT 3.990 103.040 142.660 105.040 ;
        RECT 4.400 101.640 142.660 103.040 ;
        RECT 3.990 99.640 142.660 101.640 ;
        RECT 4.400 98.240 142.660 99.640 ;
        RECT 3.990 96.240 142.660 98.240 ;
        RECT 4.400 94.840 142.260 96.240 ;
        RECT 3.990 86.040 142.660 94.840 ;
        RECT 4.400 84.640 142.660 86.040 ;
        RECT 3.990 75.840 142.660 84.640 ;
        RECT 4.400 74.440 142.660 75.840 ;
        RECT 3.990 72.440 142.660 74.440 ;
        RECT 3.990 71.040 142.260 72.440 ;
        RECT 3.990 69.040 142.660 71.040 ;
        RECT 4.400 67.640 142.660 69.040 ;
        RECT 3.990 58.840 142.660 67.640 ;
        RECT 4.400 57.440 142.660 58.840 ;
        RECT 3.990 31.640 142.660 57.440 ;
        RECT 3.990 30.240 142.260 31.640 ;
        RECT 3.990 28.240 142.660 30.240 ;
        RECT 3.990 26.840 142.260 28.240 ;
        RECT 3.990 24.840 142.660 26.840 ;
        RECT 3.990 23.440 142.260 24.840 ;
        RECT 3.990 10.715 142.660 23.440 ;
      LAYER met4 ;
        RECT 62.855 23.975 124.825 114.745 ;
  END
END sample_proj
END LIBRARY

