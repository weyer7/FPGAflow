VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fpga
  CLASS BLOCK ;
  FOREIGN fpga ;
  ORIGIN -8.000 -8.000 ;
  SIZE 442.000 BY 436.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 198.070 440.000 198.350 444.000 ;
    END
  END clk
  PIN config_data_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 8.000 225.640 12.000 226.240 ;
    END
  END config_data_in
  PIN config_data_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 235.840 450.000 236.440 ;
    END
  END config_data_out
  PIN config_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.860700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 188.410 440.000 188.690 444.000 ;
    END
  END config_en
  PIN io_east_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 150.840 450.000 151.440 ;
    END
  END io_east_in[0]
  PIN io_east_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 205.240 450.000 205.840 ;
    END
  END io_east_in[10]
  PIN io_east_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 212.040 450.000 212.640 ;
    END
  END io_east_in[11]
  PIN io_east_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 218.840 450.000 219.440 ;
    END
  END io_east_in[12]
  PIN io_east_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 222.240 450.000 222.840 ;
    END
  END io_east_in[13]
  PIN io_east_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.090 8.000 8.370 12.000 ;
    END
  END io_east_in[14]
  PIN io_east_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.310 8.000 11.590 12.000 ;
    END
  END io_east_in[15]
  PIN io_east_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 334.440 450.000 335.040 ;
    END
  END io_east_in[16]
  PIN io_east_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 337.840 450.000 338.440 ;
    END
  END io_east_in[17]
  PIN io_east_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 344.640 450.000 345.240 ;
    END
  END io_east_in[18]
  PIN io_east_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 351.440 450.000 352.040 ;
    END
  END io_east_in[19]
  PIN io_east_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 157.640 450.000 158.240 ;
    END
  END io_east_in[1]
  PIN io_east_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 354.840 450.000 355.440 ;
    END
  END io_east_in[20]
  PIN io_east_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 361.640 450.000 362.240 ;
    END
  END io_east_in[21]
  PIN io_east_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 365.040 450.000 365.640 ;
    END
  END io_east_in[22]
  PIN io_east_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 371.840 450.000 372.440 ;
    END
  END io_east_in[23]
  PIN io_east_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 378.640 450.000 379.240 ;
    END
  END io_east_in[24]
  PIN io_east_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 382.040 450.000 382.640 ;
    END
  END io_east_in[25]
  PIN io_east_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 388.840 450.000 389.440 ;
    END
  END io_east_in[26]
  PIN io_east_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 392.240 450.000 392.840 ;
    END
  END io_east_in[27]
  PIN io_east_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 399.040 450.000 399.640 ;
    END
  END io_east_in[28]
  PIN io_east_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 405.840 450.000 406.440 ;
    END
  END io_east_in[29]
  PIN io_east_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 164.440 450.000 165.040 ;
    END
  END io_east_in[2]
  PIN io_east_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.530 8.000 14.810 12.000 ;
    END
  END io_east_in[30]
  PIN io_east_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.750 8.000 18.030 12.000 ;
    END
  END io_east_in[31]
  PIN io_east_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 167.840 450.000 168.440 ;
    END
  END io_east_in[3]
  PIN io_east_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 174.640 450.000 175.240 ;
    END
  END io_east_in[4]
  PIN io_east_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 178.040 450.000 178.640 ;
    END
  END io_east_in[5]
  PIN io_east_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 184.840 450.000 185.440 ;
    END
  END io_east_in[6]
  PIN io_east_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 191.640 450.000 192.240 ;
    END
  END io_east_in[7]
  PIN io_east_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 195.040 450.000 195.640 ;
    END
  END io_east_in[8]
  PIN io_east_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 201.840 450.000 202.440 ;
    END
  END io_east_in[9]
  PIN io_east_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 76.040 450.000 76.640 ;
    END
  END io_east_out[0]
  PIN io_east_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 130.440 450.000 131.040 ;
    END
  END io_east_out[10]
  PIN io_east_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 137.240 450.000 137.840 ;
    END
  END io_east_out[11]
  PIN io_east_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 140.640 450.000 141.240 ;
    END
  END io_east_out[12]
  PIN io_east_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 147.440 450.000 148.040 ;
    END
  END io_east_out[13]
  PIN io_east_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.810 440.000 253.090 444.000 ;
    END
  END io_east_out[14]
  PIN io_east_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.590 440.000 249.870 444.000 ;
    END
  END io_east_out[15]
  PIN io_east_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 256.240 450.000 256.840 ;
    END
  END io_east_out[16]
  PIN io_east_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 263.040 450.000 263.640 ;
    END
  END io_east_out[17]
  PIN io_east_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 269.840 450.000 270.440 ;
    END
  END io_east_out[18]
  PIN io_east_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 273.240 450.000 273.840 ;
    END
  END io_east_out[19]
  PIN io_east_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 82.840 450.000 83.440 ;
    END
  END io_east_out[1]
  PIN io_east_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 280.040 450.000 280.640 ;
    END
  END io_east_out[20]
  PIN io_east_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 283.440 450.000 284.040 ;
    END
  END io_east_out[21]
  PIN io_east_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 290.240 450.000 290.840 ;
    END
  END io_east_out[22]
  PIN io_east_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 297.040 450.000 297.640 ;
    END
  END io_east_out[23]
  PIN io_east_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 300.440 450.000 301.040 ;
    END
  END io_east_out[24]
  PIN io_east_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 307.240 450.000 307.840 ;
    END
  END io_east_out[25]
  PIN io_east_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 310.640 450.000 311.240 ;
    END
  END io_east_out[26]
  PIN io_east_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 317.440 450.000 318.040 ;
    END
  END io_east_out[27]
  PIN io_east_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 324.240 450.000 324.840 ;
    END
  END io_east_out[28]
  PIN io_east_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 327.640 450.000 328.240 ;
    END
  END io_east_out[29]
  PIN io_east_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 86.240 450.000 86.840 ;
    END
  END io_east_out[2]
  PIN io_east_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.710 440.000 236.990 444.000 ;
    END
  END io_east_out[30]
  PIN io_east_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.170 440.000 214.450 444.000 ;
    END
  END io_east_out[31]
  PIN io_east_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 93.040 450.000 93.640 ;
    END
  END io_east_out[3]
  PIN io_east_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 96.440 450.000 97.040 ;
    END
  END io_east_out[4]
  PIN io_east_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 103.240 450.000 103.840 ;
    END
  END io_east_out[5]
  PIN io_east_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 110.040 450.000 110.640 ;
    END
  END io_east_out[6]
  PIN io_east_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 113.440 450.000 114.040 ;
    END
  END io_east_out[7]
  PIN io_east_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 120.240 450.000 120.840 ;
    END
  END io_east_out[8]
  PIN io_east_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 446.000 123.640 450.000 124.240 ;
    END
  END io_east_out[9]
  PIN io_north_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 75.710 440.000 75.990 444.000 ;
    END
  END io_north_in[0]
  PIN io_north_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 130.450 440.000 130.730 444.000 ;
    END
  END io_north_in[10]
  PIN io_north_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 136.890 440.000 137.170 444.000 ;
    END
  END io_north_in[11]
  PIN io_north_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 140.110 440.000 140.390 444.000 ;
    END
  END io_north_in[12]
  PIN io_north_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 146.550 440.000 146.830 444.000 ;
    END
  END io_north_in[13]
  PIN io_north_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.970 8.000 21.250 12.000 ;
    END
  END io_north_in[14]
  PIN io_north_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.190 8.000 24.470 12.000 ;
    END
  END io_north_in[15]
  PIN io_north_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 262.470 440.000 262.750 444.000 ;
    END
  END io_north_in[16]
  PIN io_north_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 268.910 440.000 269.190 444.000 ;
    END
  END io_north_in[17]
  PIN io_north_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 272.130 440.000 272.410 444.000 ;
    END
  END io_north_in[18]
  PIN io_north_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 278.570 440.000 278.850 444.000 ;
    END
  END io_north_in[19]
  PIN io_north_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 78.930 440.000 79.210 444.000 ;
    END
  END io_north_in[1]
  PIN io_north_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 285.010 440.000 285.290 444.000 ;
    END
  END io_north_in[20]
  PIN io_north_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 288.230 440.000 288.510 444.000 ;
    END
  END io_north_in[21]
  PIN io_north_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 294.670 440.000 294.950 444.000 ;
    END
  END io_north_in[22]
  PIN io_north_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 301.110 440.000 301.390 444.000 ;
    END
  END io_north_in[23]
  PIN io_north_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 307.550 440.000 307.830 444.000 ;
    END
  END io_north_in[24]
  PIN io_north_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 310.770 440.000 311.050 444.000 ;
    END
  END io_north_in[25]
  PIN io_north_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 317.210 440.000 317.490 444.000 ;
    END
  END io_north_in[26]
  PIN io_north_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 323.650 440.000 323.930 444.000 ;
    END
  END io_north_in[27]
  PIN io_north_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 326.870 440.000 327.150 444.000 ;
    END
  END io_north_in[28]
  PIN io_north_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 333.310 440.000 333.590 444.000 ;
    END
  END io_north_in[29]
  PIN io_north_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 85.370 440.000 85.650 444.000 ;
    END
  END io_north_in[2]
  PIN io_north_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.410 8.000 27.690 12.000 ;
    END
  END io_north_in[30]
  PIN io_north_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.630 8.000 30.910 12.000 ;
    END
  END io_north_in[31]
  PIN io_north_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 91.810 440.000 92.090 444.000 ;
    END
  END io_north_in[3]
  PIN io_north_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 98.250 440.000 98.530 444.000 ;
    END
  END io_north_in[4]
  PIN io_north_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 101.470 440.000 101.750 444.000 ;
    END
  END io_north_in[5]
  PIN io_north_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 107.910 440.000 108.190 444.000 ;
    END
  END io_north_in[6]
  PIN io_north_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 114.350 440.000 114.630 444.000 ;
    END
  END io_north_in[7]
  PIN io_north_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 117.570 440.000 117.850 444.000 ;
    END
  END io_north_in[8]
  PIN io_north_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 124.010 440.000 124.290 444.000 ;
    END
  END io_north_in[9]
  PIN io_north_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 152.990 440.000 153.270 444.000 ;
    END
  END io_north_out[0]
  PIN io_north_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 207.730 440.000 208.010 444.000 ;
    END
  END io_north_out[10]
  PIN io_north_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 210.950 440.000 211.230 444.000 ;
    END
  END io_north_out[11]
  PIN io_north_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 217.390 440.000 217.670 444.000 ;
    END
  END io_north_out[12]
  PIN io_north_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 220.610 440.000 220.890 444.000 ;
    END
  END io_north_out[13]
  PIN io_north_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.150 440.000 243.430 444.000 ;
    END
  END io_north_out[14]
  PIN io_north_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 239.240 450.000 239.840 ;
    END
  END io_north_out[15]
  PIN io_north_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 339.750 440.000 340.030 444.000 ;
    END
  END io_north_out[16]
  PIN io_north_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 346.190 440.000 346.470 444.000 ;
    END
  END io_north_out[17]
  PIN io_north_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 349.410 440.000 349.690 444.000 ;
    END
  END io_north_out[18]
  PIN io_north_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 355.850 440.000 356.130 444.000 ;
    END
  END io_north_out[19]
  PIN io_north_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 156.210 440.000 156.490 444.000 ;
    END
  END io_north_out[1]
  PIN io_north_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 362.290 440.000 362.570 444.000 ;
    END
  END io_north_out[20]
  PIN io_north_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 365.510 440.000 365.790 444.000 ;
    END
  END io_north_out[21]
  PIN io_north_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 371.950 440.000 372.230 444.000 ;
    END
  END io_north_out[22]
  PIN io_north_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 378.390 440.000 378.670 444.000 ;
    END
  END io_north_out[23]
  PIN io_north_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 384.830 440.000 385.110 444.000 ;
    END
  END io_north_out[24]
  PIN io_north_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 388.050 440.000 388.330 444.000 ;
    END
  END io_north_out[25]
  PIN io_north_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 394.490 440.000 394.770 444.000 ;
    END
  END io_north_out[26]
  PIN io_north_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 400.930 440.000 401.210 444.000 ;
    END
  END io_north_out[27]
  PIN io_north_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 404.150 440.000 404.430 444.000 ;
    END
  END io_north_out[28]
  PIN io_north_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 410.590 440.000 410.870 444.000 ;
    END
  END io_north_out[29]
  PIN io_north_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 162.650 440.000 162.930 444.000 ;
    END
  END io_north_out[2]
  PIN io_north_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 229.040 450.000 229.640 ;
    END
  END io_north_out[30]
  PIN io_north_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.830 440.000 224.110 444.000 ;
    END
  END io_north_out[31]
  PIN io_north_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 169.090 440.000 169.370 444.000 ;
    END
  END io_north_out[3]
  PIN io_north_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 175.530 440.000 175.810 444.000 ;
    END
  END io_north_out[4]
  PIN io_north_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 178.750 440.000 179.030 444.000 ;
    END
  END io_north_out[5]
  PIN io_north_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 185.190 440.000 185.470 444.000 ;
    END
  END io_north_out[6]
  PIN io_north_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 191.630 440.000 191.910 444.000 ;
    END
  END io_north_out[7]
  PIN io_north_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 194.850 440.000 195.130 444.000 ;
    END
  END io_north_out[8]
  PIN io_north_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 201.290 440.000 201.570 444.000 ;
    END
  END io_north_out[9]
  PIN io_south_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 152.990 8.000 153.270 12.000 ;
    END
  END io_south_in[0]
  PIN io_south_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 207.730 8.000 208.010 12.000 ;
    END
  END io_south_in[10]
  PIN io_south_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 214.170 8.000 214.450 12.000 ;
    END
  END io_south_in[11]
  PIN io_south_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 217.390 8.000 217.670 12.000 ;
    END
  END io_south_in[12]
  PIN io_south_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 223.830 8.000 224.110 12.000 ;
    END
  END io_south_in[13]
  PIN io_south_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.850 8.000 34.130 12.000 ;
    END
  END io_south_in[14]
  PIN io_south_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.070 8.000 37.350 12.000 ;
    END
  END io_south_in[15]
  PIN io_south_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 339.750 8.000 340.030 12.000 ;
    END
  END io_south_in[16]
  PIN io_south_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 346.190 8.000 346.470 12.000 ;
    END
  END io_south_in[17]
  PIN io_south_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 349.410 8.000 349.690 12.000 ;
    END
  END io_south_in[18]
  PIN io_south_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 355.850 8.000 356.130 12.000 ;
    END
  END io_south_in[19]
  PIN io_south_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 156.210 8.000 156.490 12.000 ;
    END
  END io_south_in[1]
  PIN io_south_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 362.290 8.000 362.570 12.000 ;
    END
  END io_south_in[20]
  PIN io_south_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 365.510 8.000 365.790 12.000 ;
    END
  END io_south_in[21]
  PIN io_south_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 371.950 8.000 372.230 12.000 ;
    END
  END io_south_in[22]
  PIN io_south_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 378.390 8.000 378.670 12.000 ;
    END
  END io_south_in[23]
  PIN io_south_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 384.830 8.000 385.110 12.000 ;
    END
  END io_south_in[24]
  PIN io_south_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 388.050 8.000 388.330 12.000 ;
    END
  END io_south_in[25]
  PIN io_south_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 394.490 8.000 394.770 12.000 ;
    END
  END io_south_in[26]
  PIN io_south_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 400.930 8.000 401.210 12.000 ;
    END
  END io_south_in[27]
  PIN io_south_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 48.840 450.000 49.440 ;
    END
  END io_south_in[28]
  PIN io_south_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 52.240 450.000 52.840 ;
    END
  END io_south_in[29]
  PIN io_south_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 162.650 8.000 162.930 12.000 ;
    END
  END io_south_in[2]
  PIN io_south_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.290 8.000 40.570 12.000 ;
    END
  END io_south_in[30]
  PIN io_south_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.510 8.000 43.790 12.000 ;
    END
  END io_south_in[31]
  PIN io_south_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 169.090 8.000 169.370 12.000 ;
    END
  END io_south_in[3]
  PIN io_south_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 175.530 8.000 175.810 12.000 ;
    END
  END io_south_in[4]
  PIN io_south_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 178.750 8.000 179.030 12.000 ;
    END
  END io_south_in[5]
  PIN io_south_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 185.190 8.000 185.470 12.000 ;
    END
  END io_south_in[6]
  PIN io_south_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 191.630 8.000 191.910 12.000 ;
    END
  END io_south_in[7]
  PIN io_south_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 194.850 8.000 195.130 12.000 ;
    END
  END io_south_in[8]
  PIN io_south_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 201.290 8.000 201.570 12.000 ;
    END
  END io_south_in[9]
  PIN io_south_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 75.710 8.000 75.990 12.000 ;
    END
  END io_south_out[0]
  PIN io_south_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 130.450 8.000 130.730 12.000 ;
    END
  END io_south_out[10]
  PIN io_south_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 136.890 8.000 137.170 12.000 ;
    END
  END io_south_out[11]
  PIN io_south_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 140.110 8.000 140.390 12.000 ;
    END
  END io_south_out[12]
  PIN io_south_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 146.550 8.000 146.830 12.000 ;
    END
  END io_south_out[13]
  PIN io_south_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.050 440.000 227.330 444.000 ;
    END
  END io_south_out[14]
  PIN io_south_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.490 440.000 233.770 444.000 ;
    END
  END io_south_out[15]
  PIN io_south_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 262.470 8.000 262.750 12.000 ;
    END
  END io_south_out[16]
  PIN io_south_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 268.910 8.000 269.190 12.000 ;
    END
  END io_south_out[17]
  PIN io_south_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 272.130 8.000 272.410 12.000 ;
    END
  END io_south_out[18]
  PIN io_south_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 278.570 8.000 278.850 12.000 ;
    END
  END io_south_out[19]
  PIN io_south_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 78.930 8.000 79.210 12.000 ;
    END
  END io_south_out[1]
  PIN io_south_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 285.010 8.000 285.290 12.000 ;
    END
  END io_south_out[20]
  PIN io_south_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 288.230 8.000 288.510 12.000 ;
    END
  END io_south_out[21]
  PIN io_south_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 294.670 8.000 294.950 12.000 ;
    END
  END io_south_out[22]
  PIN io_south_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 301.110 8.000 301.390 12.000 ;
    END
  END io_south_out[23]
  PIN io_south_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 307.550 8.000 307.830 12.000 ;
    END
  END io_south_out[24]
  PIN io_south_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 310.770 8.000 311.050 12.000 ;
    END
  END io_south_out[25]
  PIN io_south_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 317.210 8.000 317.490 12.000 ;
    END
  END io_south_out[26]
  PIN io_south_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 323.650 8.000 323.930 12.000 ;
    END
  END io_south_out[27]
  PIN io_south_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 326.870 8.000 327.150 12.000 ;
    END
  END io_south_out[28]
  PIN io_south_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 333.310 8.000 333.590 12.000 ;
    END
  END io_south_out[29]
  PIN io_south_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 85.370 8.000 85.650 12.000 ;
    END
  END io_south_out[2]
  PIN io_south_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 225.640 450.000 226.240 ;
    END
  END io_south_out[30]
  PIN io_south_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 232.440 450.000 233.040 ;
    END
  END io_south_out[31]
  PIN io_south_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 91.810 8.000 92.090 12.000 ;
    END
  END io_south_out[3]
  PIN io_south_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 98.250 8.000 98.530 12.000 ;
    END
  END io_south_out[4]
  PIN io_south_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 101.470 8.000 101.750 12.000 ;
    END
  END io_south_out[5]
  PIN io_south_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 107.910 8.000 108.190 12.000 ;
    END
  END io_south_out[6]
  PIN io_south_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 114.350 8.000 114.630 12.000 ;
    END
  END io_south_out[7]
  PIN io_south_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 117.570 8.000 117.850 12.000 ;
    END
  END io_south_out[8]
  PIN io_south_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 124.010 8.000 124.290 12.000 ;
    END
  END io_south_out[9]
  PIN io_west_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 8.000 76.040 12.000 76.640 ;
    END
  END io_west_in[0]
  PIN io_west_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 8.000 130.440 12.000 131.040 ;
    END
  END io_west_in[10]
  PIN io_west_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 8.000 137.240 12.000 137.840 ;
    END
  END io_west_in[11]
  PIN io_west_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 8.000 140.640 12.000 141.240 ;
    END
  END io_west_in[12]
  PIN io_west_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 8.000 147.440 12.000 148.040 ;
    END
  END io_west_in[13]
  PIN io_west_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.730 8.000 47.010 12.000 ;
    END
  END io_west_in[14]
  PIN io_west_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.950 8.000 50.230 12.000 ;
    END
  END io_west_in[15]
  PIN io_west_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 8.000 256.240 12.000 256.840 ;
    END
  END io_west_in[16]
  PIN io_west_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 8.000 263.040 12.000 263.640 ;
    END
  END io_west_in[17]
  PIN io_west_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 8.000 269.840 12.000 270.440 ;
    END
  END io_west_in[18]
  PIN io_west_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 8.000 273.240 12.000 273.840 ;
    END
  END io_west_in[19]
  PIN io_west_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 8.000 82.840 12.000 83.440 ;
    END
  END io_west_in[1]
  PIN io_west_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 8.000 280.040 12.000 280.640 ;
    END
  END io_west_in[20]
  PIN io_west_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 8.000 283.440 12.000 284.040 ;
    END
  END io_west_in[21]
  PIN io_west_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 8.000 290.240 12.000 290.840 ;
    END
  END io_west_in[22]
  PIN io_west_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 8.000 297.040 12.000 297.640 ;
    END
  END io_west_in[23]
  PIN io_west_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 8.000 300.440 12.000 301.040 ;
    END
  END io_west_in[24]
  PIN io_west_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 8.000 307.240 12.000 307.840 ;
    END
  END io_west_in[25]
  PIN io_west_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 8.000 310.640 12.000 311.240 ;
    END
  END io_west_in[26]
  PIN io_west_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 8.000 317.440 12.000 318.040 ;
    END
  END io_west_in[27]
  PIN io_west_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 8.000 324.240 12.000 324.840 ;
    END
  END io_west_in[28]
  PIN io_west_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 8.000 327.640 12.000 328.240 ;
    END
  END io_west_in[29]
  PIN io_west_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 8.000 86.240 12.000 86.840 ;
    END
  END io_west_in[2]
  PIN io_west_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.170 8.000 53.450 12.000 ;
    END
  END io_west_in[30]
  PIN io_west_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.390 8.000 56.670 12.000 ;
    END
  END io_west_in[31]
  PIN io_west_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 8.000 93.040 12.000 93.640 ;
    END
  END io_west_in[3]
  PIN io_west_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 8.000 96.440 12.000 97.040 ;
    END
  END io_west_in[4]
  PIN io_west_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 8.000 103.240 12.000 103.840 ;
    END
  END io_west_in[5]
  PIN io_west_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 8.000 110.040 12.000 110.640 ;
    END
  END io_west_in[6]
  PIN io_west_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 8.000 113.440 12.000 114.040 ;
    END
  END io_west_in[7]
  PIN io_west_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 8.000 120.240 12.000 120.840 ;
    END
  END io_west_in[8]
  PIN io_west_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 8.000 123.640 12.000 124.240 ;
    END
  END io_west_in[9]
  PIN io_west_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 150.840 12.000 151.440 ;
    END
  END io_west_out[0]
  PIN io_west_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 205.240 12.000 205.840 ;
    END
  END io_west_out[10]
  PIN io_west_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 212.040 12.000 212.640 ;
    END
  END io_west_out[11]
  PIN io_west_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 218.840 12.000 219.440 ;
    END
  END io_west_out[12]
  PIN io_west_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 222.240 12.000 222.840 ;
    END
  END io_west_out[13]
  PIN io_west_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.270 440.000 230.550 444.000 ;
    END
  END io_west_out[14]
  PIN io_west_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 446.000 242.640 450.000 243.240 ;
    END
  END io_west_out[15]
  PIN io_west_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 334.440 12.000 335.040 ;
    END
  END io_west_out[16]
  PIN io_west_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 337.840 12.000 338.440 ;
    END
  END io_west_out[17]
  PIN io_west_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 344.640 12.000 345.240 ;
    END
  END io_west_out[18]
  PIN io_west_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 351.440 12.000 352.040 ;
    END
  END io_west_out[19]
  PIN io_west_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 157.640 12.000 158.240 ;
    END
  END io_west_out[1]
  PIN io_west_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 354.840 12.000 355.440 ;
    END
  END io_west_out[20]
  PIN io_west_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 361.640 12.000 362.240 ;
    END
  END io_west_out[21]
  PIN io_west_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 365.040 12.000 365.640 ;
    END
  END io_west_out[22]
  PIN io_west_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 371.840 12.000 372.440 ;
    END
  END io_west_out[23]
  PIN io_west_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 378.640 12.000 379.240 ;
    END
  END io_west_out[24]
  PIN io_west_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 382.040 12.000 382.640 ;
    END
  END io_west_out[25]
  PIN io_west_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 388.840 12.000 389.440 ;
    END
  END io_west_out[26]
  PIN io_west_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 392.240 12.000 392.840 ;
    END
  END io_west_out[27]
  PIN io_west_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 399.040 12.000 399.640 ;
    END
  END io_west_out[28]
  PIN io_west_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 53.170 440.000 53.450 444.000 ;
    END
  END io_west_out[29]
  PIN io_west_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 164.440 12.000 165.040 ;
    END
  END io_west_out[2]
  PIN io_west_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.370 440.000 246.650 444.000 ;
    END
  END io_west_out[30]
  PIN io_west_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.930 440.000 240.210 444.000 ;
    END
  END io_west_out[31]
  PIN io_west_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 167.840 12.000 168.440 ;
    END
  END io_west_out[3]
  PIN io_west_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 174.640 12.000 175.240 ;
    END
  END io_west_out[4]
  PIN io_west_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 178.040 12.000 178.640 ;
    END
  END io_west_out[5]
  PIN io_west_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 184.840 12.000 185.440 ;
    END
  END io_west_out[6]
  PIN io_west_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 191.640 12.000 192.240 ;
    END
  END io_west_out[7]
  PIN io_west_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 195.040 12.000 195.640 ;
    END
  END io_west_out[8]
  PIN io_west_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 8.000 201.840 12.000 202.440 ;
    END
  END io_west_out[9]
  PIN le_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 62.440 450.000 63.040 ;
    END
  END le_clk
  PIN le_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 65.840 450.000 66.440 ;
    END
  END le_en
  PIN le_nrst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 446.000 72.640 450.000 73.240 ;
    END
  END le_nrst
  PIN nrst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.860700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 204.510 440.000 204.790 444.000 ;
    END
  END nrst
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 16.780 16.880 18.380 445.520 ;
    END
    PORT
      LAYER met5 ;
        RECT 16.780 16.880 450.580 18.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 16.780 443.920 450.580 445.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 448.980 16.880 450.580 445.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 88.580 13.580 90.180 50.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 88.580 405.145 90.180 448.820 ;
    END
    PORT
      LAYER met4 ;
        RECT 180.580 13.580 182.180 50.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 180.580 405.145 182.180 448.820 ;
    END
    PORT
      LAYER met4 ;
        RECT 272.580 13.580 274.180 50.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 272.580 405.145 274.180 448.820 ;
    END
    PORT
      LAYER met4 ;
        RECT 364.580 13.580 366.180 50.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 364.580 405.145 366.180 448.820 ;
    END
    PORT
      LAYER met5 ;
        RECT 13.480 88.680 453.880 90.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 13.480 180.680 453.880 182.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 13.480 272.680 453.880 274.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 13.480 364.680 453.880 366.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 29.740 35.120 31.340 424.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 432.700 35.120 434.300 424.560 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 13.480 13.580 15.080 448.820 ;
    END
    PORT
      LAYER met5 ;
        RECT 13.480 13.580 453.880 15.180 ;
    END
    PORT
      LAYER met5 ;
        RECT 13.480 447.220 453.880 448.820 ;
    END
    PORT
      LAYER met4 ;
        RECT 452.280 13.580 453.880 448.820 ;
    END
    PORT
      LAYER met4 ;
        RECT 91.880 13.580 93.480 50.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 91.880 405.145 93.480 448.820 ;
    END
    PORT
      LAYER met4 ;
        RECT 183.880 13.580 185.480 50.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 183.880 405.145 185.480 448.820 ;
    END
    PORT
      LAYER met4 ;
        RECT 275.880 13.580 277.480 50.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 275.880 405.145 277.480 448.820 ;
    END
    PORT
      LAYER met4 ;
        RECT 367.880 13.580 369.480 50.935 ;
    END
    PORT
      LAYER met4 ;
        RECT 367.880 405.145 369.480 448.820 ;
    END
    PORT
      LAYER met5 ;
        RECT 13.480 91.980 453.880 93.580 ;
    END
    PORT
      LAYER met5 ;
        RECT 13.480 183.980 453.880 185.580 ;
    END
    PORT
      LAYER met5 ;
        RECT 13.480 275.980 453.880 277.580 ;
    END
    PORT
      LAYER met5 ;
        RECT 13.480 367.980 453.880 369.580 ;
    END
    PORT
      LAYER met4 ;
        RECT 33.420 35.120 35.020 424.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 436.380 35.120 437.980 424.560 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 24.190 24.395 443.170 438.005 ;
      LAYER li1 ;
        RECT 24.380 24.395 442.980 438.005 ;
      LAYER met1 ;
        RECT 13.590 24.240 444.930 438.160 ;
      LAYER met2 ;
        RECT 13.610 439.720 52.890 440.000 ;
        RECT 53.730 439.720 75.430 440.000 ;
        RECT 76.270 439.720 78.650 440.000 ;
        RECT 79.490 439.720 85.090 440.000 ;
        RECT 85.930 439.720 91.530 440.000 ;
        RECT 92.370 439.720 97.970 440.000 ;
        RECT 98.810 439.720 101.190 440.000 ;
        RECT 102.030 439.720 107.630 440.000 ;
        RECT 108.470 439.720 114.070 440.000 ;
        RECT 114.910 439.720 117.290 440.000 ;
        RECT 118.130 439.720 123.730 440.000 ;
        RECT 124.570 439.720 130.170 440.000 ;
        RECT 131.010 439.720 136.610 440.000 ;
        RECT 137.450 439.720 139.830 440.000 ;
        RECT 140.670 439.720 146.270 440.000 ;
        RECT 147.110 439.720 152.710 440.000 ;
        RECT 153.550 439.720 155.930 440.000 ;
        RECT 156.770 439.720 162.370 440.000 ;
        RECT 163.210 439.720 168.810 440.000 ;
        RECT 169.650 439.720 175.250 440.000 ;
        RECT 176.090 439.720 178.470 440.000 ;
        RECT 179.310 439.720 184.910 440.000 ;
        RECT 185.750 439.720 188.130 440.000 ;
        RECT 188.970 439.720 191.350 440.000 ;
        RECT 192.190 439.720 194.570 440.000 ;
        RECT 195.410 439.720 197.790 440.000 ;
        RECT 198.630 439.720 201.010 440.000 ;
        RECT 201.850 439.720 204.230 440.000 ;
        RECT 205.070 439.720 207.450 440.000 ;
        RECT 208.290 439.720 210.670 440.000 ;
        RECT 211.510 439.720 213.890 440.000 ;
        RECT 214.730 439.720 217.110 440.000 ;
        RECT 217.950 439.720 220.330 440.000 ;
        RECT 221.170 439.720 223.550 440.000 ;
        RECT 224.390 439.720 226.770 440.000 ;
        RECT 227.610 439.720 229.990 440.000 ;
        RECT 230.830 439.720 233.210 440.000 ;
        RECT 234.050 439.720 236.430 440.000 ;
        RECT 237.270 439.720 239.650 440.000 ;
        RECT 240.490 439.720 242.870 440.000 ;
        RECT 243.710 439.720 246.090 440.000 ;
        RECT 246.930 439.720 249.310 440.000 ;
        RECT 250.150 439.720 252.530 440.000 ;
        RECT 253.370 439.720 262.190 440.000 ;
        RECT 263.030 439.720 268.630 440.000 ;
        RECT 269.470 439.720 271.850 440.000 ;
        RECT 272.690 439.720 278.290 440.000 ;
        RECT 279.130 439.720 284.730 440.000 ;
        RECT 285.570 439.720 287.950 440.000 ;
        RECT 288.790 439.720 294.390 440.000 ;
        RECT 295.230 439.720 300.830 440.000 ;
        RECT 301.670 439.720 307.270 440.000 ;
        RECT 308.110 439.720 310.490 440.000 ;
        RECT 311.330 439.720 316.930 440.000 ;
        RECT 317.770 439.720 323.370 440.000 ;
        RECT 324.210 439.720 326.590 440.000 ;
        RECT 327.430 439.720 333.030 440.000 ;
        RECT 333.870 439.720 339.470 440.000 ;
        RECT 340.310 439.720 345.910 440.000 ;
        RECT 346.750 439.720 349.130 440.000 ;
        RECT 349.970 439.720 355.570 440.000 ;
        RECT 356.410 439.720 362.010 440.000 ;
        RECT 362.850 439.720 365.230 440.000 ;
        RECT 366.070 439.720 371.670 440.000 ;
        RECT 372.510 439.720 378.110 440.000 ;
        RECT 378.950 439.720 384.550 440.000 ;
        RECT 385.390 439.720 387.770 440.000 ;
        RECT 388.610 439.720 394.210 440.000 ;
        RECT 395.050 439.720 400.650 440.000 ;
        RECT 401.490 439.720 403.870 440.000 ;
        RECT 404.710 439.720 410.310 440.000 ;
        RECT 411.150 439.720 444.910 440.000 ;
        RECT 13.610 12.280 444.910 439.720 ;
        RECT 13.610 12.000 14.250 12.280 ;
        RECT 15.090 12.000 17.470 12.280 ;
        RECT 18.310 12.000 20.690 12.280 ;
        RECT 21.530 12.000 23.910 12.280 ;
        RECT 24.750 12.000 27.130 12.280 ;
        RECT 27.970 12.000 30.350 12.280 ;
        RECT 31.190 12.000 33.570 12.280 ;
        RECT 34.410 12.000 36.790 12.280 ;
        RECT 37.630 12.000 40.010 12.280 ;
        RECT 40.850 12.000 43.230 12.280 ;
        RECT 44.070 12.000 46.450 12.280 ;
        RECT 47.290 12.000 49.670 12.280 ;
        RECT 50.510 12.000 52.890 12.280 ;
        RECT 53.730 12.000 56.110 12.280 ;
        RECT 56.950 12.000 75.430 12.280 ;
        RECT 76.270 12.000 78.650 12.280 ;
        RECT 79.490 12.000 85.090 12.280 ;
        RECT 85.930 12.000 91.530 12.280 ;
        RECT 92.370 12.000 97.970 12.280 ;
        RECT 98.810 12.000 101.190 12.280 ;
        RECT 102.030 12.000 107.630 12.280 ;
        RECT 108.470 12.000 114.070 12.280 ;
        RECT 114.910 12.000 117.290 12.280 ;
        RECT 118.130 12.000 123.730 12.280 ;
        RECT 124.570 12.000 130.170 12.280 ;
        RECT 131.010 12.000 136.610 12.280 ;
        RECT 137.450 12.000 139.830 12.280 ;
        RECT 140.670 12.000 146.270 12.280 ;
        RECT 147.110 12.000 152.710 12.280 ;
        RECT 153.550 12.000 155.930 12.280 ;
        RECT 156.770 12.000 162.370 12.280 ;
        RECT 163.210 12.000 168.810 12.280 ;
        RECT 169.650 12.000 175.250 12.280 ;
        RECT 176.090 12.000 178.470 12.280 ;
        RECT 179.310 12.000 184.910 12.280 ;
        RECT 185.750 12.000 191.350 12.280 ;
        RECT 192.190 12.000 194.570 12.280 ;
        RECT 195.410 12.000 201.010 12.280 ;
        RECT 201.850 12.000 207.450 12.280 ;
        RECT 208.290 12.000 213.890 12.280 ;
        RECT 214.730 12.000 217.110 12.280 ;
        RECT 217.950 12.000 223.550 12.280 ;
        RECT 224.390 12.000 262.190 12.280 ;
        RECT 263.030 12.000 268.630 12.280 ;
        RECT 269.470 12.000 271.850 12.280 ;
        RECT 272.690 12.000 278.290 12.280 ;
        RECT 279.130 12.000 284.730 12.280 ;
        RECT 285.570 12.000 287.950 12.280 ;
        RECT 288.790 12.000 294.390 12.280 ;
        RECT 295.230 12.000 300.830 12.280 ;
        RECT 301.670 12.000 307.270 12.280 ;
        RECT 308.110 12.000 310.490 12.280 ;
        RECT 311.330 12.000 316.930 12.280 ;
        RECT 317.770 12.000 323.370 12.280 ;
        RECT 324.210 12.000 326.590 12.280 ;
        RECT 327.430 12.000 333.030 12.280 ;
        RECT 333.870 12.000 339.470 12.280 ;
        RECT 340.310 12.000 345.910 12.280 ;
        RECT 346.750 12.000 349.130 12.280 ;
        RECT 349.970 12.000 355.570 12.280 ;
        RECT 356.410 12.000 362.010 12.280 ;
        RECT 362.850 12.000 365.230 12.280 ;
        RECT 366.070 12.000 371.670 12.280 ;
        RECT 372.510 12.000 378.110 12.280 ;
        RECT 378.950 12.000 384.550 12.280 ;
        RECT 385.390 12.000 387.770 12.280 ;
        RECT 388.610 12.000 394.210 12.280 ;
        RECT 395.050 12.000 400.650 12.280 ;
        RECT 401.490 12.000 444.910 12.280 ;
      LAYER met3 ;
        RECT 12.000 406.840 446.000 438.085 ;
        RECT 12.000 405.440 445.600 406.840 ;
        RECT 12.000 400.040 446.000 405.440 ;
        RECT 12.400 398.640 445.600 400.040 ;
        RECT 12.000 393.240 446.000 398.640 ;
        RECT 12.400 391.840 445.600 393.240 ;
        RECT 12.000 389.840 446.000 391.840 ;
        RECT 12.400 388.440 445.600 389.840 ;
        RECT 12.000 383.040 446.000 388.440 ;
        RECT 12.400 381.640 445.600 383.040 ;
        RECT 12.000 379.640 446.000 381.640 ;
        RECT 12.400 378.240 445.600 379.640 ;
        RECT 12.000 372.840 446.000 378.240 ;
        RECT 12.400 371.440 445.600 372.840 ;
        RECT 12.000 366.040 446.000 371.440 ;
        RECT 12.400 364.640 445.600 366.040 ;
        RECT 12.000 362.640 446.000 364.640 ;
        RECT 12.400 361.240 445.600 362.640 ;
        RECT 12.000 355.840 446.000 361.240 ;
        RECT 12.400 354.440 445.600 355.840 ;
        RECT 12.000 352.440 446.000 354.440 ;
        RECT 12.400 351.040 445.600 352.440 ;
        RECT 12.000 345.640 446.000 351.040 ;
        RECT 12.400 344.240 445.600 345.640 ;
        RECT 12.000 338.840 446.000 344.240 ;
        RECT 12.400 337.440 445.600 338.840 ;
        RECT 12.000 335.440 446.000 337.440 ;
        RECT 12.400 334.040 445.600 335.440 ;
        RECT 12.000 328.640 446.000 334.040 ;
        RECT 12.400 327.240 445.600 328.640 ;
        RECT 12.000 325.240 446.000 327.240 ;
        RECT 12.400 323.840 445.600 325.240 ;
        RECT 12.000 318.440 446.000 323.840 ;
        RECT 12.400 317.040 445.600 318.440 ;
        RECT 12.000 311.640 446.000 317.040 ;
        RECT 12.400 310.240 445.600 311.640 ;
        RECT 12.000 308.240 446.000 310.240 ;
        RECT 12.400 306.840 445.600 308.240 ;
        RECT 12.000 301.440 446.000 306.840 ;
        RECT 12.400 300.040 445.600 301.440 ;
        RECT 12.000 298.040 446.000 300.040 ;
        RECT 12.400 296.640 445.600 298.040 ;
        RECT 12.000 291.240 446.000 296.640 ;
        RECT 12.400 289.840 445.600 291.240 ;
        RECT 12.000 284.440 446.000 289.840 ;
        RECT 12.400 283.040 445.600 284.440 ;
        RECT 12.000 281.040 446.000 283.040 ;
        RECT 12.400 279.640 445.600 281.040 ;
        RECT 12.000 274.240 446.000 279.640 ;
        RECT 12.400 272.840 445.600 274.240 ;
        RECT 12.000 270.840 446.000 272.840 ;
        RECT 12.400 269.440 445.600 270.840 ;
        RECT 12.000 264.040 446.000 269.440 ;
        RECT 12.400 262.640 445.600 264.040 ;
        RECT 12.000 257.240 446.000 262.640 ;
        RECT 12.400 255.840 445.600 257.240 ;
        RECT 12.000 243.640 446.000 255.840 ;
        RECT 12.000 242.240 445.600 243.640 ;
        RECT 12.000 240.240 446.000 242.240 ;
        RECT 12.000 238.840 445.600 240.240 ;
        RECT 12.000 236.840 446.000 238.840 ;
        RECT 12.000 235.440 445.600 236.840 ;
        RECT 12.000 233.440 446.000 235.440 ;
        RECT 12.000 232.040 445.600 233.440 ;
        RECT 12.000 230.040 446.000 232.040 ;
        RECT 12.000 228.640 445.600 230.040 ;
        RECT 12.000 226.640 446.000 228.640 ;
        RECT 12.400 225.240 445.600 226.640 ;
        RECT 12.000 223.240 446.000 225.240 ;
        RECT 12.400 221.840 445.600 223.240 ;
        RECT 12.000 219.840 446.000 221.840 ;
        RECT 12.400 218.440 445.600 219.840 ;
        RECT 12.000 213.040 446.000 218.440 ;
        RECT 12.400 211.640 445.600 213.040 ;
        RECT 12.000 206.240 446.000 211.640 ;
        RECT 12.400 204.840 445.600 206.240 ;
        RECT 12.000 202.840 446.000 204.840 ;
        RECT 12.400 201.440 445.600 202.840 ;
        RECT 12.000 196.040 446.000 201.440 ;
        RECT 12.400 194.640 445.600 196.040 ;
        RECT 12.000 192.640 446.000 194.640 ;
        RECT 12.400 191.240 445.600 192.640 ;
        RECT 12.000 185.840 446.000 191.240 ;
        RECT 12.400 184.440 445.600 185.840 ;
        RECT 12.000 179.040 446.000 184.440 ;
        RECT 12.400 177.640 445.600 179.040 ;
        RECT 12.000 175.640 446.000 177.640 ;
        RECT 12.400 174.240 445.600 175.640 ;
        RECT 12.000 168.840 446.000 174.240 ;
        RECT 12.400 167.440 445.600 168.840 ;
        RECT 12.000 165.440 446.000 167.440 ;
        RECT 12.400 164.040 445.600 165.440 ;
        RECT 12.000 158.640 446.000 164.040 ;
        RECT 12.400 157.240 445.600 158.640 ;
        RECT 12.000 151.840 446.000 157.240 ;
        RECT 12.400 150.440 445.600 151.840 ;
        RECT 12.000 148.440 446.000 150.440 ;
        RECT 12.400 147.040 445.600 148.440 ;
        RECT 12.000 141.640 446.000 147.040 ;
        RECT 12.400 140.240 445.600 141.640 ;
        RECT 12.000 138.240 446.000 140.240 ;
        RECT 12.400 136.840 445.600 138.240 ;
        RECT 12.000 131.440 446.000 136.840 ;
        RECT 12.400 130.040 445.600 131.440 ;
        RECT 12.000 124.640 446.000 130.040 ;
        RECT 12.400 123.240 445.600 124.640 ;
        RECT 12.000 121.240 446.000 123.240 ;
        RECT 12.400 119.840 445.600 121.240 ;
        RECT 12.000 114.440 446.000 119.840 ;
        RECT 12.400 113.040 445.600 114.440 ;
        RECT 12.000 111.040 446.000 113.040 ;
        RECT 12.400 109.640 445.600 111.040 ;
        RECT 12.000 104.240 446.000 109.640 ;
        RECT 12.400 102.840 445.600 104.240 ;
        RECT 12.000 97.440 446.000 102.840 ;
        RECT 12.400 96.040 445.600 97.440 ;
        RECT 12.000 94.040 446.000 96.040 ;
        RECT 12.400 92.640 445.600 94.040 ;
        RECT 12.000 87.240 446.000 92.640 ;
        RECT 12.400 85.840 445.600 87.240 ;
        RECT 12.000 83.840 446.000 85.840 ;
        RECT 12.400 82.440 445.600 83.840 ;
        RECT 12.000 77.040 446.000 82.440 ;
        RECT 12.400 75.640 445.600 77.040 ;
        RECT 12.000 73.640 446.000 75.640 ;
        RECT 12.000 72.240 445.600 73.640 ;
        RECT 12.000 66.840 446.000 72.240 ;
        RECT 12.000 65.440 445.600 66.840 ;
        RECT 12.000 63.440 446.000 65.440 ;
        RECT 12.000 62.040 445.600 63.440 ;
        RECT 12.000 53.240 446.000 62.040 ;
        RECT 12.000 51.840 445.600 53.240 ;
        RECT 12.000 49.840 446.000 51.840 ;
        RECT 12.000 48.440 445.600 49.840 ;
        RECT 12.000 24.315 446.000 48.440 ;
      LAYER met4 ;
        RECT 51.535 404.745 88.180 436.905 ;
        RECT 90.580 404.745 91.480 436.905 ;
        RECT 93.880 404.745 180.180 436.905 ;
        RECT 182.580 404.745 183.480 436.905 ;
        RECT 185.880 404.745 272.180 436.905 ;
        RECT 274.580 404.745 275.480 436.905 ;
        RECT 277.880 404.745 364.180 436.905 ;
        RECT 366.580 404.745 367.480 436.905 ;
        RECT 369.880 404.745 407.320 436.905 ;
        RECT 51.535 51.535 407.320 404.745 ;
      LAYER met5 ;
        RECT 52.420 371.180 412.960 404.540 ;
        RECT 52.420 279.180 412.960 363.080 ;
        RECT 52.420 187.180 412.960 271.080 ;
        RECT 52.420 95.180 412.960 179.080 ;
        RECT 52.420 54.640 412.960 87.080 ;
  END
END fpga
END LIBRARY

